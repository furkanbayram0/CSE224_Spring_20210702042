magic
tech sky130A
magscale 1 2
timestamp 1745718357
<< checkpaint >>
rect -3932 -3244 10778 14940
<< viali >>
rect 1409 9605 1443 9639
rect 1777 9605 1811 9639
rect 2237 9537 2271 9571
rect 2053 9401 2087 9435
rect 1869 9129 1903 9163
rect 1501 9061 1535 9095
rect 1685 8925 1719 8959
rect 2053 8925 2087 8959
rect 6469 8925 6503 8959
rect 6285 8789 6319 8823
rect 1409 8449 1443 8483
rect 2145 8449 2179 8483
rect 2329 8449 2363 8483
rect 1593 8313 1627 8347
rect 2329 8313 2363 8347
rect 1685 7837 1719 7871
rect 1501 7701 1535 7735
rect 3341 7429 3375 7463
rect 1409 7361 1443 7395
rect 2237 7361 2271 7395
rect 2421 7361 2455 7395
rect 2513 7361 2547 7395
rect 3617 7361 3651 7395
rect 3525 7293 3559 7327
rect 1593 7225 1627 7259
rect 2329 7225 2363 7259
rect 2697 7157 2731 7191
rect 3341 7157 3375 7191
rect 3801 7157 3835 7191
rect 3157 6885 3191 6919
rect 3801 6885 3835 6919
rect 2789 6817 2823 6851
rect 4261 6817 4295 6851
rect 5089 6817 5123 6851
rect 4169 6749 4203 6783
rect 4997 6749 5031 6783
rect 5181 6749 5215 6783
rect 3249 6613 3283 6647
rect 1593 6409 1627 6443
rect 1409 6273 1443 6307
rect 5917 6273 5951 6307
rect 6009 6273 6043 6307
rect 5733 6069 5767 6103
rect 1593 5865 1627 5899
rect 1409 5661 1443 5695
rect 1409 5185 1443 5219
rect 1869 5185 1903 5219
rect 2053 5185 2087 5219
rect 5549 5185 5583 5219
rect 5641 5117 5675 5151
rect 1593 5049 1627 5083
rect 5181 5049 5215 5083
rect 2237 4981 2271 5015
rect 4445 4777 4479 4811
rect 4905 4777 4939 4811
rect 1593 4709 1627 4743
rect 4537 4641 4571 4675
rect 5549 4641 5583 4675
rect 6009 4641 6043 4675
rect 1409 4573 1443 4607
rect 4445 4573 4479 4607
rect 4721 4573 4755 4607
rect 5917 4573 5951 4607
rect 1961 4097 1995 4131
rect 2237 4097 2271 4131
rect 2421 4097 2455 4131
rect 3157 4097 3191 4131
rect 3341 4097 3375 4131
rect 3433 4097 3467 4131
rect 3525 4097 3559 4131
rect 6193 4097 6227 4131
rect 2099 3961 2133 3995
rect 2973 3961 3007 3995
rect 6009 3961 6043 3995
rect 2329 3893 2363 3927
rect 4813 3689 4847 3723
rect 1501 3621 1535 3655
rect 1685 3485 1719 3519
rect 4537 3485 4571 3519
rect 4629 3485 4663 3519
rect 5917 3145 5951 3179
rect 1685 3009 1719 3043
rect 2053 3009 2087 3043
rect 2145 3009 2179 3043
rect 5825 3009 5859 3043
rect 6009 3009 6043 3043
rect 2329 2873 2363 2907
rect 1501 2805 1535 2839
rect 1869 2805 1903 2839
rect 1685 2465 1719 2499
rect 1409 2397 1443 2431
<< metal1 >>
rect 1104 9818 6808 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 6808 9818
rect 1104 9744 6808 9766
rect 1394 9596 1400 9648
rect 1452 9596 1458 9648
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 5074 9636 5080 9648
rect 1811 9608 5080 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 3418 9568 3424 9580
rect 2271 9540 3424 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 2038 9392 2044 9444
rect 2096 9392 2102 9444
rect 1104 9274 6808 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6808 9274
rect 1104 9200 6808 9222
rect 1118 9120 1124 9172
rect 1176 9160 1182 9172
rect 1857 9163 1915 9169
rect 1857 9160 1869 9163
rect 1176 9132 1869 9160
rect 1176 9120 1182 9132
rect 1857 9129 1869 9132
rect 1903 9129 1915 9163
rect 1857 9123 1915 9129
rect 842 9052 848 9104
rect 900 9092 906 9104
rect 1489 9095 1547 9101
rect 1489 9092 1501 9095
rect 900 9064 1501 9092
rect 900 9052 906 9064
rect 1489 9061 1501 9064
rect 1535 9061 1547 9095
rect 1489 9055 1547 9061
rect 1670 8916 1676 8968
rect 1728 8916 1734 8968
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8956 2099 8959
rect 2958 8956 2964 8968
rect 2087 8928 2964 8956
rect 2087 8925 2099 8928
rect 2041 8919 2099 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 6273 8823 6331 8829
rect 6273 8820 6285 8823
rect 5868 8792 6285 8820
rect 5868 8780 5874 8792
rect 6273 8789 6285 8792
rect 6319 8789 6331 8823
rect 6273 8783 6331 8789
rect 1104 8730 6808 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 6808 8730
rect 1104 8656 6808 8678
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2148 8412 2176 8443
rect 2314 8440 2320 8492
rect 2372 8440 2378 8492
rect 2498 8412 2504 8424
rect 2148 8384 2504 8412
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 1762 8344 1768 8356
rect 1627 8316 1768 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 2317 8347 2375 8353
rect 2317 8313 2329 8347
rect 2363 8344 2375 8347
rect 4062 8344 4068 8356
rect 2363 8316 4068 8344
rect 2363 8313 2375 8316
rect 2317 8307 2375 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 1104 8186 6808 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6808 8186
rect 1104 8112 6808 8134
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 3786 7868 3792 7880
rect 1719 7840 3792 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 1489 7735 1547 7741
rect 1489 7732 1501 7735
rect 900 7704 1501 7732
rect 900 7692 906 7704
rect 1489 7701 1501 7704
rect 1535 7701 1547 7735
rect 1489 7695 1547 7701
rect 1104 7642 6808 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 6808 7642
rect 1104 7568 6808 7590
rect 3329 7463 3387 7469
rect 3329 7460 3341 7463
rect 2240 7432 3341 7460
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 2240 7401 2268 7432
rect 3329 7429 3341 7432
rect 3375 7429 3387 7463
rect 3329 7423 3387 7429
rect 2225 7395 2283 7401
rect 2225 7392 2237 7395
rect 1636 7364 2237 7392
rect 1636 7352 1642 7364
rect 2225 7361 2237 7364
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2314 7352 2320 7404
rect 2372 7392 2378 7404
rect 2409 7395 2467 7401
rect 2409 7392 2421 7395
rect 2372 7364 2421 7392
rect 2372 7352 2378 7364
rect 2409 7361 2421 7364
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 2556 7364 3617 7392
rect 2556 7352 2562 7364
rect 3605 7361 3617 7364
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 3513 7327 3571 7333
rect 3513 7324 3525 7327
rect 2332 7296 3525 7324
rect 2332 7265 2360 7296
rect 3513 7293 3525 7296
rect 3559 7324 3571 7327
rect 4154 7324 4160 7336
rect 3559 7296 4160 7324
rect 3559 7293 3571 7296
rect 3513 7287 3571 7293
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 2317 7259 2375 7265
rect 2317 7256 2329 7259
rect 1627 7228 2329 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 2317 7225 2329 7228
rect 2363 7225 2375 7259
rect 2317 7219 2375 7225
rect 2406 7216 2412 7268
rect 2464 7256 2470 7268
rect 2464 7228 3372 7256
rect 2464 7216 2470 7228
rect 2685 7191 2743 7197
rect 2685 7157 2697 7191
rect 2731 7188 2743 7191
rect 2774 7188 2780 7200
rect 2731 7160 2780 7188
rect 2731 7157 2743 7160
rect 2685 7151 2743 7157
rect 2774 7148 2780 7160
rect 2832 7148 2838 7200
rect 3344 7197 3372 7228
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7157 3387 7191
rect 3329 7151 3387 7157
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3789 7191 3847 7197
rect 3789 7188 3801 7191
rect 3568 7160 3801 7188
rect 3568 7148 3574 7160
rect 3789 7157 3801 7160
rect 3835 7157 3847 7191
rect 3789 7151 3847 7157
rect 1104 7098 6808 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6808 7098
rect 1104 7024 6808 7046
rect 3142 6876 3148 6928
rect 3200 6916 3206 6928
rect 3510 6916 3516 6928
rect 3200 6888 3516 6916
rect 3200 6876 3206 6888
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 3786 6876 3792 6928
rect 3844 6876 3850 6928
rect 2774 6808 2780 6860
rect 2832 6808 2838 6860
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4249 6851 4307 6857
rect 4249 6848 4261 6851
rect 4120 6820 4261 6848
rect 4120 6808 4126 6820
rect 4249 6817 4261 6820
rect 4295 6817 4307 6851
rect 4249 6811 4307 6817
rect 5074 6808 5080 6860
rect 5132 6808 5138 6860
rect 4154 6740 4160 6792
rect 4212 6740 4218 6792
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6780 5227 6783
rect 5902 6780 5908 6792
rect 5215 6752 5908 6780
rect 5215 6749 5227 6752
rect 5169 6743 5227 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 6454 6644 6460 6656
rect 3283 6616 6460 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 1104 6554 6808 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 6808 6554
rect 1104 6480 6808 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1854 6440 1860 6452
rect 1627 6412 1860 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1854 6400 1860 6412
rect 1912 6440 1918 6452
rect 2498 6440 2504 6452
rect 1912 6412 2504 6440
rect 1912 6400 1918 6412
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5905 6307 5963 6313
rect 5905 6304 5917 6307
rect 5684 6276 5917 6304
rect 5684 6264 5690 6276
rect 5905 6273 5917 6276
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 5994 6264 6000 6316
rect 6052 6264 6058 6316
rect 5718 6060 5724 6112
rect 5776 6060 5782 6112
rect 1104 6010 6808 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6808 6010
rect 1104 5936 6808 5958
rect 1578 5856 1584 5908
rect 1636 5856 1642 5908
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1104 5466 6808 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 6808 5466
rect 1104 5392 6808 5414
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1854 5176 1860 5228
rect 1912 5176 1918 5228
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 2004 5188 2053 5216
rect 2004 5176 2010 5188
rect 2041 5185 2053 5188
rect 2087 5216 2099 5219
rect 2314 5216 2320 5228
rect 2087 5188 2320 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 4488 5188 5549 5216
rect 4488 5176 4494 5188
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5902 5148 5908 5160
rect 5675 5120 5908 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5080 1639 5083
rect 2406 5080 2412 5092
rect 1627 5052 2412 5080
rect 1627 5049 1639 5052
rect 1581 5043 1639 5049
rect 2406 5040 2412 5052
rect 2464 5040 2470 5092
rect 5166 5040 5172 5092
rect 5224 5040 5230 5092
rect 2225 5015 2283 5021
rect 2225 4981 2237 5015
rect 2271 5012 2283 5015
rect 3326 5012 3332 5024
rect 2271 4984 3332 5012
rect 2271 4981 2283 4984
rect 2225 4975 2283 4981
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 1104 4922 6808 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6808 4922
rect 1104 4848 6808 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 4430 4808 4436 4820
rect 1820 4780 4436 4808
rect 1820 4768 1826 4780
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 5994 4808 6000 4820
rect 4939 4780 6000 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 1627 4712 5948 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 2406 4632 2412 4684
rect 2464 4672 2470 4684
rect 4525 4675 4583 4681
rect 4525 4672 4537 4675
rect 2464 4644 4537 4672
rect 2464 4632 2470 4644
rect 4525 4641 4537 4644
rect 4571 4641 4583 4675
rect 4525 4635 4583 4641
rect 5534 4632 5540 4684
rect 5592 4632 5598 4684
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 900 4576 1409 4604
rect 900 4564 906 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3970 4604 3976 4616
rect 3200 4576 3976 4604
rect 3200 4564 3206 4576
rect 3970 4564 3976 4576
rect 4028 4604 4034 4616
rect 5920 4613 5948 4712
rect 5994 4632 6000 4684
rect 6052 4632 6058 4684
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4028 4576 4445 4604
rect 4028 4564 4034 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 4433 4567 4491 4573
rect 4540 4576 4721 4604
rect 4540 4548 4568 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 4522 4496 4528 4548
rect 4580 4496 4586 4548
rect 1104 4378 6808 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 6808 4378
rect 1104 4304 6808 4326
rect 3142 4264 3148 4276
rect 2792 4236 3148 4264
rect 2792 4196 2820 4236
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 2332 4168 2820 4196
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2332 4128 2360 4168
rect 2271 4100 2360 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 1964 4060 1992 4091
rect 2406 4088 2412 4140
rect 2464 4088 2470 4140
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3160 4060 3188 4091
rect 3326 4088 3332 4140
rect 3384 4088 3390 4140
rect 3418 4088 3424 4140
rect 3476 4088 3482 4140
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 4062 4128 4068 4140
rect 3559 4100 4068 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 6178 4088 6184 4140
rect 6236 4088 6242 4140
rect 5718 4060 5724 4072
rect 1964 4032 3096 4060
rect 3160 4032 5724 4060
rect 1762 3952 1768 4004
rect 1820 3992 1826 4004
rect 2087 3995 2145 4001
rect 2087 3992 2099 3995
rect 1820 3964 2099 3992
rect 1820 3952 1826 3964
rect 2087 3961 2099 3964
rect 2133 3961 2145 3995
rect 2087 3955 2145 3961
rect 2958 3952 2964 4004
rect 3016 3952 3022 4004
rect 3068 3992 3096 4032
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 4522 3992 4528 4004
rect 3068 3964 4528 3992
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 5997 3995 6055 4001
rect 5997 3992 6009 3995
rect 4764 3964 6009 3992
rect 4764 3952 4770 3964
rect 5997 3961 6009 3964
rect 6043 3961 6055 3995
rect 5997 3955 6055 3961
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 5626 3924 5632 3936
rect 2363 3896 5632 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 1104 3834 6808 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6808 3834
rect 1104 3760 6808 3782
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 4706 3720 4712 3732
rect 1728 3692 4712 3720
rect 1728 3680 1734 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 4801 3723 4859 3729
rect 4801 3689 4813 3723
rect 4847 3720 4859 3723
rect 4982 3720 4988 3732
rect 4847 3692 4988 3720
rect 4847 3689 4859 3692
rect 4801 3683 4859 3689
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 842 3612 848 3664
rect 900 3652 906 3664
rect 1489 3655 1547 3661
rect 1489 3652 1501 3655
rect 900 3624 1501 3652
rect 900 3612 906 3624
rect 1489 3621 1501 3624
rect 1535 3621 1547 3655
rect 1489 3615 1547 3621
rect 1762 3612 1768 3664
rect 1820 3652 1826 3664
rect 6178 3652 6184 3664
rect 1820 3624 6184 3652
rect 1820 3612 1826 3624
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 5534 3584 5540 3596
rect 1688 3556 5540 3584
rect 1688 3525 1716 3556
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 4632 3448 4660 3479
rect 4028 3420 4660 3448
rect 4028 3408 4034 3420
rect 1104 3290 6808 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 6808 3290
rect 1104 3216 6808 3238
rect 5810 3176 5816 3188
rect 1688 3148 5816 3176
rect 1688 3049 1716 3148
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 5902 3136 5908 3188
rect 5960 3136 5966 3188
rect 5166 3108 5172 3120
rect 2056 3080 5172 3108
rect 2056 3049 2084 3080
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 1118 2932 1124 2984
rect 1176 2972 1182 2984
rect 2148 2972 2176 3003
rect 3970 3000 3976 3052
rect 4028 3040 4034 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 4028 3012 5825 3040
rect 4028 3000 4034 3012
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 4522 2972 4528 2984
rect 1176 2944 2176 2972
rect 2332 2944 4528 2972
rect 1176 2932 1182 2944
rect 2332 2913 2360 2944
rect 4522 2932 4528 2944
rect 4580 2972 4586 2984
rect 6012 2972 6040 3003
rect 4580 2944 6040 2972
rect 4580 2932 4586 2944
rect 2317 2907 2375 2913
rect 2317 2873 2329 2907
rect 2363 2873 2375 2907
rect 2317 2867 2375 2873
rect 1486 2796 1492 2848
rect 1544 2796 1550 2848
rect 1854 2796 1860 2848
rect 1912 2796 1918 2848
rect 1104 2746 6808 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6808 2746
rect 1104 2672 6808 2694
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 1762 2496 1768 2508
rect 1719 2468 1768 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 1762 2456 1768 2468
rect 1820 2456 1826 2508
rect 1394 2388 1400 2440
rect 1452 2388 1458 2440
rect 1104 2202 6808 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 6808 2202
rect 1104 2128 6808 2150
<< via1 >>
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 1400 9639 1452 9648
rect 1400 9605 1409 9639
rect 1409 9605 1443 9639
rect 1443 9605 1452 9639
rect 1400 9596 1452 9605
rect 5080 9596 5132 9648
rect 3424 9528 3476 9580
rect 2044 9435 2096 9444
rect 2044 9401 2053 9435
rect 2053 9401 2087 9435
rect 2087 9401 2096 9435
rect 2044 9392 2096 9401
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 1124 9120 1176 9172
rect 848 9052 900 9104
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 2964 8916 3016 8968
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 5816 8780 5868 8832
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 2504 8372 2556 8424
rect 1768 8304 1820 8356
rect 4068 8304 4120 8356
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 3792 7828 3844 7880
rect 848 7692 900 7744
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1584 7352 1636 7404
rect 2320 7352 2372 7404
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 4160 7284 4212 7336
rect 2412 7216 2464 7268
rect 2780 7148 2832 7200
rect 3516 7148 3568 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 3148 6919 3200 6928
rect 3148 6885 3157 6919
rect 3157 6885 3191 6919
rect 3191 6885 3200 6919
rect 3148 6876 3200 6885
rect 3516 6876 3568 6928
rect 3792 6919 3844 6928
rect 3792 6885 3801 6919
rect 3801 6885 3835 6919
rect 3835 6885 3844 6919
rect 3792 6876 3844 6885
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 2780 6808 2832 6817
rect 4068 6808 4120 6860
rect 5080 6851 5132 6860
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4988 6783 5040 6792
rect 4988 6749 4997 6783
rect 4997 6749 5031 6783
rect 5031 6749 5040 6783
rect 4988 6740 5040 6749
rect 5908 6740 5960 6792
rect 6460 6604 6512 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 1860 6400 1912 6452
rect 2504 6400 2556 6452
rect 848 6264 900 6316
rect 5632 6264 5684 6316
rect 6000 6307 6052 6316
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 848 5176 900 5228
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 1952 5176 2004 5228
rect 2320 5176 2372 5228
rect 4436 5176 4488 5228
rect 5908 5108 5960 5160
rect 2412 5040 2464 5092
rect 5172 5083 5224 5092
rect 5172 5049 5181 5083
rect 5181 5049 5215 5083
rect 5215 5049 5224 5083
rect 5172 5040 5224 5049
rect 3332 4972 3384 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 1768 4768 1820 4820
rect 4436 4811 4488 4820
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 6000 4768 6052 4820
rect 2412 4632 2464 4684
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 848 4564 900 4616
rect 3148 4564 3200 4616
rect 3976 4564 4028 4616
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 4528 4496 4580 4548
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 3148 4224 3200 4276
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3424 4131 3476 4140
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 3424 4088 3476 4097
rect 4068 4088 4120 4140
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 1768 3952 1820 4004
rect 2964 3995 3016 4004
rect 2964 3961 2973 3995
rect 2973 3961 3007 3995
rect 3007 3961 3016 3995
rect 2964 3952 3016 3961
rect 5724 4020 5776 4072
rect 4528 3952 4580 4004
rect 4712 3952 4764 4004
rect 5632 3884 5684 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 1676 3680 1728 3732
rect 4712 3680 4764 3732
rect 4988 3680 5040 3732
rect 848 3612 900 3664
rect 1768 3612 1820 3664
rect 6184 3612 6236 3664
rect 5540 3544 5592 3596
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 3976 3408 4028 3460
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 5816 3136 5868 3188
rect 5908 3179 5960 3188
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 5172 3068 5224 3120
rect 1124 2932 1176 2984
rect 3976 3000 4028 3052
rect 4528 2932 4580 2984
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 1768 2456 1820 2508
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1412 9654 1440 10911
rect 2042 10296 2098 10305
rect 2042 10231 2098 10240
rect 1400 9648 1452 9654
rect 1122 9616 1178 9625
rect 1400 9590 1452 9596
rect 1122 9551 1178 9560
rect 1136 9178 1164 9551
rect 2056 9450 2084 10231
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 1124 9172 1176 9178
rect 1124 9114 1176 9120
rect 848 9104 900 9110
rect 846 9072 848 9081
rect 900 9072 902 9081
rect 846 9007 902 9016
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 848 7744 900 7750
rect 846 7712 848 7721
rect 900 7712 902 7721
rect 846 7647 902 7656
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1412 6905 1440 7346
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1596 5914 1624 7346
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5001 888 5170
rect 846 4992 902 5001
rect 846 4927 902 4936
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 860 4321 888 4558
rect 846 4312 902 4321
rect 846 4247 902 4256
rect 1688 3738 1716 8910
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1780 4826 1808 8298
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2332 7410 2360 8434
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2516 7410 2544 8366
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2332 7290 2360 7346
rect 2332 7274 2452 7290
rect 2332 7268 2464 7274
rect 2332 7262 2412 7268
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1872 5234 1900 6394
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2332 5234 2360 7262
rect 2412 7210 2464 7216
rect 2516 6458 2544 7346
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6866 2820 7142
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 1964 5114 1992 5170
rect 1872 5086 1992 5114
rect 2412 5092 2464 5098
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1780 4010 1808 4762
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 1872 3890 1900 5086
rect 2412 5034 2464 5040
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2424 4690 2452 5034
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2424 4146 2452 4626
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2976 4010 3004 8910
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3160 4622 3188 6870
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3160 4282 3188 4558
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3344 4146 3372 4966
rect 3436 4146 3464 9522
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 6934 3556 7142
rect 3804 6934 3832 7822
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3792 6928 3844 6934
rect 3792 6870 3844 6876
rect 4080 6866 4108 8298
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 1780 3862 1900 3890
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1780 3670 1808 3862
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 848 3664 900 3670
rect 846 3632 848 3641
rect 1768 3664 1820 3670
rect 900 3632 902 3641
rect 1768 3606 1820 3612
rect 846 3567 902 3576
rect 1124 2984 1176 2990
rect 1124 2926 1176 2932
rect 1136 2825 1164 2926
rect 1492 2848 1544 2854
rect 1122 2816 1178 2825
rect 1492 2790 1544 2796
rect 1122 2751 1178 2760
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 785 1440 2382
rect 1504 1465 1532 2790
rect 1780 2514 1808 3606
rect 3988 3466 4016 4558
rect 4080 4146 4108 6802
rect 4172 6798 4200 7278
rect 5092 6866 5120 9590
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4448 4826 4476 5170
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4540 4010 4568 4490
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4540 3534 4568 3946
rect 4724 3738 4752 3946
rect 5000 3738 5028 6734
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 3988 3058 4016 3402
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4540 2990 4568 3470
rect 5184 3126 5212 5034
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5552 3602 5580 4626
rect 5644 3942 5672 6258
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 4078 5764 6054
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5828 3194 5856 8774
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 5166 5948 6734
rect 6472 6662 6500 8910
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 3194 5948 5102
rect 6012 4826 6040 6258
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6012 4690 6040 4762
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6196 3670 6224 4082
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 1872 2145 1900 2790
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 1858 2136 1914 2145
rect 2610 2139 2918 2148
rect 1858 2071 1914 2080
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 1398 776 1454 785
rect 1398 711 1454 720
<< via2 >>
rect 1398 10920 1454 10976
rect 2042 10240 2098 10296
rect 1122 9560 1178 9616
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 846 9052 848 9072
rect 848 9052 900 9072
rect 900 9052 902 9072
rect 846 9016 902 9052
rect 1398 8200 1454 8256
rect 846 7692 848 7712
rect 848 7692 900 7712
rect 900 7692 902 7712
rect 846 7656 902 7692
rect 1398 6840 1454 6896
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 1398 5480 1454 5536
rect 846 4936 902 4992
rect 846 4256 902 4312
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 846 3612 848 3632
rect 848 3612 900 3632
rect 900 3612 902 3632
rect 846 3576 902 3612
rect 1122 2760 1178 2816
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1858 2080 1914 2136
rect 1490 1400 1546 1456
rect 1398 720 1454 776
<< metal3 >>
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 0 10298 800 10328
rect 2037 10298 2103 10301
rect 0 10296 2103 10298
rect 0 10240 2042 10296
rect 2098 10240 2103 10296
rect 0 10238 2103 10240
rect 0 10208 800 10238
rect 2037 10235 2103 10238
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 0 9618 800 9648
rect 1117 9618 1183 9621
rect 0 9616 1183 9618
rect 0 9560 1122 9616
rect 1178 9560 1183 9616
rect 0 9558 1183 9560
rect 0 9528 800 9558
rect 1117 9555 1183 9558
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 0 8848 800 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 0 7488 800 7518
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 0 6128 800 6158
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 0 4768 800 4798
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 841 4314 907 4317
rect 798 4312 907 4314
rect 798 4256 846 4312
rect 902 4256 907 4312
rect 798 4251 907 4256
rect 798 4208 858 4251
rect 0 4118 858 4208
rect 0 4088 800 4118
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 0 3408 800 3438
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 0 2818 800 2848
rect 1117 2818 1183 2821
rect 0 2816 1183 2818
rect 0 2760 1122 2816
rect 1178 2760 1183 2816
rect 0 2758 1183 2760
rect 0 2728 800 2758
rect 1117 2755 1183 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 2606 2208 2922 2209
rect 0 2138 800 2168
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 1853 2138 1919 2141
rect 0 2136 1919 2138
rect 0 2080 1858 2136
rect 1914 2080 1919 2136
rect 0 2078 1919 2080
rect 0 2048 800 2078
rect 1853 2075 1919 2078
rect 0 1458 800 1488
rect 1485 1458 1551 1461
rect 0 1456 1551 1458
rect 0 1400 1490 1456
rect 1546 1400 1551 1456
rect 0 1398 1551 1400
rect 0 1368 800 1398
rect 1485 1395 1551 1398
rect 0 778 800 808
rect 1393 778 1459 781
rect 0 776 1459 778
rect 0 720 1398 776
rect 1454 720 1459 776
rect 0 718 1459 720
rect 0 688 800 718
rect 1393 715 1459 718
<< via3 >>
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9840
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 9824 2924 9840
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8736 2924 9760
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform -1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _11_
timestamp 0
transform -1 0 4416 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _12_
timestamp 0
transform -1 0 2760 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _13_
timestamp 0
transform 1 0 3312 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _14_
timestamp 0
transform 1 0 2760 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 0
transform 1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _16_
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _17_
timestamp 0
transform 1 0 4416 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 0
transform 1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _19_
timestamp 0
transform -1 0 5796 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _20_
timestamp 0
transform 1 0 4416 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _21_
timestamp 0
transform 1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform -1 0 6164 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform 1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _24_
timestamp 0
transform -1 0 6164 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _25_
timestamp 0
transform 1 0 1840 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _26_
timestamp 0
transform 1 0 3312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 0
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_13
timestamp 0
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 0
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_14
timestamp 0
transform 1 0 2392 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_26
timestamp 0
transform 1 0 3496 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_38
timestamp 0
transform 1 0 4600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_50
timestamp 0
transform 1 0 5704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 0
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_7
timestamp 0
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 0
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_35
timestamp 0
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_19
timestamp 0
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_23
timestamp 0
transform 1 0 3220 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 0
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 0
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 0
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_35
timestamp 0
transform 1 0 4324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_42
timestamp 0
transform 1 0 4968 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_55
timestamp 0
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_6
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_13
timestamp 0
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_25
timestamp 0
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_37
timestamp 0
transform 1 0 4508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_43
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_6
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_18
timestamp 0
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_30
timestamp 0
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_42
timestamp 0
transform 1 0 4968 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_24
timestamp 0
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_36
timestamp 0
transform 1 0 4416 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_45
timestamp 0
transform 1 0 5244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_57
timestamp 0
transform 1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_6
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_10
timestamp 0
transform 1 0 2024 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_18
timestamp 0
transform 1 0 2760 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_31
timestamp 0
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_43
timestamp 0
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_7
timestamp 0
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_19
timestamp 0
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_6
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_10
timestamp 0
transform 1 0 2024 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_14
timestamp 0
transform 1 0 2392 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_26
timestamp 0
transform 1 0 3496 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_38
timestamp 0
transform 1 0 4600 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_50
timestamp 0
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_11
timestamp 0
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_23
timestamp 0
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_13
timestamp 0
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_25
timestamp 0
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_29
timestamp 0
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 0
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 0
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform -1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 0
transform -1 0 1932 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform -1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_14
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_15
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_16
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_17
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_18
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_19
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_20
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_21
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_22
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_23
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_24
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_25
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 6808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_26
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_27
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 6808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_30
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_31
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_32
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_33
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_34
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_35
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_36
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_37
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_38
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_39
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_40
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_41
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_42
timestamp 0
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_43
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
<< labels >>
rlabel metal1 s 3956 9792 3956 9792 4 VGND
rlabel metal1 s 3956 9248 3956 9248 4 VPWR
rlabel metal1 s 3818 4114 3818 4114 4 _00_
rlabel metal1 s 2760 7174 2760 7174 4 _01_
rlabel metal1 s 3818 4590 3818 4590 4 _02_
rlabel metal1 s 4876 6630 4876 6630 4 _03_
rlabel metal1 s 5796 5134 5796 5134 4 _04_
rlabel metal1 s 4922 3706 4922 3706 4 _05_
rlabel metal2 s 6026 5474 6026 5474 4 _06_
rlabel metal1 s 4002 3910 4002 3910 4 _07_
rlabel metal1 s 3174 4080 3174 4080 4 _08_
rlabel metal2 s 3358 4556 3358 4556 4 _09_
rlabel metal3 s 1050 748 1050 748 4 in[0]
rlabel metal3 s 0 6128 800 6248 4 in[1]
port 4 nsew
rlabel metal3 s 1050 6868 1050 6868 4 in[2]
rlabel metal3 s 1050 5508 1050 5508 4 in[3]
rlabel metal3 s 912 2788 912 2788 4 in[4]
rlabel metal3 s 1050 8228 1050 8228 4 in[5]
rlabel metal3 s 0 4768 800 4888 4 in[6]
port 9 nsew
rlabel metal3 s 0 4088 800 4208 4 in[7]
port 10 nsew
rlabel metal1 s 2024 5202 2024 5202 4 net1
rlabel metal1 s 2852 9554 2852 9554 4 net10
rlabel metal2 s 3818 7378 3818 7378 4 net11
rlabel metal1 s 3772 3162 3772 3162 4 net12
rlabel metal1 s 3450 9622 3450 9622 4 net13
rlabel metal1 s 2070 3060 2070 3060 4 net14
rlabel metal1 s 2530 8942 2530 8942 4 net15
rlabel metal1 s 1702 3536 1702 3536 4 net16
rlabel metal1 s 2070 6426 2070 6426 4 net2
rlabel metal1 s 3864 7310 3864 7310 4 net3
rlabel metal1 s 1932 7378 1932 7378 4 net4
rlabel metal2 s 4554 3230 4554 3230 4 net5
rlabel metal1 s 1955 3978 1955 3978 4 net6
rlabel metal2 s 2438 4590 2438 4590 4 net7
rlabel metal1 s 5934 4658 5934 4658 4 net8
rlabel metal1 s 5382 3978 5382 3978 4 net9
rlabel metal3 s 0 8848 800 8968 4 out[0]
port 11 nsew
rlabel metal2 s 2070 9843 2070 9843 4 out[1]
rlabel metal3 s 0 7488 800 7608 4 out[2]
port 13 nsew
rlabel metal3 s 1096 1428 1096 1428 4 out[3]
rlabel metal3 s 1050 10948 1050 10948 4 out[4]
rlabel metal3 s 1280 2108 1280 2108 4 out[5]
rlabel metal1 s 1518 9146 1518 9146 4 out[6]
rlabel metal3 s 0 3408 800 3528 4 out[7]
port 18 nsew
flabel metal4 s 2604 2128 2924 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1944 2128 2264 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 688 800 808 0 FreeSans 600 0 0 0 in[0]
port 3 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 in[1]
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 in[2]
port 5 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 in[3]
port 6 nsew
flabel metal3 s 0 2728 800 2848 0 FreeSans 600 0 0 0 in[4]
port 7 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 in[5]
port 8 nsew
flabel metal3 s 400 4828 400 4828 0 FreeSans 600 0 0 0 in[6]
flabel metal3 s 400 4148 400 4148 0 FreeSans 600 0 0 0 in[7]
flabel metal3 s 400 8908 400 8908 0 FreeSans 600 0 0 0 out[0]
flabel metal3 s 0 10208 800 10328 0 FreeSans 600 0 0 0 out[1]
port 12 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 out[2]
flabel metal3 s 0 1368 800 1488 0 FreeSans 600 0 0 0 out[3]
port 14 nsew
flabel metal3 s 0 10888 800 11008 0 FreeSans 600 0 0 0 out[4]
port 15 nsew
flabel metal3 s 0 2048 800 2168 0 FreeSans 600 0 0 0 out[5]
port 16 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 out[6]
port 17 nsew
flabel metal3 s 400 3468 400 3468 0 FreeSans 600 0 0 0 out[7]
<< properties >>
string FIXED_BBOX 0 0 8000 12000
<< end >>
