magic
tech sky130A
magscale 1 2
timestamp 1747871253
<< checkpaint >>
rect -3932 -2836 19932 20380
<< viali >>
rect 9597 15657 9631 15691
rect 10517 15589 10551 15623
rect 8309 15521 8343 15555
rect 13093 15521 13127 15555
rect 14197 15521 14231 15555
rect 4077 15453 4111 15487
rect 4261 15453 4295 15487
rect 4537 15453 4571 15487
rect 8585 15453 8619 15487
rect 9505 15453 9539 15487
rect 10333 15453 10367 15487
rect 14289 15453 14323 15487
rect 12541 15385 12575 15419
rect 12725 15385 12759 15419
rect 12817 15385 12851 15419
rect 2421 15317 2455 15351
rect 2789 15317 2823 15351
rect 3893 15317 3927 15351
rect 6837 15317 6871 15351
rect 12449 15317 12483 15351
rect 12909 15317 12943 15351
rect 13369 15317 13403 15351
rect 13921 15317 13955 15351
rect 6653 15113 6687 15147
rect 7205 15113 7239 15147
rect 10977 15113 11011 15147
rect 14013 15113 14047 15147
rect 6837 15045 6871 15079
rect 12265 15045 12299 15079
rect 1593 14977 1627 15011
rect 1869 14977 1903 15011
rect 2053 14977 2087 15011
rect 5549 14977 5583 15011
rect 5733 14977 5767 15011
rect 7021 14977 7055 15011
rect 7113 14977 7147 15011
rect 10793 14977 10827 15011
rect 11069 14977 11103 15011
rect 11713 14977 11747 15011
rect 11989 14977 12023 15011
rect 14473 14977 14507 15011
rect 4261 14909 4295 14943
rect 4537 14909 4571 14943
rect 1961 14841 1995 14875
rect 11805 14841 11839 14875
rect 2513 14773 2547 14807
rect 2789 14773 2823 14807
rect 5365 14773 5399 14807
rect 5641 14773 5675 14807
rect 7665 14773 7699 14807
rect 10333 14773 10367 14807
rect 10793 14773 10827 14807
rect 11621 14773 11655 14807
rect 1593 14569 1627 14603
rect 10977 14569 11011 14603
rect 2973 14501 3007 14535
rect 5457 14433 5491 14467
rect 5733 14433 5767 14467
rect 12817 14433 12851 14467
rect 2053 14365 2087 14399
rect 8953 14365 8987 14399
rect 11345 14365 11379 14399
rect 1409 14297 1443 14331
rect 1625 14297 1659 14331
rect 9229 14297 9263 14331
rect 1777 14229 1811 14263
rect 2605 14229 2639 14263
rect 3985 14229 4019 14263
rect 10701 14229 10735 14263
rect 11713 14229 11747 14263
rect 13277 14229 13311 14263
rect 13829 14229 13863 14263
rect 14473 14229 14507 14263
rect 1593 14025 1627 14059
rect 8493 14025 8527 14059
rect 9505 14025 9539 14059
rect 12633 14025 12667 14059
rect 2053 13957 2087 13991
rect 8125 13957 8159 13991
rect 8341 13957 8375 13991
rect 9137 13957 9171 13991
rect 9353 13957 9387 13991
rect 13001 13957 13035 13991
rect 14013 13957 14047 13991
rect 1409 13889 1443 13923
rect 1961 13889 1995 13923
rect 2237 13889 2271 13923
rect 4353 13889 4387 13923
rect 4537 13889 4571 13923
rect 5917 13889 5951 13923
rect 6561 13889 6595 13923
rect 8953 13889 8987 13923
rect 11713 13889 11747 13923
rect 12725 13889 12759 13923
rect 13185 13889 13219 13923
rect 13277 13889 13311 13923
rect 13461 13889 13495 13923
rect 14197 13889 14231 13923
rect 2329 13821 2363 13855
rect 7113 13821 7147 13855
rect 13369 13821 13403 13855
rect 14381 13821 14415 13855
rect 2237 13753 2271 13787
rect 4721 13753 4755 13787
rect 6009 13753 6043 13787
rect 4089 13685 4123 13719
rect 4997 13685 5031 13719
rect 8309 13685 8343 13719
rect 9321 13685 9355 13719
rect 12357 13685 12391 13719
rect 13921 13685 13955 13719
rect 4077 13481 4111 13515
rect 4537 13481 4571 13515
rect 4721 13481 4755 13515
rect 11897 13481 11931 13515
rect 13829 13481 13863 13515
rect 2329 13413 2363 13447
rect 7573 13413 7607 13447
rect 3985 13345 4019 13379
rect 7205 13345 7239 13379
rect 11069 13345 11103 13379
rect 12081 13345 12115 13379
rect 1961 13277 1995 13311
rect 2789 13277 2823 13311
rect 3617 13277 3651 13311
rect 3893 13277 3927 13311
rect 5089 13277 5123 13311
rect 7297 13277 7331 13311
rect 7573 13277 7607 13311
rect 7941 13277 7975 13311
rect 11805 13277 11839 13311
rect 11989 13277 12023 13311
rect 14105 13277 14139 13311
rect 2605 13209 2639 13243
rect 4353 13209 4387 13243
rect 5181 13209 5215 13243
rect 6929 13209 6963 13243
rect 8677 13209 8711 13243
rect 10793 13209 10827 13243
rect 12357 13209 12391 13243
rect 14197 13209 14231 13243
rect 1869 13141 1903 13175
rect 2973 13141 3007 13175
rect 4261 13141 4295 13175
rect 4563 13141 4597 13175
rect 7389 13141 7423 13175
rect 9321 13141 9355 13175
rect 11437 13141 11471 13175
rect 3617 12937 3651 12971
rect 6193 12937 6227 12971
rect 6929 12937 6963 12971
rect 14105 12937 14139 12971
rect 3801 12869 3835 12903
rect 4001 12869 4035 12903
rect 9045 12869 9079 12903
rect 4629 12801 4663 12835
rect 5181 12801 5215 12835
rect 6009 12801 6043 12835
rect 6193 12801 6227 12835
rect 6561 12801 6595 12835
rect 6745 12801 6779 12835
rect 8585 12801 8619 12835
rect 8767 12801 8801 12835
rect 11713 12801 11747 12835
rect 12449 12801 12483 12835
rect 14197 12801 14231 12835
rect 4169 12665 4203 12699
rect 4537 12665 4571 12699
rect 5825 12665 5859 12699
rect 7297 12665 7331 12699
rect 8953 12665 8987 12699
rect 11989 12665 12023 12699
rect 12265 12665 12299 12699
rect 3985 12597 4019 12631
rect 4721 12597 4755 12631
rect 10333 12597 10367 12631
rect 11621 12597 11655 12631
rect 13185 12597 13219 12631
rect 14381 12597 14415 12631
rect 3617 12393 3651 12427
rect 10425 12393 10459 12427
rect 12541 12393 12575 12427
rect 13277 12393 13311 12427
rect 11529 12325 11563 12359
rect 4353 12257 4387 12291
rect 6469 12257 6503 12291
rect 13645 12257 13679 12291
rect 6377 12189 6411 12223
rect 10149 12189 10183 12223
rect 10793 12189 10827 12223
rect 12173 12189 12207 12223
rect 12725 12189 12759 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 13553 12189 13587 12223
rect 6101 12121 6135 12155
rect 8217 12121 8251 12155
rect 9137 12121 9171 12155
rect 13461 12121 13495 12155
rect 10241 12053 10275 12087
rect 10425 12053 10459 12087
rect 11069 12053 11103 12087
rect 11805 12053 11839 12087
rect 13093 12053 13127 12087
rect 13261 12053 13295 12087
rect 14473 12053 14507 12087
rect 3249 11849 3283 11883
rect 3709 11849 3743 11883
rect 4169 11849 4203 11883
rect 11805 11849 11839 11883
rect 12081 11849 12115 11883
rect 13001 11849 13035 11883
rect 4721 11781 4755 11815
rect 5181 11781 5215 11815
rect 6561 11781 6595 11815
rect 12449 11781 12483 11815
rect 2789 11713 2823 11747
rect 3308 11713 3342 11747
rect 3525 11713 3559 11747
rect 3801 11713 3835 11747
rect 4537 11713 4571 11747
rect 4629 11713 4663 11747
rect 5825 11713 5859 11747
rect 6469 11713 6503 11747
rect 6745 11713 6779 11747
rect 7113 11713 7147 11747
rect 7205 11713 7239 11747
rect 8953 11713 8987 11747
rect 11345 11713 11379 11747
rect 11713 11713 11747 11747
rect 11897 11713 11931 11747
rect 6929 11645 6963 11679
rect 8493 11645 8527 11679
rect 8744 11645 8778 11679
rect 8861 11645 8895 11679
rect 9229 11645 9263 11679
rect 9321 11645 9355 11679
rect 9597 11645 9631 11679
rect 2881 11577 2915 11611
rect 11529 11577 11563 11611
rect 2697 11509 2731 11543
rect 3433 11509 3467 11543
rect 3525 11509 3559 11543
rect 5733 11509 5767 11543
rect 7573 11509 7607 11543
rect 8585 11509 8619 11543
rect 13369 11509 13403 11543
rect 8953 11305 8987 11339
rect 3985 11237 4019 11271
rect 4077 11237 4111 11271
rect 6653 11237 6687 11271
rect 13001 11237 13035 11271
rect 3801 11169 3835 11203
rect 4537 11169 4571 11203
rect 10701 11169 10735 11203
rect 11437 11169 11471 11203
rect 12449 11169 12483 11203
rect 4077 11101 4111 11135
rect 6653 11101 6687 11135
rect 6929 11101 6963 11135
rect 7573 11101 7607 11135
rect 8125 11101 8159 11135
rect 12633 11101 12667 11135
rect 13093 11101 13127 11135
rect 13185 11101 13219 11135
rect 13369 11101 13403 11135
rect 13737 11101 13771 11135
rect 3249 11033 3283 11067
rect 4813 11033 4847 11067
rect 6561 11033 6595 11067
rect 6837 11033 6871 11067
rect 8493 11033 8527 11067
rect 10425 11033 10459 11067
rect 12817 11033 12851 11067
rect 14473 11033 14507 11067
rect 3157 10965 3191 10999
rect 7205 10965 7239 10999
rect 8033 10965 8067 10999
rect 2421 10761 2455 10795
rect 3341 10761 3375 10795
rect 3709 10761 3743 10795
rect 5089 10761 5123 10795
rect 5273 10761 5307 10795
rect 5641 10761 5675 10795
rect 12081 10761 12115 10795
rect 14381 10761 14415 10795
rect 2145 10693 2179 10727
rect 7449 10693 7483 10727
rect 7665 10693 7699 10727
rect 10241 10693 10275 10727
rect 12357 10693 12391 10727
rect 2237 10625 2271 10659
rect 2421 10625 2455 10659
rect 3157 10625 3191 10659
rect 3341 10625 3375 10659
rect 6193 10625 6227 10659
rect 7205 10625 7239 10659
rect 9999 10625 10033 10659
rect 12449 10625 12483 10659
rect 12541 10625 12575 10659
rect 12725 10625 12759 10659
rect 13001 10625 13035 10659
rect 13461 10625 13495 10659
rect 14197 10625 14231 10659
rect 14473 10625 14507 10659
rect 4905 10557 4939 10591
rect 4997 10557 5031 10591
rect 5365 10557 5399 10591
rect 5457 10557 5491 10591
rect 9597 10557 9631 10591
rect 9689 10557 9723 10591
rect 13737 10557 13771 10591
rect 6009 10489 6043 10523
rect 7297 10489 7331 10523
rect 12541 10489 12575 10523
rect 2789 10421 2823 10455
rect 7481 10421 7515 10455
rect 11805 10421 11839 10455
rect 14013 10421 14047 10455
rect 10425 10217 10459 10251
rect 13001 10217 13035 10251
rect 13369 10217 13403 10251
rect 13645 10217 13679 10251
rect 3341 10149 3375 10183
rect 6561 10081 6595 10115
rect 6837 10081 6871 10115
rect 13001 10081 13035 10115
rect 9965 10013 9999 10047
rect 10241 10013 10275 10047
rect 10425 10013 10459 10047
rect 10517 10013 10551 10047
rect 10977 10013 11011 10047
rect 12081 10013 12115 10047
rect 12449 10013 12483 10047
rect 12725 10013 12759 10047
rect 13185 10013 13219 10047
rect 12909 9945 12943 9979
rect 8309 9877 8343 9911
rect 9689 9877 9723 9911
rect 9873 9877 9907 9911
rect 10609 9877 10643 9911
rect 12265 9877 12299 9911
rect 12633 9877 12667 9911
rect 14473 9877 14507 9911
rect 3709 9673 3743 9707
rect 6561 9673 6595 9707
rect 6745 9673 6779 9707
rect 6377 9605 6411 9639
rect 8125 9605 8159 9639
rect 9413 9605 9447 9639
rect 9873 9605 9907 9639
rect 12633 9605 12667 9639
rect 13921 9605 13955 9639
rect 2973 9537 3007 9571
rect 3157 9537 3191 9571
rect 3525 9537 3559 9571
rect 3801 9537 3835 9571
rect 4353 9537 4387 9571
rect 4445 9537 4479 9571
rect 6653 9537 6687 9571
rect 7481 9537 7515 9571
rect 7573 9537 7607 9571
rect 7665 9537 7699 9571
rect 9045 9537 9079 9571
rect 9137 9537 9171 9571
rect 9229 9537 9263 9571
rect 9597 9537 9631 9571
rect 11529 9537 11563 9571
rect 11989 9537 12023 9571
rect 12547 9537 12581 9571
rect 12725 9537 12759 9571
rect 14381 9537 14415 9571
rect 2329 9469 2363 9503
rect 2697 9469 2731 9503
rect 4708 9469 4742 9503
rect 7389 9469 7423 9503
rect 7849 9469 7883 9503
rect 11621 9469 11655 9503
rect 2421 9401 2455 9435
rect 2881 9401 2915 9435
rect 11345 9401 11379 9435
rect 2789 9333 2823 9367
rect 3341 9333 3375 9367
rect 4169 9333 4203 9367
rect 6193 9333 6227 9367
rect 6929 9333 6963 9367
rect 8861 9333 8895 9367
rect 12449 9333 12483 9367
rect 13001 9333 13035 9367
rect 13461 9333 13495 9367
rect 5917 9129 5951 9163
rect 13001 9129 13035 9163
rect 2421 9061 2455 9095
rect 9321 9061 9355 9095
rect 11713 9061 11747 9095
rect 5457 8993 5491 9027
rect 5733 8993 5767 9027
rect 2237 8925 2271 8959
rect 5825 8925 5859 8959
rect 6377 8925 6411 8959
rect 9137 8925 9171 8959
rect 9413 8925 9447 8959
rect 11621 8925 11655 8959
rect 11805 8925 11839 8959
rect 13185 8925 13219 8959
rect 13369 8925 13403 8959
rect 13645 8925 13679 8959
rect 7021 8857 7055 8891
rect 9689 8857 9723 8891
rect 3433 8789 3467 8823
rect 3985 8789 4019 8823
rect 8309 8789 8343 8823
rect 11161 8789 11195 8823
rect 13277 8789 13311 8823
rect 14473 8789 14507 8823
rect 11253 8585 11287 8619
rect 12081 8585 12115 8619
rect 13921 8585 13955 8619
rect 14105 8585 14139 8619
rect 14257 8517 14291 8551
rect 14473 8517 14507 8551
rect 5733 8449 5767 8483
rect 6653 8449 6687 8483
rect 8677 8449 8711 8483
rect 10517 8449 10551 8483
rect 10701 8449 10735 8483
rect 11529 8449 11563 8483
rect 12265 8449 12299 8483
rect 14013 8449 14047 8483
rect 3525 8381 3559 8415
rect 3801 8381 3835 8415
rect 5641 8381 5675 8415
rect 8953 8381 8987 8415
rect 10425 8381 10459 8415
rect 11805 8381 11839 8415
rect 13369 8381 13403 8415
rect 5273 8313 5307 8347
rect 6469 8313 6503 8347
rect 10885 8313 10919 8347
rect 3433 8245 3467 8279
rect 6101 8245 6135 8279
rect 13737 8245 13771 8279
rect 14289 8245 14323 8279
rect 4537 8041 4571 8075
rect 6929 8041 6963 8075
rect 10701 8041 10735 8075
rect 11069 8041 11103 8075
rect 10885 7973 10919 8007
rect 5457 7905 5491 7939
rect 6285 7905 6319 7939
rect 2237 7837 2271 7871
rect 2421 7837 2455 7871
rect 3893 7837 3927 7871
rect 4077 7837 4111 7871
rect 4169 7837 4203 7871
rect 4351 7837 4385 7871
rect 4813 7837 4847 7871
rect 5089 7837 5123 7871
rect 5273 7837 5307 7871
rect 5549 7837 5583 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 11437 7837 11471 7871
rect 12081 7837 12115 7871
rect 14289 7837 14323 7871
rect 3249 7769 3283 7803
rect 3617 7769 3651 7803
rect 4629 7769 4663 7803
rect 4997 7769 5031 7803
rect 2329 7701 2363 7735
rect 3985 7701 4019 7735
rect 5273 7701 5307 7735
rect 7205 7701 7239 7735
rect 11069 7701 11103 7735
rect 11713 7701 11747 7735
rect 13829 7701 13863 7735
rect 14473 7701 14507 7735
rect 2421 7497 2455 7531
rect 6745 7497 6779 7531
rect 6837 7497 6871 7531
rect 7297 7497 7331 7531
rect 10057 7497 10091 7531
rect 13461 7497 13495 7531
rect 14381 7497 14415 7531
rect 3893 7429 3927 7463
rect 4537 7429 4571 7463
rect 7665 7429 7699 7463
rect 10333 7429 10367 7463
rect 10517 7429 10551 7463
rect 10793 7429 10827 7463
rect 11805 7429 11839 7463
rect 1409 7361 1443 7395
rect 1593 7361 1627 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 8033 7361 8067 7395
rect 10241 7361 10275 7395
rect 11161 7361 11195 7395
rect 11345 7361 11379 7395
rect 13553 7361 13587 7395
rect 14013 7361 14047 7395
rect 14289 7361 14323 7395
rect 4169 7293 4203 7327
rect 4261 7293 4295 7327
rect 7113 7293 7147 7327
rect 11529 7293 11563 7327
rect 6929 7225 6963 7259
rect 7941 7225 7975 7259
rect 13277 7225 13311 7259
rect 13921 7225 13955 7259
rect 1501 7157 1535 7191
rect 6009 7157 6043 7191
rect 10241 7157 10275 7191
rect 11253 7157 11287 7191
rect 14197 7157 14231 7191
rect 2881 6953 2915 6987
rect 5089 6953 5123 6987
rect 11437 6953 11471 6987
rect 12436 6953 12470 6987
rect 3065 6817 3099 6851
rect 4721 6817 4755 6851
rect 9137 6817 9171 6851
rect 13921 6817 13955 6851
rect 2973 6749 3007 6783
rect 3801 6749 3835 6783
rect 4169 6749 4203 6783
rect 4286 6749 4320 6783
rect 4629 6749 4663 6783
rect 5273 6749 5307 6783
rect 5733 6749 5767 6783
rect 5917 6749 5951 6783
rect 6193 6749 6227 6783
rect 9229 6749 9263 6783
rect 12173 6749 12207 6783
rect 14105 6749 14139 6783
rect 7757 6681 7791 6715
rect 10149 6681 10183 6715
rect 3617 6613 3651 6647
rect 4077 6613 4111 6647
rect 4445 6613 4479 6647
rect 5457 6613 5491 6647
rect 5549 6613 5583 6647
rect 9597 6613 9631 6647
rect 14197 6613 14231 6647
rect 3525 6409 3559 6443
rect 6025 6409 6059 6443
rect 11989 6409 12023 6443
rect 5089 6341 5123 6375
rect 5825 6341 5859 6375
rect 7573 6341 7607 6375
rect 8769 6341 8803 6375
rect 10241 6341 10275 6375
rect 10701 6341 10735 6375
rect 14289 6341 14323 6375
rect 4353 6273 4387 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 6469 6273 6503 6307
rect 6745 6273 6779 6307
rect 6929 6273 6963 6307
rect 7297 6273 7331 6307
rect 10333 6273 10367 6307
rect 10793 6273 10827 6307
rect 11345 6273 11379 6307
rect 11805 6273 11839 6307
rect 12265 6273 12299 6307
rect 4813 6205 4847 6239
rect 7205 6205 7239 6239
rect 7757 6205 7791 6239
rect 8493 6205 8527 6239
rect 11621 6205 11655 6239
rect 12541 6205 12575 6239
rect 6193 6137 6227 6171
rect 10517 6137 10551 6171
rect 5365 6069 5399 6103
rect 6009 6069 6043 6103
rect 6561 6069 6595 6103
rect 8033 6069 8067 6103
rect 11161 6069 11195 6103
rect 2789 5865 2823 5899
rect 3985 5865 4019 5899
rect 4169 5865 4203 5899
rect 4537 5865 4571 5899
rect 7297 5865 7331 5899
rect 9229 5865 9263 5899
rect 10885 5865 10919 5899
rect 14289 5865 14323 5899
rect 1869 5797 1903 5831
rect 4353 5797 4387 5831
rect 4997 5797 5031 5831
rect 7757 5797 7791 5831
rect 8401 5797 8435 5831
rect 14105 5797 14139 5831
rect 3341 5729 3375 5763
rect 5273 5729 5307 5763
rect 11897 5729 11931 5763
rect 12173 5729 12207 5763
rect 13921 5729 13955 5763
rect 1685 5661 1719 5695
rect 2973 5661 3007 5695
rect 3065 5661 3099 5695
rect 4445 5661 4479 5695
rect 4629 5661 4663 5695
rect 4905 5661 4939 5695
rect 5089 5661 5123 5695
rect 7389 5661 7423 5695
rect 8033 5661 8067 5695
rect 8309 5661 8343 5695
rect 8401 5661 8435 5695
rect 8677 5661 8711 5695
rect 11621 5661 11655 5695
rect 11805 5661 11839 5695
rect 2237 5593 2271 5627
rect 3801 5593 3835 5627
rect 4813 5593 4847 5627
rect 5549 5593 5583 5627
rect 7757 5593 7791 5627
rect 8125 5593 8159 5627
rect 14257 5593 14291 5627
rect 14473 5593 14507 5627
rect 3157 5525 3191 5559
rect 4011 5525 4045 5559
rect 7021 5525 7055 5559
rect 7941 5525 7975 5559
rect 9505 5525 9539 5559
rect 11437 5525 11471 5559
rect 11621 5525 11655 5559
rect 3249 5321 3283 5355
rect 3617 5321 3651 5355
rect 4353 5321 4387 5355
rect 5473 5321 5507 5355
rect 5089 5253 5123 5287
rect 5273 5253 5307 5287
rect 5825 5253 5859 5287
rect 6041 5253 6075 5287
rect 6745 5253 6779 5287
rect 11805 5253 11839 5287
rect 11989 5253 12023 5287
rect 12725 5253 12759 5287
rect 14473 5253 14507 5287
rect 6561 5185 6595 5219
rect 8769 5185 8803 5219
rect 9321 5185 9355 5219
rect 9505 5185 9539 5219
rect 9597 5185 9631 5219
rect 12449 5185 12483 5219
rect 4813 5117 4847 5151
rect 6377 5117 6411 5151
rect 8493 5117 8527 5151
rect 9873 5117 9907 5151
rect 11345 5117 11379 5151
rect 5641 5049 5675 5083
rect 6193 5049 6227 5083
rect 7021 5049 7055 5083
rect 5457 4981 5491 5015
rect 6009 4981 6043 5015
rect 9137 4981 9171 5015
rect 9321 4981 9355 5015
rect 11621 4981 11655 5015
rect 11805 4981 11839 5015
rect 12265 4981 12299 5015
rect 1961 4777 1995 4811
rect 3525 4777 3559 4811
rect 7849 4777 7883 4811
rect 8033 4777 8067 4811
rect 8401 4777 8435 4811
rect 9965 4777 9999 4811
rect 11161 4777 11195 4811
rect 13645 4777 13679 4811
rect 14473 4777 14507 4811
rect 2329 4709 2363 4743
rect 2881 4709 2915 4743
rect 5365 4709 5399 4743
rect 8953 4709 8987 4743
rect 7573 4641 7607 4675
rect 12357 4641 12391 4675
rect 1777 4573 1811 4607
rect 1961 4573 1995 4607
rect 2145 4573 2179 4607
rect 2329 4573 2363 4607
rect 2697 4573 2731 4607
rect 3249 4573 3283 4607
rect 3617 4573 3651 4607
rect 5181 4573 5215 4607
rect 5825 4573 5859 4607
rect 8309 4573 8343 4607
rect 9229 4573 9263 4607
rect 9321 4573 9355 4607
rect 9413 4573 9447 4607
rect 9597 4573 9631 4607
rect 11575 4573 11609 4607
rect 11713 4573 11747 4607
rect 11805 4573 11839 4607
rect 11989 4573 12023 4607
rect 12541 4573 12575 4607
rect 12633 4573 12667 4607
rect 13737 4573 13771 4607
rect 14289 4573 14323 4607
rect 6101 4505 6135 4539
rect 8217 4505 8251 4539
rect 10793 4505 10827 4539
rect 10977 4505 11011 4539
rect 11345 4505 11379 4539
rect 1685 4437 1719 4471
rect 3065 4437 3099 4471
rect 4077 4437 4111 4471
rect 5733 4437 5767 4471
rect 8017 4437 8051 4471
rect 10609 4437 10643 4471
rect 13093 4437 13127 4471
rect 13921 4437 13955 4471
rect 2973 4233 3007 4267
rect 3433 4233 3467 4267
rect 13921 4233 13955 4267
rect 8401 4165 8435 4199
rect 12817 4165 12851 4199
rect 2513 4097 2547 4131
rect 6929 4097 6963 4131
rect 11805 4097 11839 4131
rect 11989 4097 12023 4131
rect 13737 4097 13771 4131
rect 14013 4097 14047 4131
rect 14289 4097 14323 4131
rect 14381 4097 14415 4131
rect 6101 4029 6135 4063
rect 7021 4029 7055 4063
rect 9137 4029 9171 4063
rect 12173 4029 12207 4063
rect 13185 4029 13219 4063
rect 2697 3961 2731 3995
rect 5733 3961 5767 3995
rect 6561 3961 6595 3995
rect 7757 3961 7791 3995
rect 11253 3961 11287 3995
rect 13461 3961 13495 3995
rect 14105 3961 14139 3995
rect 8769 3893 8803 3927
rect 1501 3689 1535 3723
rect 2513 3689 2547 3723
rect 6837 3689 6871 3723
rect 7665 3689 7699 3723
rect 9505 3689 9539 3723
rect 10057 3689 10091 3723
rect 11713 3689 11747 3723
rect 13737 3689 13771 3723
rect 14289 3689 14323 3723
rect 8585 3621 8619 3655
rect 9689 3621 9723 3655
rect 14105 3621 14139 3655
rect 9137 3553 9171 3587
rect 1501 3485 1535 3519
rect 1777 3485 1811 3519
rect 6929 3485 6963 3519
rect 7021 3485 7055 3519
rect 7113 3485 7147 3519
rect 7297 3485 7331 3519
rect 8033 3485 8067 3519
rect 8217 3485 8251 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 13001 3485 13035 3519
rect 13093 3485 13127 3519
rect 6745 3417 6779 3451
rect 9321 3417 9355 3451
rect 9537 3417 9571 3451
rect 11437 3417 11471 3451
rect 11897 3417 11931 3451
rect 14473 3417 14507 3451
rect 1685 3349 1719 3383
rect 2145 3349 2179 3383
rect 11529 3349 11563 3383
rect 11697 3349 11731 3383
rect 12449 3349 12483 3383
rect 12817 3349 12851 3383
rect 14273 3349 14307 3383
rect 3157 3145 3191 3179
rect 3801 3145 3835 3179
rect 7849 3145 7883 3179
rect 8861 3145 8895 3179
rect 9505 3145 9539 3179
rect 9873 3145 9907 3179
rect 10609 3145 10643 3179
rect 11897 3145 11931 3179
rect 3433 3077 3467 3111
rect 8677 3077 8711 3111
rect 12265 3077 12299 3111
rect 14289 3077 14323 3111
rect 3157 3009 3191 3043
rect 3249 3009 3283 3043
rect 8953 3009 8987 3043
rect 9045 3009 9079 3043
rect 10149 3009 10183 3043
rect 10424 3009 10458 3043
rect 10885 3009 10919 3043
rect 11989 3009 12023 3043
rect 13829 3009 13863 3043
rect 14013 3009 14047 3043
rect 14197 3009 14231 3043
rect 10241 2941 10275 2975
rect 10333 2941 10367 2975
rect 11253 2941 11287 2975
rect 8677 2873 8711 2907
rect 9137 2873 9171 2907
rect 14105 2873 14139 2907
rect 13737 2805 13771 2839
rect 1593 2601 1627 2635
rect 9229 2601 9263 2635
rect 12909 2601 12943 2635
rect 14289 2601 14323 2635
rect 11529 2533 11563 2567
rect 3065 2465 3099 2499
rect 3341 2465 3375 2499
rect 10701 2465 10735 2499
rect 13277 2465 13311 2499
rect 9045 2397 9079 2431
rect 9137 2397 9171 2431
rect 9413 2397 9447 2431
rect 11069 2397 11103 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 13461 2397 13495 2431
rect 13737 2397 13771 2431
rect 14473 2397 14507 2431
rect 8769 2329 8803 2363
rect 9505 2329 9539 2363
rect 9781 2329 9815 2363
rect 10885 2329 10919 2363
rect 10977 2329 11011 2363
rect 9597 2261 9631 2295
rect 10149 2261 10183 2295
rect 11253 2261 11287 2295
rect 12541 2261 12575 2295
rect 13645 2261 13679 2295
rect 13921 2261 13955 2295
<< metal1 >>
rect 6638 15920 6644 15972
rect 6696 15960 6702 15972
rect 14734 15960 14740 15972
rect 6696 15932 14740 15960
rect 6696 15920 6702 15932
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 658 15852 664 15904
rect 716 15892 722 15904
rect 9674 15892 9680 15904
rect 716 15864 9680 15892
rect 716 15852 722 15864
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 1104 15802 14812 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 14812 15802
rect 1104 15728 14812 15750
rect 9585 15691 9643 15697
rect 9585 15657 9597 15691
rect 9631 15688 9643 15691
rect 14550 15688 14556 15700
rect 9631 15660 14556 15688
rect 9631 15657 9643 15660
rect 9585 15651 9643 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 10505 15623 10563 15629
rect 10505 15589 10517 15623
rect 10551 15620 10563 15623
rect 14366 15620 14372 15632
rect 10551 15592 14372 15620
rect 10551 15589 10563 15592
rect 10505 15583 10563 15589
rect 14366 15580 14372 15592
rect 14424 15580 14430 15632
rect 8202 15552 8208 15564
rect 4080 15524 8208 15552
rect 4080 15493 4108 15524
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15552 8355 15555
rect 10594 15552 10600 15564
rect 8343 15524 10600 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 13081 15555 13139 15561
rect 13081 15521 13093 15555
rect 13127 15552 13139 15555
rect 13722 15552 13728 15564
rect 13127 15524 13728 15552
rect 13127 15521 13139 15524
rect 13081 15515 13139 15521
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 14182 15512 14188 15564
rect 14240 15512 14246 15564
rect 4065 15487 4123 15493
rect 4065 15453 4077 15487
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15484 4307 15487
rect 4525 15487 4583 15493
rect 4525 15484 4537 15487
rect 4295 15456 4537 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 4525 15453 4537 15456
rect 4571 15484 4583 15487
rect 4890 15484 4896 15496
rect 4571 15456 4896 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15484 8631 15487
rect 8938 15484 8944 15496
rect 8619 15456 8944 15484
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 9180 15456 9505 15484
rect 9180 15444 9186 15456
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 10318 15444 10324 15496
rect 10376 15444 10382 15496
rect 12728 15456 13308 15484
rect 5994 15376 6000 15428
rect 6052 15416 6058 15428
rect 6052 15388 7130 15416
rect 6052 15376 6058 15388
rect 10134 15376 10140 15428
rect 10192 15416 10198 15428
rect 12728 15425 12756 15456
rect 12529 15419 12587 15425
rect 12529 15416 12541 15419
rect 10192 15388 12541 15416
rect 10192 15376 10198 15388
rect 12529 15385 12541 15388
rect 12575 15385 12587 15419
rect 12529 15379 12587 15385
rect 12713 15419 12771 15425
rect 12713 15385 12725 15419
rect 12759 15385 12771 15419
rect 12713 15379 12771 15385
rect 12805 15419 12863 15425
rect 12805 15385 12817 15419
rect 12851 15416 12863 15419
rect 13280 15416 13308 15456
rect 14274 15444 14280 15496
rect 14332 15444 14338 15496
rect 15286 15416 15292 15428
rect 12851 15388 13216 15416
rect 13280 15388 15292 15416
rect 12851 15385 12863 15388
rect 12805 15379 12863 15385
rect 13188 15360 13216 15388
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 2406 15308 2412 15360
rect 2464 15308 2470 15360
rect 2777 15351 2835 15357
rect 2777 15317 2789 15351
rect 2823 15348 2835 15351
rect 3234 15348 3240 15360
rect 2823 15320 3240 15348
rect 2823 15317 2835 15320
rect 2777 15311 2835 15317
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 3881 15351 3939 15357
rect 3881 15317 3893 15351
rect 3927 15348 3939 15351
rect 5074 15348 5080 15360
rect 3927 15320 5080 15348
rect 3927 15317 3939 15320
rect 3881 15311 3939 15317
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 6822 15308 6828 15360
rect 6880 15308 6886 15360
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 12492 15320 12909 15348
rect 12492 15308 12498 15320
rect 12897 15317 12909 15320
rect 12943 15317 12955 15351
rect 12897 15311 12955 15317
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 13357 15351 13415 15357
rect 13357 15348 13369 15351
rect 13228 15320 13369 15348
rect 13228 15308 13234 15320
rect 13357 15317 13369 15320
rect 13403 15317 13415 15351
rect 13357 15311 13415 15317
rect 13906 15308 13912 15360
rect 13964 15308 13970 15360
rect 1104 15258 14812 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 14812 15258
rect 1104 15184 14812 15206
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 3878 15144 3884 15156
rect 2464 15116 3884 15144
rect 2464 15104 2470 15116
rect 3878 15104 3884 15116
rect 3936 15104 3942 15156
rect 6546 15144 6552 15156
rect 4264 15116 6552 15144
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 1596 14940 1624 14971
rect 1854 14968 1860 15020
rect 1912 14968 1918 15020
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 2424 15008 2452 15104
rect 4264 15076 4292 15116
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 6638 15104 6644 15156
rect 6696 15104 6702 15156
rect 7193 15147 7251 15153
rect 6748 15116 7144 15144
rect 3818 15048 4292 15076
rect 4338 15036 4344 15088
rect 4396 15076 4402 15088
rect 6748 15076 6776 15116
rect 4396 15048 6776 15076
rect 6825 15079 6883 15085
rect 4396 15036 4402 15048
rect 6825 15045 6837 15079
rect 6871 15076 6883 15079
rect 6914 15076 6920 15088
rect 6871 15048 6920 15076
rect 6871 15045 6883 15048
rect 6825 15039 6883 15045
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 7116 15076 7144 15116
rect 7193 15113 7205 15147
rect 7239 15144 7251 15147
rect 8110 15144 8116 15156
rect 7239 15116 8116 15144
rect 7239 15113 7251 15116
rect 7193 15107 7251 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 10965 15147 11023 15153
rect 10965 15144 10977 15147
rect 10836 15116 10977 15144
rect 10836 15104 10842 15116
rect 10965 15113 10977 15116
rect 11011 15113 11023 15147
rect 10965 15107 11023 15113
rect 14001 15147 14059 15153
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14274 15144 14280 15156
rect 14047 15116 14280 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14274 15104 14280 15116
rect 14332 15144 14338 15156
rect 14918 15144 14924 15156
rect 14332 15116 14924 15144
rect 14332 15104 14338 15116
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 7116 15048 7236 15076
rect 2087 14980 2452 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 5350 14968 5356 15020
rect 5408 15008 5414 15020
rect 5537 15011 5595 15017
rect 5537 15008 5549 15011
rect 5408 14980 5549 15008
rect 5408 14968 5414 14980
rect 5537 14977 5549 14980
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 5721 15011 5779 15017
rect 5721 14977 5733 15011
rect 5767 15008 5779 15011
rect 5902 15008 5908 15020
rect 5767 14980 5908 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 3234 14940 3240 14952
rect 1596 14912 3240 14940
rect 3234 14900 3240 14912
rect 3292 14900 3298 14952
rect 4246 14900 4252 14952
rect 4304 14900 4310 14952
rect 4522 14900 4528 14952
rect 4580 14900 4586 14952
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14872 2007 14875
rect 3142 14872 3148 14884
rect 1995 14844 3148 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 3142 14832 3148 14844
rect 3200 14832 3206 14884
rect 4540 14872 4568 14900
rect 5166 14872 5172 14884
rect 4540 14844 5172 14872
rect 5166 14832 5172 14844
rect 5224 14872 5230 14884
rect 5718 14872 5724 14884
rect 5224 14844 5724 14872
rect 5224 14832 5230 14844
rect 5718 14832 5724 14844
rect 5776 14832 5782 14884
rect 7024 14872 7052 14971
rect 7098 14968 7104 15020
rect 7156 14968 7162 15020
rect 7208 15008 7236 15048
rect 7282 15036 7288 15088
rect 7340 15076 7346 15088
rect 10686 15076 10692 15088
rect 7340 15048 10692 15076
rect 7340 15036 7346 15048
rect 10686 15036 10692 15048
rect 10744 15036 10750 15088
rect 10870 15036 10876 15088
rect 10928 15076 10934 15088
rect 12253 15079 12311 15085
rect 12253 15076 12265 15079
rect 10928 15048 11100 15076
rect 10928 15036 10934 15048
rect 10502 15008 10508 15020
rect 7208 14980 10508 15008
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 15008 10839 15011
rect 10962 15008 10968 15020
rect 10827 14980 10968 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 11072 15017 11100 15048
rect 11716 15048 12265 15076
rect 11716 15020 11744 15048
rect 12253 15045 12265 15048
rect 12299 15045 12311 15079
rect 12253 15039 12311 15045
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 14977 11115 15011
rect 11057 14971 11115 14977
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 14977 12035 15011
rect 11977 14971 12035 14977
rect 8478 14900 8484 14952
rect 8536 14940 8542 14952
rect 11992 14940 12020 14971
rect 14458 14968 14464 15020
rect 14516 14968 14522 15020
rect 8536 14912 12020 14940
rect 8536 14900 8542 14912
rect 7024 14844 10916 14872
rect 1486 14764 1492 14816
rect 1544 14804 1550 14816
rect 1854 14804 1860 14816
rect 1544 14776 1860 14804
rect 1544 14764 1550 14776
rect 1854 14764 1860 14776
rect 1912 14804 1918 14816
rect 2501 14807 2559 14813
rect 2501 14804 2513 14807
rect 1912 14776 2513 14804
rect 1912 14764 1918 14776
rect 2501 14773 2513 14776
rect 2547 14773 2559 14807
rect 2501 14767 2559 14773
rect 2777 14807 2835 14813
rect 2777 14773 2789 14807
rect 2823 14804 2835 14807
rect 3234 14804 3240 14816
rect 2823 14776 3240 14804
rect 2823 14773 2835 14776
rect 2777 14767 2835 14773
rect 3234 14764 3240 14776
rect 3292 14764 3298 14816
rect 5350 14764 5356 14816
rect 5408 14764 5414 14816
rect 5626 14764 5632 14816
rect 5684 14764 5690 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7653 14807 7711 14813
rect 7653 14804 7665 14807
rect 7156 14776 7665 14804
rect 7156 14764 7162 14776
rect 7653 14773 7665 14776
rect 7699 14804 7711 14807
rect 8386 14804 8392 14816
rect 7699 14776 8392 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 8386 14764 8392 14776
rect 8444 14764 8450 14816
rect 10318 14764 10324 14816
rect 10376 14764 10382 14816
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 10781 14807 10839 14813
rect 10781 14804 10793 14807
rect 10468 14776 10793 14804
rect 10468 14764 10474 14776
rect 10781 14773 10793 14776
rect 10827 14773 10839 14807
rect 10888 14804 10916 14844
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 11793 14875 11851 14881
rect 11793 14872 11805 14875
rect 11112 14844 11805 14872
rect 11112 14832 11118 14844
rect 11793 14841 11805 14844
rect 11839 14841 11851 14875
rect 11793 14835 11851 14841
rect 12342 14832 12348 14884
rect 12400 14872 12406 14884
rect 12526 14872 12532 14884
rect 12400 14844 12532 14872
rect 12400 14832 12406 14844
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 11514 14804 11520 14816
rect 10888 14776 11520 14804
rect 10781 14767 10839 14773
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 11606 14764 11612 14816
rect 11664 14764 11670 14816
rect 1104 14714 14812 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 14812 14714
rect 1104 14640 14812 14662
rect 1578 14560 1584 14612
rect 1636 14560 1642 14612
rect 4706 14600 4712 14612
rect 1688 14572 4712 14600
rect 934 14492 940 14544
rect 992 14532 998 14544
rect 1688 14532 1716 14572
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5316 14572 5672 14600
rect 5316 14560 5322 14572
rect 2961 14535 3019 14541
rect 2961 14532 2973 14535
rect 992 14504 1716 14532
rect 2746 14504 2973 14532
rect 992 14492 998 14504
rect 1946 14424 1952 14476
rect 2004 14464 2010 14476
rect 2746 14464 2774 14504
rect 2961 14501 2973 14504
rect 3007 14532 3019 14535
rect 4338 14532 4344 14544
rect 3007 14504 4344 14532
rect 3007 14501 3019 14504
rect 2961 14495 3019 14501
rect 4338 14492 4344 14504
rect 4396 14492 4402 14544
rect 5644 14532 5672 14572
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 10778 14600 10784 14612
rect 7524 14572 10784 14600
rect 7524 14560 7530 14572
rect 10778 14560 10784 14572
rect 10836 14600 10842 14612
rect 10965 14603 11023 14609
rect 10965 14600 10977 14603
rect 10836 14572 10977 14600
rect 10836 14560 10842 14572
rect 10965 14569 10977 14572
rect 11011 14569 11023 14603
rect 10965 14563 11023 14569
rect 8294 14532 8300 14544
rect 5644 14504 8300 14532
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 12342 14532 12348 14544
rect 10244 14504 12348 14532
rect 2004 14436 2774 14464
rect 2004 14424 2010 14436
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 5445 14467 5503 14473
rect 5445 14464 5457 14467
rect 3844 14436 5457 14464
rect 3844 14424 3850 14436
rect 5445 14433 5457 14436
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 5718 14424 5724 14476
rect 5776 14424 5782 14476
rect 10244 14464 10272 14504
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 5828 14436 10272 14464
rect 12406 14436 12817 14464
rect 2041 14399 2099 14405
rect 2041 14396 2053 14399
rect 1412 14368 2053 14396
rect 1412 14337 1440 14368
rect 2041 14365 2053 14368
rect 2087 14396 2099 14399
rect 4154 14396 4160 14408
rect 2087 14368 4160 14396
rect 2087 14365 2099 14368
rect 2041 14359 2099 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 1397 14331 1455 14337
rect 1397 14297 1409 14331
rect 1443 14297 1455 14331
rect 1397 14291 1455 14297
rect 1613 14331 1671 14337
rect 1613 14297 1625 14331
rect 1659 14328 1671 14331
rect 1854 14328 1860 14340
rect 1659 14300 1860 14328
rect 1659 14297 1671 14300
rect 1613 14291 1671 14297
rect 1854 14288 1860 14300
rect 1912 14288 1918 14340
rect 5014 14300 5396 14328
rect 1762 14220 1768 14272
rect 1820 14220 1826 14272
rect 2593 14263 2651 14269
rect 2593 14229 2605 14263
rect 2639 14260 2651 14263
rect 2958 14260 2964 14272
rect 2639 14232 2964 14260
rect 2639 14229 2651 14232
rect 2593 14223 2651 14229
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 3973 14263 4031 14269
rect 3973 14229 3985 14263
rect 4019 14260 4031 14263
rect 4430 14260 4436 14272
rect 4019 14232 4436 14260
rect 4019 14229 4031 14232
rect 3973 14223 4031 14229
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 4614 14220 4620 14272
rect 4672 14260 4678 14272
rect 5258 14260 5264 14272
rect 4672 14232 5264 14260
rect 4672 14220 4678 14232
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5368 14260 5396 14300
rect 5828 14260 5856 14436
rect 12406 14408 12434 14436
rect 12805 14433 12817 14436
rect 12851 14464 12863 14467
rect 13262 14464 13268 14476
rect 12851 14436 13268 14464
rect 12851 14433 12863 14436
rect 12805 14427 12863 14433
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 6546 14356 6552 14408
rect 6604 14396 6610 14408
rect 8754 14396 8760 14408
rect 6604 14368 8760 14396
rect 6604 14356 6610 14368
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 8938 14356 8944 14408
rect 8996 14356 9002 14408
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 11333 14399 11391 14405
rect 11333 14396 11345 14399
rect 11020 14368 11345 14396
rect 11020 14356 11026 14368
rect 11333 14365 11345 14368
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 12342 14356 12348 14408
rect 12400 14368 12434 14408
rect 12400 14356 12406 14368
rect 9214 14288 9220 14340
rect 9272 14288 9278 14340
rect 13906 14328 13912 14340
rect 10442 14300 13912 14328
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 5368 14232 5856 14260
rect 6086 14220 6092 14272
rect 6144 14260 6150 14272
rect 9858 14260 9864 14272
rect 6144 14232 9864 14260
rect 6144 14220 6150 14232
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 9950 14220 9956 14272
rect 10008 14260 10014 14272
rect 10689 14263 10747 14269
rect 10689 14260 10701 14263
rect 10008 14232 10701 14260
rect 10008 14220 10014 14232
rect 10689 14229 10701 14232
rect 10735 14229 10747 14263
rect 10689 14223 10747 14229
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 11701 14263 11759 14269
rect 11701 14260 11713 14263
rect 10928 14232 11713 14260
rect 10928 14220 10934 14232
rect 11701 14229 11713 14232
rect 11747 14229 11759 14263
rect 11701 14223 11759 14229
rect 13265 14263 13323 14269
rect 13265 14229 13277 14263
rect 13311 14260 13323 14263
rect 13538 14260 13544 14272
rect 13311 14232 13544 14260
rect 13311 14229 13323 14232
rect 13265 14223 13323 14229
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 13814 14220 13820 14272
rect 13872 14220 13878 14272
rect 14458 14220 14464 14272
rect 14516 14220 14522 14272
rect 1104 14170 14812 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 14812 14170
rect 1104 14096 14812 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1627 14028 4016 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 2041 13991 2099 13997
rect 2041 13957 2053 13991
rect 2087 13988 2099 13991
rect 2774 13988 2780 14000
rect 2087 13960 2780 13988
rect 2087 13957 2099 13960
rect 2041 13951 2099 13957
rect 2774 13948 2780 13960
rect 2832 13948 2838 14000
rect 3602 13948 3608 14000
rect 3660 13948 3666 14000
rect 3988 13988 4016 14028
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 6822 14056 6828 14068
rect 4212 14028 6828 14056
rect 4212 14016 4218 14028
rect 6822 14016 6828 14028
rect 6880 14056 6886 14068
rect 6880 14028 8294 14056
rect 6880 14016 6886 14028
rect 4614 13988 4620 14000
rect 3988 13960 4620 13988
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 4798 13948 4804 14000
rect 4856 13988 4862 14000
rect 8113 13991 8171 13997
rect 8113 13988 8125 13991
rect 4856 13960 8125 13988
rect 4856 13948 4862 13960
rect 8113 13957 8125 13960
rect 8159 13957 8171 13991
rect 8113 13951 8171 13957
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 1946 13880 1952 13932
rect 2004 13880 2010 13932
rect 2222 13880 2228 13932
rect 2280 13880 2286 13932
rect 4338 13880 4344 13932
rect 4396 13880 4402 13932
rect 4522 13880 4528 13932
rect 4580 13880 4586 13932
rect 4706 13880 4712 13932
rect 4764 13880 4770 13932
rect 5718 13880 5724 13932
rect 5776 13920 5782 13932
rect 5905 13923 5963 13929
rect 5905 13920 5917 13923
rect 5776 13892 5917 13920
rect 5776 13880 5782 13892
rect 5905 13889 5917 13892
rect 5951 13920 5963 13923
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 5951 13892 6561 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 8266 13920 8294 14028
rect 8478 14016 8484 14068
rect 8536 14016 8542 14068
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 11330 14056 11336 14068
rect 9539 14028 11336 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 12584 14028 12633 14056
rect 12584 14016 12590 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 12621 14019 12679 14025
rect 8329 13991 8387 13997
rect 8329 13957 8341 13991
rect 8375 13988 8387 13991
rect 9030 13988 9036 14000
rect 8375 13960 9036 13988
rect 8375 13957 8387 13960
rect 8329 13951 8387 13957
rect 9030 13948 9036 13960
rect 9088 13948 9094 14000
rect 9125 13991 9183 13997
rect 9125 13957 9137 13991
rect 9171 13957 9183 13991
rect 9125 13951 9183 13957
rect 9341 13991 9399 13997
rect 9341 13957 9353 13991
rect 9387 13988 9399 13991
rect 9582 13988 9588 14000
rect 9387 13960 9588 13988
rect 9387 13957 9399 13960
rect 9341 13951 9399 13957
rect 8941 13923 8999 13929
rect 8941 13920 8953 13923
rect 8266 13892 8953 13920
rect 6549 13883 6607 13889
rect 8941 13889 8953 13892
rect 8987 13920 8999 13923
rect 9140 13920 9168 13951
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 9674 13948 9680 14000
rect 9732 13988 9738 14000
rect 12989 13991 13047 13997
rect 12989 13988 13001 13991
rect 9732 13960 13001 13988
rect 9732 13948 9738 13960
rect 12989 13957 13001 13960
rect 13035 13957 13047 13991
rect 13538 13988 13544 14000
rect 12989 13951 13047 13957
rect 13096 13960 13544 13988
rect 8987 13892 9168 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 11701 13923 11759 13929
rect 11701 13920 11713 13923
rect 9916 13892 11713 13920
rect 9916 13880 9922 13892
rect 11701 13889 11713 13892
rect 11747 13920 11759 13923
rect 12342 13920 12348 13932
rect 11747 13892 12348 13920
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13920 12771 13923
rect 13096 13920 13124 13960
rect 13538 13948 13544 13960
rect 13596 13948 13602 14000
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 13998 13988 14004 14000
rect 13872 13960 14004 13988
rect 13872 13948 13878 13960
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 12759 13892 13124 13920
rect 13173 13923 13231 13929
rect 12759 13889 12771 13892
rect 12713 13883 12771 13889
rect 13173 13889 13185 13923
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 1762 13812 1768 13864
rect 1820 13852 1826 13864
rect 2317 13855 2375 13861
rect 1820 13824 2268 13852
rect 1820 13812 1826 13824
rect 2240 13793 2268 13824
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 3510 13852 3516 13864
rect 2363 13824 3516 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 4724 13793 4752 13880
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 6730 13852 6736 13864
rect 5408 13824 6736 13852
rect 5408 13812 5414 13824
rect 6730 13812 6736 13824
rect 6788 13852 6794 13864
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 6788 13824 7113 13852
rect 6788 13812 6794 13824
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 9306 13852 9312 13864
rect 8352 13824 9312 13852
rect 8352 13812 8358 13824
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 13188 13852 13216 13883
rect 13262 13880 13268 13932
rect 13320 13880 13326 13932
rect 13446 13880 13452 13932
rect 13504 13880 13510 13932
rect 14182 13880 14188 13932
rect 14240 13880 14246 13932
rect 12360 13824 13216 13852
rect 2225 13787 2283 13793
rect 2225 13753 2237 13787
rect 2271 13753 2283 13787
rect 2225 13747 2283 13753
rect 4709 13787 4767 13793
rect 4709 13753 4721 13787
rect 4755 13753 4767 13787
rect 4709 13747 4767 13753
rect 5994 13744 6000 13796
rect 6052 13744 6058 13796
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 8076 13756 9352 13784
rect 8076 13744 8082 13756
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 2130 13716 2136 13728
rect 1728 13688 2136 13716
rect 1728 13676 1734 13688
rect 2130 13676 2136 13688
rect 2188 13676 2194 13728
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4077 13719 4135 13725
rect 4077 13716 4089 13719
rect 4028 13688 4089 13716
rect 4028 13676 4034 13688
rect 4077 13685 4089 13688
rect 4123 13685 4135 13719
rect 4077 13679 4135 13685
rect 4614 13676 4620 13728
rect 4672 13716 4678 13728
rect 4985 13719 5043 13725
rect 4985 13716 4997 13719
rect 4672 13688 4997 13716
rect 4672 13676 4678 13688
rect 4985 13685 4997 13688
rect 5031 13716 5043 13719
rect 5350 13716 5356 13728
rect 5031 13688 5356 13716
rect 5031 13685 5043 13688
rect 4985 13679 5043 13685
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 5442 13676 5448 13728
rect 5500 13716 5506 13728
rect 7558 13716 7564 13728
rect 5500 13688 7564 13716
rect 5500 13676 5506 13688
rect 7558 13676 7564 13688
rect 7616 13676 7622 13728
rect 8294 13676 8300 13728
rect 8352 13676 8358 13728
rect 9324 13725 9352 13756
rect 9309 13719 9367 13725
rect 9309 13685 9321 13719
rect 9355 13685 9367 13719
rect 9309 13679 9367 13685
rect 9398 13676 9404 13728
rect 9456 13716 9462 13728
rect 11146 13716 11152 13728
rect 9456 13688 11152 13716
rect 9456 13676 9462 13688
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 12360 13725 12388 13824
rect 13354 13812 13360 13864
rect 13412 13812 13418 13864
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 15654 13852 15660 13864
rect 14415 13824 15660 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 12345 13719 12403 13725
rect 12345 13716 12357 13719
rect 11848 13688 12357 13716
rect 11848 13676 11854 13688
rect 12345 13685 12357 13688
rect 12391 13685 12403 13719
rect 12345 13679 12403 13685
rect 13538 13676 13544 13728
rect 13596 13716 13602 13728
rect 13909 13719 13967 13725
rect 13909 13716 13921 13719
rect 13596 13688 13921 13716
rect 13596 13676 13602 13688
rect 13909 13685 13921 13688
rect 13955 13716 13967 13719
rect 14090 13716 14096 13728
rect 13955 13688 14096 13716
rect 13955 13685 13967 13688
rect 13909 13679 13967 13685
rect 14090 13676 14096 13688
rect 14148 13676 14154 13728
rect 1104 13626 14812 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 14812 13626
rect 1104 13552 14812 13574
rect 4062 13472 4068 13524
rect 4120 13472 4126 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 4614 13512 4620 13524
rect 4571 13484 4620 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 4709 13515 4767 13521
rect 4709 13481 4721 13515
rect 4755 13512 4767 13515
rect 6454 13512 6460 13524
rect 4755 13484 6460 13512
rect 4755 13481 4767 13484
rect 4709 13475 4767 13481
rect 6454 13472 6460 13484
rect 6512 13472 6518 13524
rect 7116 13484 8984 13512
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 5534 13444 5540 13456
rect 2363 13416 5540 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 2332 13308 2360 13407
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 3510 13336 3516 13388
rect 3568 13376 3574 13388
rect 3973 13379 4031 13385
rect 3973 13376 3985 13379
rect 3568 13348 3985 13376
rect 3568 13336 3574 13348
rect 3973 13345 3985 13348
rect 4019 13345 4031 13379
rect 7116 13376 7144 13484
rect 7561 13447 7619 13453
rect 7561 13413 7573 13447
rect 7607 13444 7619 13447
rect 8110 13444 8116 13456
rect 7607 13416 8116 13444
rect 7607 13413 7619 13416
rect 7561 13407 7619 13413
rect 8110 13404 8116 13416
rect 8168 13404 8174 13456
rect 8202 13404 8208 13456
rect 8260 13444 8266 13456
rect 8478 13444 8484 13456
rect 8260 13416 8484 13444
rect 8260 13404 8266 13416
rect 8478 13404 8484 13416
rect 8536 13404 8542 13456
rect 8956 13444 8984 13484
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 11885 13515 11943 13521
rect 11885 13512 11897 13515
rect 9088 13484 11897 13512
rect 9088 13472 9094 13484
rect 11885 13481 11897 13484
rect 11931 13481 11943 13515
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 11885 13475 11943 13481
rect 11992 13484 13829 13512
rect 9766 13444 9772 13456
rect 8956 13416 9772 13444
rect 9766 13404 9772 13416
rect 9824 13404 9830 13456
rect 11146 13404 11152 13456
rect 11204 13444 11210 13456
rect 11992 13444 12020 13484
rect 13817 13481 13829 13484
rect 13863 13481 13875 13515
rect 13817 13475 13875 13481
rect 11204 13416 12020 13444
rect 11204 13404 11210 13416
rect 3973 13339 4031 13345
rect 4264 13348 7144 13376
rect 7193 13379 7251 13385
rect 2777 13311 2835 13317
rect 2777 13308 2789 13311
rect 1995 13280 2360 13308
rect 2608 13280 2789 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 1118 13200 1124 13252
rect 1176 13240 1182 13252
rect 2608 13249 2636 13280
rect 2777 13277 2789 13280
rect 2823 13277 2835 13311
rect 2777 13271 2835 13277
rect 2866 13268 2872 13320
rect 2924 13308 2930 13320
rect 3602 13308 3608 13320
rect 2924 13280 3608 13308
rect 2924 13268 2930 13280
rect 3602 13268 3608 13280
rect 3660 13308 3666 13320
rect 3881 13311 3939 13317
rect 3881 13308 3893 13311
rect 3660 13280 3893 13308
rect 3660 13268 3666 13280
rect 3881 13277 3893 13280
rect 3927 13277 3939 13311
rect 3881 13271 3939 13277
rect 2593 13243 2651 13249
rect 2593 13240 2605 13243
rect 1176 13212 2605 13240
rect 1176 13200 1182 13212
rect 2593 13209 2605 13212
rect 2639 13209 2651 13243
rect 4264 13240 4292 13348
rect 7193 13345 7205 13379
rect 7239 13376 7251 13379
rect 8570 13376 8576 13388
rect 7239 13348 8576 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 8570 13336 8576 13348
rect 8628 13376 8634 13388
rect 8938 13376 8944 13388
rect 8628 13348 8944 13376
rect 8628 13336 8634 13348
rect 8938 13336 8944 13348
rect 8996 13376 9002 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 8996 13348 11069 13376
rect 8996 13336 9002 13348
rect 11057 13345 11069 13348
rect 11103 13376 11115 13379
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11103 13348 12081 13376
rect 11103 13345 11115 13348
rect 11057 13339 11115 13345
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4356 13280 5089 13308
rect 4356 13252 4384 13280
rect 5077 13277 5089 13280
rect 5123 13308 5135 13311
rect 5442 13308 5448 13320
rect 5123 13280 5448 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7616 13280 7941 13308
rect 7616 13268 7622 13280
rect 7929 13277 7941 13280
rect 7975 13308 7987 13311
rect 9398 13308 9404 13320
rect 7975 13280 9404 13308
rect 7975 13277 7987 13280
rect 7929 13271 7987 13277
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11790 13308 11796 13320
rect 11480 13280 11796 13308
rect 11480 13268 11486 13280
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 11977 13311 12035 13317
rect 11977 13277 11989 13311
rect 12023 13308 12035 13311
rect 12023 13280 12112 13308
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 2593 13203 2651 13209
rect 2976 13212 4292 13240
rect 1302 13132 1308 13184
rect 1360 13172 1366 13184
rect 2976 13181 3004 13212
rect 4338 13200 4344 13252
rect 4396 13200 4402 13252
rect 5169 13243 5227 13249
rect 5169 13209 5181 13243
rect 5215 13240 5227 13243
rect 5258 13240 5264 13252
rect 5215 13212 5264 13240
rect 5215 13209 5227 13212
rect 5169 13203 5227 13209
rect 5258 13200 5264 13212
rect 5316 13200 5322 13252
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 6917 13243 6975 13249
rect 5408 13212 5750 13240
rect 5408 13200 5414 13212
rect 6917 13209 6929 13243
rect 6963 13240 6975 13243
rect 7392 13240 7420 13268
rect 6963 13212 7420 13240
rect 6963 13209 6975 13212
rect 6917 13203 6975 13209
rect 8294 13200 8300 13252
rect 8352 13240 8358 13252
rect 8665 13243 8723 13249
rect 8665 13240 8677 13243
rect 8352 13212 8677 13240
rect 8352 13200 8358 13212
rect 8665 13209 8677 13212
rect 8711 13240 8723 13243
rect 8711 13212 9444 13240
rect 10350 13212 10732 13240
rect 8711 13209 8723 13212
rect 8665 13203 8723 13209
rect 1857 13175 1915 13181
rect 1857 13172 1869 13175
rect 1360 13144 1869 13172
rect 1360 13132 1366 13144
rect 1857 13141 1869 13144
rect 1903 13141 1915 13175
rect 1857 13135 1915 13141
rect 2961 13175 3019 13181
rect 2961 13141 2973 13175
rect 3007 13141 3019 13175
rect 2961 13135 3019 13141
rect 4246 13132 4252 13184
rect 4304 13132 4310 13184
rect 4551 13175 4609 13181
rect 4551 13141 4563 13175
rect 4597 13172 4609 13175
rect 4706 13172 4712 13184
rect 4597 13144 4712 13172
rect 4597 13141 4609 13144
rect 4551 13135 4609 13141
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 6730 13132 6736 13184
rect 6788 13172 6794 13184
rect 7377 13175 7435 13181
rect 7377 13172 7389 13175
rect 6788 13144 7389 13172
rect 6788 13132 6794 13144
rect 7377 13141 7389 13144
rect 7423 13141 7435 13175
rect 7377 13135 7435 13141
rect 9030 13132 9036 13184
rect 9088 13172 9094 13184
rect 9309 13175 9367 13181
rect 9309 13172 9321 13175
rect 9088 13144 9321 13172
rect 9088 13132 9094 13144
rect 9309 13141 9321 13144
rect 9355 13141 9367 13175
rect 9416 13172 9444 13212
rect 9858 13172 9864 13184
rect 9416 13144 9864 13172
rect 9309 13135 9367 13141
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 10704 13172 10732 13212
rect 10778 13200 10784 13252
rect 10836 13200 10842 13252
rect 12084 13240 12112 13280
rect 14090 13268 14096 13320
rect 14148 13308 14154 13320
rect 14642 13308 14648 13320
rect 14148 13280 14648 13308
rect 14148 13268 14154 13280
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 12250 13240 12256 13252
rect 10888 13212 12020 13240
rect 12084 13212 12256 13240
rect 10888 13172 10916 13212
rect 10704 13144 10916 13172
rect 11422 13132 11428 13184
rect 11480 13132 11486 13184
rect 11992 13172 12020 13212
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 12342 13200 12348 13252
rect 12400 13200 12406 13252
rect 12434 13200 12440 13252
rect 12492 13240 12498 13252
rect 14185 13243 14243 13249
rect 14185 13240 14197 13243
rect 12492 13212 12834 13240
rect 13648 13212 14197 13240
rect 12492 13200 12498 13212
rect 13648 13172 13676 13212
rect 14185 13209 14197 13212
rect 14231 13209 14243 13243
rect 14185 13203 14243 13209
rect 11992 13144 13676 13172
rect 1104 13082 14812 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 14812 13082
rect 1104 13008 14812 13030
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3510 12968 3516 12980
rect 3108 12940 3516 12968
rect 3108 12928 3114 12940
rect 3510 12928 3516 12940
rect 3568 12968 3574 12980
rect 3605 12971 3663 12977
rect 3605 12968 3617 12971
rect 3568 12940 3617 12968
rect 3568 12928 3574 12940
rect 3605 12937 3617 12940
rect 3651 12937 3663 12971
rect 3605 12931 3663 12937
rect 6178 12928 6184 12980
rect 6236 12928 6242 12980
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12968 6975 12971
rect 13262 12968 13268 12980
rect 6963 12940 13268 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 14090 12928 14096 12980
rect 14148 12928 14154 12980
rect 2406 12860 2412 12912
rect 2464 12900 2470 12912
rect 3789 12903 3847 12909
rect 3789 12900 3801 12903
rect 2464 12872 3801 12900
rect 2464 12860 2470 12872
rect 3789 12869 3801 12872
rect 3835 12869 3847 12903
rect 3989 12903 4047 12909
rect 3989 12900 4001 12903
rect 3789 12863 3847 12869
rect 3896 12872 4001 12900
rect 2498 12792 2504 12844
rect 2556 12832 2562 12844
rect 3896 12832 3924 12872
rect 3989 12869 4001 12872
rect 4035 12869 4047 12903
rect 6270 12900 6276 12912
rect 3989 12863 4047 12869
rect 4172 12872 6276 12900
rect 2556 12804 3924 12832
rect 2556 12792 2562 12804
rect 1210 12724 1216 12776
rect 1268 12764 1274 12776
rect 1268 12736 2774 12764
rect 1268 12724 1274 12736
rect 2746 12696 2774 12736
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 4172 12764 4200 12872
rect 6270 12860 6276 12872
rect 6328 12900 6334 12912
rect 6328 12872 6914 12900
rect 6328 12860 6334 12872
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 4663 12804 5181 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5169 12801 5181 12804
rect 5215 12832 5227 12835
rect 5718 12832 5724 12844
rect 5215 12804 5724 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 5994 12792 6000 12844
rect 6052 12792 6058 12844
rect 6178 12792 6184 12844
rect 6236 12792 6242 12844
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6512 12804 6561 12832
rect 6512 12792 6518 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 6886 12832 6914 12872
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 9033 12903 9091 12909
rect 9033 12900 9045 12903
rect 8352 12872 9045 12900
rect 8352 12860 8358 12872
rect 9033 12869 9045 12872
rect 9079 12869 9091 12903
rect 9033 12863 9091 12869
rect 9214 12860 9220 12912
rect 9272 12900 9278 12912
rect 12342 12900 12348 12912
rect 9272 12872 12348 12900
rect 9272 12860 9278 12872
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 6886 12804 8585 12832
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 8754 12792 8760 12844
rect 8812 12792 8818 12844
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 9180 12804 11284 12832
rect 9180 12792 9186 12804
rect 3200 12736 4200 12764
rect 3200 12724 3206 12736
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 4304 12736 8708 12764
rect 4304 12724 4310 12736
rect 4157 12699 4215 12705
rect 4157 12696 4169 12699
rect 2746 12668 4169 12696
rect 4157 12665 4169 12668
rect 4203 12665 4215 12699
rect 4157 12659 4215 12665
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12696 4583 12699
rect 4571 12668 4844 12696
rect 4571 12665 4583 12668
rect 4525 12659 4583 12665
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4540 12628 4568 12659
rect 4019 12600 4568 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4706 12588 4712 12640
rect 4764 12588 4770 12640
rect 4816 12628 4844 12668
rect 4890 12656 4896 12708
rect 4948 12696 4954 12708
rect 5813 12699 5871 12705
rect 5813 12696 5825 12699
rect 4948 12668 5825 12696
rect 4948 12656 4954 12668
rect 5813 12665 5825 12668
rect 5859 12696 5871 12699
rect 5994 12696 6000 12708
rect 5859 12668 6000 12696
rect 5859 12665 5871 12668
rect 5813 12659 5871 12665
rect 5994 12656 6000 12668
rect 6052 12696 6058 12708
rect 6638 12696 6644 12708
rect 6052 12668 6644 12696
rect 6052 12656 6058 12668
rect 6638 12656 6644 12668
rect 6696 12656 6702 12708
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 7285 12699 7343 12705
rect 7285 12696 7297 12699
rect 6788 12668 7297 12696
rect 6788 12656 6794 12668
rect 7285 12665 7297 12668
rect 7331 12696 7343 12699
rect 7558 12696 7564 12708
rect 7331 12668 7564 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 8202 12628 8208 12640
rect 4816 12600 8208 12628
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 8680 12628 8708 12736
rect 9306 12724 9312 12776
rect 9364 12764 9370 12776
rect 11146 12764 11152 12776
rect 9364 12736 11152 12764
rect 9364 12724 9370 12736
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 11256 12764 11284 12804
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12832 12495 12835
rect 14090 12832 14096 12844
rect 12483 12804 14096 12832
rect 12483 12801 12495 12804
rect 12437 12795 12495 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14200 12764 14228 12795
rect 11256 12736 14228 12764
rect 8941 12699 8999 12705
rect 8941 12665 8953 12699
rect 8987 12696 8999 12699
rect 9490 12696 9496 12708
rect 8987 12668 9496 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 11698 12696 11704 12708
rect 9640 12668 11704 12696
rect 9640 12656 9646 12668
rect 11698 12656 11704 12668
rect 11756 12696 11762 12708
rect 11977 12699 12035 12705
rect 11977 12696 11989 12699
rect 11756 12668 11989 12696
rect 11756 12656 11762 12668
rect 11977 12665 11989 12668
rect 12023 12665 12035 12699
rect 11977 12659 12035 12665
rect 12250 12656 12256 12708
rect 12308 12656 12314 12708
rect 9122 12628 9128 12640
rect 8680 12600 9128 12628
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9306 12588 9312 12640
rect 9364 12628 9370 12640
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9364 12600 10333 12628
rect 9364 12588 9370 12600
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 10321 12591 10379 12597
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 11296 12600 11621 12628
rect 11296 12588 11302 12600
rect 11609 12597 11621 12600
rect 11655 12597 11667 12631
rect 11609 12591 11667 12597
rect 13170 12588 13176 12640
rect 13228 12588 13234 12640
rect 14369 12631 14427 12637
rect 14369 12597 14381 12631
rect 14415 12628 14427 12631
rect 14826 12628 14832 12640
rect 14415 12600 14832 12628
rect 14415 12597 14427 12600
rect 14369 12591 14427 12597
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 1104 12538 14812 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 14812 12538
rect 1104 12464 14812 12486
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 3605 12427 3663 12433
rect 3605 12424 3617 12427
rect 3476 12396 3617 12424
rect 3476 12384 3482 12396
rect 3605 12393 3617 12396
rect 3651 12424 3663 12427
rect 4522 12424 4528 12436
rect 3651 12396 4528 12424
rect 3651 12393 3663 12396
rect 3605 12387 3663 12393
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 8386 12424 8392 12436
rect 5500 12396 8392 12424
rect 5500 12384 5506 12396
rect 8386 12384 8392 12396
rect 8444 12424 8450 12436
rect 9582 12424 9588 12436
rect 8444 12396 9588 12424
rect 8444 12384 8450 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 10413 12427 10471 12433
rect 10413 12393 10425 12427
rect 10459 12424 10471 12427
rect 10870 12424 10876 12436
rect 10459 12396 10876 12424
rect 10459 12393 10471 12396
rect 10413 12387 10471 12393
rect 10870 12384 10876 12396
rect 10928 12424 10934 12436
rect 10928 12396 11560 12424
rect 10928 12384 10934 12396
rect 8110 12316 8116 12368
rect 8168 12356 8174 12368
rect 8294 12356 8300 12368
rect 8168 12328 8300 12356
rect 8168 12316 8174 12328
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 8846 12316 8852 12368
rect 8904 12356 8910 12368
rect 10134 12356 10140 12368
rect 8904 12328 10140 12356
rect 8904 12316 8910 12328
rect 10134 12316 10140 12328
rect 10192 12316 10198 12368
rect 11532 12365 11560 12396
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12529 12427 12587 12433
rect 12529 12424 12541 12427
rect 12032 12396 12541 12424
rect 12032 12384 12038 12396
rect 12529 12393 12541 12396
rect 12575 12393 12587 12427
rect 12529 12387 12587 12393
rect 13262 12384 13268 12436
rect 13320 12384 13326 12436
rect 11517 12359 11575 12365
rect 11517 12325 11529 12359
rect 11563 12356 11575 12359
rect 15010 12356 15016 12368
rect 11563 12328 15016 12356
rect 11563 12325 11575 12328
rect 11517 12319 11575 12325
rect 15010 12316 15016 12328
rect 15068 12316 15074 12368
rect 4338 12248 4344 12300
rect 4396 12288 4402 12300
rect 4522 12288 4528 12300
rect 4396 12260 4528 12288
rect 4396 12248 4402 12260
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 5684 12260 6469 12288
rect 5684 12248 5690 12260
rect 6380 12229 6408 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 6788 12260 8984 12288
rect 6788 12248 6794 12260
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6411 12192 6445 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 8386 12220 8392 12232
rect 6604 12192 8392 12220
rect 6604 12180 6610 12192
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 8956 12220 8984 12260
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 13633 12291 13691 12297
rect 13633 12288 13645 12291
rect 9732 12260 13645 12288
rect 9732 12248 9738 12260
rect 13633 12257 13645 12260
rect 13679 12257 13691 12291
rect 13633 12251 13691 12257
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 8956 12192 10149 12220
rect 10137 12189 10149 12192
rect 10183 12220 10195 12223
rect 10318 12220 10324 12232
rect 10183 12192 10324 12220
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 10318 12180 10324 12192
rect 10376 12220 10382 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 10376 12192 10793 12220
rect 10376 12180 10382 12192
rect 10781 12189 10793 12192
rect 10827 12220 10839 12223
rect 10962 12220 10968 12232
rect 10827 12192 10968 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 11572 12192 12173 12220
rect 11572 12180 11578 12192
rect 12161 12189 12173 12192
rect 12207 12220 12219 12223
rect 12526 12220 12532 12232
rect 12207 12192 12532 12220
rect 12207 12189 12219 12192
rect 12161 12183 12219 12189
rect 12526 12180 12532 12192
rect 12584 12220 12590 12232
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 12584 12192 12725 12220
rect 12584 12180 12590 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 12894 12180 12900 12232
rect 12952 12180 12958 12232
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 4764 12124 4922 12152
rect 4764 12112 4770 12124
rect 6086 12112 6092 12164
rect 6144 12112 6150 12164
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7742 12152 7748 12164
rect 6972 12124 7748 12152
rect 6972 12112 6978 12124
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 8202 12112 8208 12164
rect 8260 12112 8266 12164
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 9125 12155 9183 12161
rect 9125 12152 9137 12155
rect 8628 12124 9137 12152
rect 8628 12112 8634 12124
rect 9125 12121 9137 12124
rect 9171 12152 9183 12155
rect 9306 12152 9312 12164
rect 9171 12124 9312 12152
rect 9171 12121 9183 12124
rect 9125 12115 9183 12121
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 10870 12152 10876 12164
rect 9416 12124 10876 12152
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 9416 12084 9444 12124
rect 10870 12112 10876 12124
rect 10928 12112 10934 12164
rect 13004 12152 13032 12183
rect 13262 12180 13268 12232
rect 13320 12220 13326 12232
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 13320 12192 13553 12220
rect 13320 12180 13326 12192
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 11808 12124 13032 12152
rect 11808 12096 11836 12124
rect 13446 12112 13452 12164
rect 13504 12112 13510 12164
rect 3660 12056 9444 12084
rect 3660 12044 3666 12056
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 10229 12087 10287 12093
rect 10229 12084 10241 12087
rect 10192 12056 10241 12084
rect 10192 12044 10198 12056
rect 10229 12053 10241 12056
rect 10275 12053 10287 12087
rect 10229 12047 10287 12053
rect 10413 12087 10471 12093
rect 10413 12053 10425 12087
rect 10459 12084 10471 12087
rect 10502 12084 10508 12096
rect 10459 12056 10508 12084
rect 10459 12053 10471 12056
rect 10413 12047 10471 12053
rect 10502 12044 10508 12056
rect 10560 12084 10566 12096
rect 10962 12084 10968 12096
rect 10560 12056 10968 12084
rect 10560 12044 10566 12056
rect 10962 12044 10968 12056
rect 11020 12084 11026 12096
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 11020 12056 11069 12084
rect 11020 12044 11026 12056
rect 11057 12053 11069 12056
rect 11103 12053 11115 12087
rect 11057 12047 11115 12053
rect 11790 12044 11796 12096
rect 11848 12044 11854 12096
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 13081 12087 13139 12093
rect 13081 12084 13093 12087
rect 13044 12056 13093 12084
rect 13044 12044 13050 12056
rect 13081 12053 13093 12056
rect 13127 12053 13139 12087
rect 13081 12047 13139 12053
rect 13249 12087 13307 12093
rect 13249 12053 13261 12087
rect 13295 12084 13307 12087
rect 13538 12084 13544 12096
rect 13295 12056 13544 12084
rect 13295 12053 13307 12056
rect 13249 12047 13307 12053
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 14458 12044 14464 12096
rect 14516 12044 14522 12096
rect 1104 11994 14812 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 14812 11994
rect 1104 11920 14812 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3237 11883 3295 11889
rect 3237 11880 3249 11883
rect 3016 11852 3249 11880
rect 3016 11840 3022 11852
rect 3237 11849 3249 11852
rect 3283 11849 3295 11883
rect 3237 11843 3295 11849
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 4157 11883 4215 11889
rect 4157 11880 4169 11883
rect 3743 11852 4169 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 4157 11849 4169 11852
rect 4203 11880 4215 11883
rect 8386 11880 8392 11892
rect 4203 11852 8392 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 11514 11880 11520 11892
rect 8628 11852 11520 11880
rect 8628 11840 8634 11852
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 11793 11883 11851 11889
rect 11793 11849 11805 11883
rect 11839 11880 11851 11883
rect 11839 11852 12020 11880
rect 11839 11849 11851 11852
rect 11793 11843 11851 11849
rect 4706 11772 4712 11824
rect 4764 11772 4770 11824
rect 4890 11772 4896 11824
rect 4948 11812 4954 11824
rect 5166 11812 5172 11824
rect 4948 11784 5172 11812
rect 4948 11772 4954 11784
rect 5166 11772 5172 11784
rect 5224 11812 5230 11824
rect 5626 11812 5632 11824
rect 5224 11784 5632 11812
rect 5224 11772 5230 11784
rect 5626 11772 5632 11784
rect 5684 11772 5690 11824
rect 6549 11815 6607 11821
rect 6549 11781 6561 11815
rect 6595 11812 6607 11815
rect 9674 11812 9680 11824
rect 6595 11784 9680 11812
rect 6595 11781 6607 11784
rect 6549 11775 6607 11781
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 10042 11772 10048 11824
rect 10100 11772 10106 11824
rect 11992 11812 12020 11852
rect 12066 11840 12072 11892
rect 12124 11840 12130 11892
rect 12989 11883 13047 11889
rect 12989 11849 13001 11883
rect 13035 11880 13047 11883
rect 13446 11880 13452 11892
rect 13035 11852 13452 11880
rect 13035 11849 13047 11852
rect 12989 11843 13047 11849
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 14918 11840 14924 11892
rect 14976 11880 14982 11892
rect 15194 11880 15200 11892
rect 14976 11852 15200 11880
rect 14976 11840 14982 11852
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 12437 11815 12495 11821
rect 12437 11812 12449 11815
rect 11348 11784 11836 11812
rect 11992 11784 12449 11812
rect 2774 11704 2780 11756
rect 2832 11704 2838 11756
rect 3296 11747 3354 11753
rect 3296 11713 3308 11747
rect 3342 11744 3354 11747
rect 3418 11744 3424 11756
rect 3342 11716 3424 11744
rect 3342 11713 3354 11716
rect 3296 11707 3354 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11744 3571 11747
rect 3602 11744 3608 11756
rect 3559 11716 3608 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 4246 11744 4252 11756
rect 3835 11716 4252 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4571 11716 4629 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4617 11713 4629 11716
rect 4663 11744 4675 11747
rect 5442 11744 5448 11756
rect 4663 11716 5448 11744
rect 4663 11713 4675 11716
rect 4617 11707 4675 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 4706 11636 4712 11688
rect 4764 11676 4770 11688
rect 5534 11676 5540 11688
rect 4764 11648 5540 11676
rect 4764 11636 4770 11648
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 4062 11608 4068 11620
rect 2915 11580 4068 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 5828 11608 5856 11707
rect 6270 11704 6276 11756
rect 6328 11744 6334 11756
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 6328 11716 6469 11744
rect 6328 11704 6334 11716
rect 6457 11713 6469 11716
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 6696 11716 6745 11744
rect 6696 11704 6702 11716
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 7098 11704 7104 11756
rect 7156 11704 7162 11756
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11744 7251 11747
rect 8294 11744 8300 11756
rect 7239 11716 8300 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 8294 11704 8300 11716
rect 8352 11704 8358 11756
rect 11348 11753 11376 11784
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8588 11716 8953 11744
rect 8588 11688 8616 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11744 11391 11747
rect 11514 11744 11520 11756
rect 11379 11716 11520 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 11698 11704 11704 11756
rect 11756 11704 11762 11756
rect 11808 11744 11836 11784
rect 12437 11781 12449 11784
rect 12483 11812 12495 11815
rect 13814 11812 13820 11824
rect 12483 11784 13820 11812
rect 12483 11781 12495 11784
rect 12437 11775 12495 11781
rect 13814 11772 13820 11784
rect 13872 11772 13878 11824
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11808 11716 11897 11744
rect 11885 11713 11897 11716
rect 11931 11744 11943 11747
rect 14274 11744 14280 11756
rect 11931 11716 14280 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 6917 11679 6975 11685
rect 6917 11645 6929 11679
rect 6963 11676 6975 11679
rect 7742 11676 7748 11688
rect 6963 11648 7748 11676
rect 6963 11645 6975 11648
rect 6917 11639 6975 11645
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 8481 11679 8539 11685
rect 8481 11645 8493 11679
rect 8527 11676 8539 11679
rect 8570 11676 8576 11688
rect 8527 11648 8576 11676
rect 8527 11645 8539 11648
rect 8481 11639 8539 11645
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 8754 11685 8760 11688
rect 8732 11679 8760 11685
rect 8732 11645 8744 11679
rect 8732 11639 8760 11645
rect 8754 11636 8760 11639
rect 8812 11636 8818 11688
rect 8846 11636 8852 11688
rect 8904 11636 8910 11688
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11645 9275 11679
rect 9217 11639 9275 11645
rect 8864 11608 8892 11636
rect 5828 11580 8892 11608
rect 2685 11543 2743 11549
rect 2685 11509 2697 11543
rect 2731 11540 2743 11543
rect 2958 11540 2964 11552
rect 2731 11512 2964 11540
rect 2731 11509 2743 11512
rect 2685 11503 2743 11509
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 3418 11500 3424 11552
rect 3476 11500 3482 11552
rect 3510 11500 3516 11552
rect 3568 11500 3574 11552
rect 4080 11540 4108 11568
rect 5534 11540 5540 11552
rect 4080 11512 5540 11540
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 6546 11540 6552 11552
rect 5776 11512 6552 11540
rect 5776 11500 5782 11512
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 7561 11543 7619 11549
rect 7561 11509 7573 11543
rect 7607 11540 7619 11543
rect 8294 11540 8300 11552
rect 7607 11512 8300 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8570 11500 8576 11552
rect 8628 11500 8634 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9232 11540 9260 11639
rect 9306 11636 9312 11688
rect 9364 11636 9370 11688
rect 9582 11636 9588 11688
rect 9640 11636 9646 11688
rect 11422 11568 11428 11620
rect 11480 11608 11486 11620
rect 11517 11611 11575 11617
rect 11517 11608 11529 11611
rect 11480 11580 11529 11608
rect 11480 11568 11486 11580
rect 11517 11577 11529 11580
rect 11563 11577 11575 11611
rect 13446 11608 13452 11620
rect 11517 11571 11575 11577
rect 12406 11580 13452 11608
rect 8904 11512 9260 11540
rect 8904 11500 8910 11512
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 12406 11540 12434 11580
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 10744 11512 12434 11540
rect 10744 11500 10750 11512
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 13262 11540 13268 11552
rect 12952 11512 13268 11540
rect 12952 11500 12958 11512
rect 13262 11500 13268 11512
rect 13320 11540 13326 11552
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 13320 11512 13369 11540
rect 13320 11500 13326 11512
rect 13357 11509 13369 11512
rect 13403 11509 13415 11543
rect 13357 11503 13415 11509
rect 1104 11450 14812 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 14812 11450
rect 1104 11376 14812 11398
rect 1486 11296 1492 11348
rect 1544 11336 1550 11348
rect 2590 11336 2596 11348
rect 1544 11308 2596 11336
rect 1544 11296 1550 11308
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3602 11336 3608 11348
rect 2832 11308 3608 11336
rect 2832 11296 2838 11308
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 5166 11336 5172 11348
rect 3804 11308 5172 11336
rect 3142 11160 3148 11212
rect 3200 11200 3206 11212
rect 3694 11200 3700 11212
rect 3200 11172 3700 11200
rect 3200 11160 3206 11172
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 3804 11209 3832 11308
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 7006 11336 7012 11348
rect 5592 11308 7012 11336
rect 5592 11296 5598 11308
rect 7006 11296 7012 11308
rect 7064 11336 7070 11348
rect 7064 11308 8800 11336
rect 7064 11296 7070 11308
rect 3970 11228 3976 11280
rect 4028 11228 4034 11280
rect 4065 11271 4123 11277
rect 4065 11237 4077 11271
rect 4111 11268 4123 11271
rect 4338 11268 4344 11280
rect 4111 11240 4344 11268
rect 4111 11237 4123 11240
rect 4065 11231 4123 11237
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 6641 11271 6699 11277
rect 6641 11237 6653 11271
rect 6687 11268 6699 11271
rect 7650 11268 7656 11280
rect 6687 11240 7656 11268
rect 6687 11237 6699 11240
rect 6641 11231 6699 11237
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 8772 11268 8800 11308
rect 8938 11296 8944 11348
rect 8996 11296 9002 11348
rect 9048 11308 13216 11336
rect 9048 11268 9076 11308
rect 7892 11240 8708 11268
rect 8772 11240 9076 11268
rect 7892 11228 7898 11240
rect 3789 11203 3847 11209
rect 3789 11169 3801 11203
rect 3835 11169 3847 11203
rect 4525 11203 4583 11209
rect 3789 11163 3847 11169
rect 3896 11172 4384 11200
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 3896 11132 3924 11172
rect 1636 11104 3924 11132
rect 4065 11135 4123 11141
rect 1636 11092 1642 11104
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4246 11132 4252 11144
rect 4111 11104 4252 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 3237 11067 3295 11073
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 4154 11064 4160 11076
rect 3283 11036 4160 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 4356 11064 4384 11172
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 4890 11200 4896 11212
rect 4571 11172 4896 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 7006 11200 7012 11212
rect 5408 11172 6684 11200
rect 5408 11160 5414 11172
rect 6656 11141 6684 11172
rect 6748 11172 7012 11200
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 4801 11067 4859 11073
rect 4801 11064 4813 11067
rect 4356 11036 4813 11064
rect 4801 11033 4813 11036
rect 4847 11033 4859 11067
rect 6454 11064 6460 11076
rect 6026 11036 6460 11064
rect 4801 11027 4859 11033
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 6549 11067 6607 11073
rect 6549 11033 6561 11067
rect 6595 11064 6607 11067
rect 6748 11064 6776 11172
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 7190 11160 7196 11212
rect 7248 11200 7254 11212
rect 8570 11200 8576 11212
rect 7248 11172 8576 11200
rect 7248 11160 7254 11172
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 7282 11132 7288 11144
rect 6963 11104 7288 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 7282 11092 7288 11104
rect 7340 11132 7346 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7340 11104 7573 11132
rect 7340 11092 7346 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8294 11132 8300 11144
rect 8159 11104 8300 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8294 11092 8300 11104
rect 8352 11132 8358 11144
rect 8680 11132 8708 11240
rect 9306 11228 9312 11280
rect 9364 11228 9370 11280
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 12894 11268 12900 11280
rect 11204 11240 12900 11268
rect 11204 11228 11210 11240
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 12989 11271 13047 11277
rect 12989 11237 13001 11271
rect 13035 11268 13047 11271
rect 13078 11268 13084 11280
rect 13035 11240 13084 11268
rect 13035 11237 13047 11240
rect 12989 11231 13047 11237
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 9324 11200 9352 11228
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 9324 11172 10701 11200
rect 10689 11169 10701 11172
rect 10735 11169 10747 11203
rect 10689 11163 10747 11169
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 11514 11200 11520 11212
rect 11471 11172 11520 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 12434 11160 12440 11212
rect 12492 11160 12498 11212
rect 12526 11160 12532 11212
rect 12584 11160 12590 11212
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 12860 11172 13124 11200
rect 12860 11160 12866 11172
rect 8352 11104 8524 11132
rect 8680 11104 9338 11132
rect 8352 11092 8358 11104
rect 8496 11076 8524 11104
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 12544 11132 12572 11160
rect 11020 11104 12572 11132
rect 12621 11135 12679 11141
rect 11020 11092 11026 11104
rect 12621 11101 12633 11135
rect 12667 11132 12679 11135
rect 12986 11132 12992 11144
rect 12667 11104 12992 11132
rect 12667 11101 12679 11104
rect 12621 11095 12679 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13096 11141 13124 11172
rect 13188 11141 13216 11308
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 6595 11036 6776 11064
rect 6825 11067 6883 11073
rect 6595 11033 6607 11036
rect 6549 11027 6607 11033
rect 6825 11033 6837 11067
rect 6871 11033 6883 11067
rect 6825 11027 6883 11033
rect 3145 10999 3203 11005
rect 3145 10965 3157 10999
rect 3191 10996 3203 10999
rect 4614 10996 4620 11008
rect 3191 10968 4620 10996
rect 3191 10965 3203 10968
rect 3145 10959 3203 10965
rect 4614 10956 4620 10968
rect 4672 10996 4678 11008
rect 4890 10996 4896 11008
rect 4672 10968 4896 10996
rect 4672 10956 4678 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 6178 10956 6184 11008
rect 6236 10996 6242 11008
rect 6638 10996 6644 11008
rect 6236 10968 6644 10996
rect 6236 10956 6242 10968
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 6840 10996 6868 11027
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7834 11064 7840 11076
rect 7064 11036 7840 11064
rect 7064 11024 7070 11036
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8478 11024 8484 11076
rect 8536 11024 8542 11076
rect 10413 11067 10471 11073
rect 10413 11033 10425 11067
rect 10459 11064 10471 11067
rect 12250 11064 12256 11076
rect 10459 11036 12256 11064
rect 10459 11033 10471 11036
rect 10413 11027 10471 11033
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12802 11024 12808 11076
rect 12860 11024 12866 11076
rect 13096 11064 13124 11095
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 13320 11104 13369 11132
rect 13320 11092 13326 11104
rect 13357 11101 13369 11104
rect 13403 11132 13415 11135
rect 13725 11135 13783 11141
rect 13725 11132 13737 11135
rect 13403 11104 13737 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 13725 11101 13737 11104
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 13538 11064 13544 11076
rect 13096 11036 13544 11064
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 13814 11064 13820 11076
rect 13688 11036 13820 11064
rect 13688 11024 13694 11036
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14458 11024 14464 11076
rect 14516 11024 14522 11076
rect 7098 10996 7104 11008
rect 6840 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10996 7162 11008
rect 7193 10999 7251 11005
rect 7193 10996 7205 10999
rect 7156 10968 7205 10996
rect 7156 10956 7162 10968
rect 7193 10965 7205 10968
rect 7239 10965 7251 10999
rect 7193 10959 7251 10965
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 8021 10999 8079 11005
rect 8021 10996 8033 10999
rect 7340 10968 8033 10996
rect 7340 10956 7346 10968
rect 8021 10965 8033 10968
rect 8067 10965 8079 10999
rect 12820 10996 12848 11024
rect 12986 10996 12992 11008
rect 12820 10968 12992 10996
rect 8021 10959 8079 10965
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 1104 10906 14812 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 14812 10906
rect 1104 10832 14812 10854
rect 2406 10752 2412 10804
rect 2464 10752 2470 10804
rect 3326 10752 3332 10804
rect 3384 10752 3390 10804
rect 3697 10795 3755 10801
rect 3697 10761 3709 10795
rect 3743 10792 3755 10795
rect 4706 10792 4712 10804
rect 3743 10764 4712 10792
rect 3743 10761 3755 10764
rect 3697 10755 3755 10761
rect 2133 10727 2191 10733
rect 2133 10693 2145 10727
rect 2179 10724 2191 10727
rect 2179 10696 3096 10724
rect 2179 10693 2191 10696
rect 2133 10687 2191 10693
rect 2240 10665 2268 10696
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2409 10659 2467 10665
rect 2271 10628 2305 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2409 10625 2421 10659
rect 2455 10656 2467 10659
rect 2774 10656 2780 10668
rect 2455 10628 2780 10656
rect 2455 10625 2467 10628
rect 2409 10619 2467 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 3068 10588 3096 10696
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10656 3387 10659
rect 3712 10656 3740 10755
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10761 5135 10795
rect 5077 10755 5135 10761
rect 5092 10724 5120 10755
rect 5258 10752 5264 10804
rect 5316 10752 5322 10804
rect 5629 10795 5687 10801
rect 5629 10761 5641 10795
rect 5675 10792 5687 10795
rect 6362 10792 6368 10804
rect 5675 10764 6368 10792
rect 5675 10761 5687 10764
rect 5629 10755 5687 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 7282 10792 7288 10804
rect 6696 10764 7288 10792
rect 6696 10752 6702 10764
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 9030 10792 9036 10804
rect 7616 10764 9036 10792
rect 7616 10752 7622 10764
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 12069 10795 12127 10801
rect 12069 10792 12081 10795
rect 10376 10764 12081 10792
rect 10376 10752 10382 10764
rect 12069 10761 12081 10764
rect 12115 10792 12127 10795
rect 12526 10792 12532 10804
rect 12115 10764 12532 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 13780 10764 14381 10792
rect 13780 10752 13786 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 14369 10755 14427 10761
rect 5902 10724 5908 10736
rect 5092 10696 5908 10724
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 6914 10684 6920 10736
rect 6972 10724 6978 10736
rect 7437 10727 7495 10733
rect 7437 10724 7449 10727
rect 6972 10696 7449 10724
rect 6972 10684 6978 10696
rect 7437 10693 7449 10696
rect 7483 10693 7495 10727
rect 7653 10727 7711 10733
rect 7653 10724 7665 10727
rect 7437 10687 7495 10693
rect 7576 10696 7665 10724
rect 3375 10628 3740 10656
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 4430 10616 4436 10668
rect 4488 10656 4494 10668
rect 4488 10628 5396 10656
rect 4488 10616 4494 10628
rect 5368 10600 5396 10628
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 5868 10628 6193 10656
rect 5868 10616 5874 10628
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6362 10616 6368 10668
rect 6420 10656 6426 10668
rect 6822 10656 6828 10668
rect 6420 10628 6828 10656
rect 6420 10616 6426 10628
rect 6822 10616 6828 10628
rect 6880 10656 6886 10668
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 6880 10654 6914 10656
rect 7024 10654 7205 10656
rect 6880 10628 7205 10654
rect 6880 10626 7052 10628
rect 6880 10616 6886 10626
rect 7193 10625 7205 10628
rect 7239 10656 7251 10659
rect 7239 10654 7420 10656
rect 7576 10654 7604 10696
rect 7653 10693 7665 10696
rect 7699 10693 7711 10727
rect 7653 10687 7711 10693
rect 9858 10684 9864 10736
rect 9916 10724 9922 10736
rect 10229 10727 10287 10733
rect 10229 10724 10241 10727
rect 9916 10696 10241 10724
rect 9916 10684 9922 10696
rect 10229 10693 10241 10696
rect 10275 10724 10287 10727
rect 10686 10724 10692 10736
rect 10275 10696 10692 10724
rect 10275 10693 10287 10696
rect 10229 10687 10287 10693
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 12342 10684 12348 10736
rect 12400 10684 12406 10736
rect 7239 10628 7604 10654
rect 7239 10625 7251 10628
rect 7392 10626 7604 10628
rect 7193 10619 7251 10625
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 7800 10628 8984 10656
rect 7800 10616 7806 10628
rect 4706 10588 4712 10600
rect 3068 10560 4712 10588
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 4985 10591 5043 10597
rect 4985 10588 4997 10591
rect 4948 10560 4997 10588
rect 4948 10548 4954 10560
rect 4985 10557 4997 10560
rect 5031 10557 5043 10591
rect 4985 10551 5043 10557
rect 5350 10548 5356 10600
rect 5408 10548 5414 10600
rect 5442 10548 5448 10600
rect 5500 10548 5506 10600
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 6730 10588 6736 10600
rect 6328 10560 6736 10588
rect 6328 10548 6334 10560
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 8846 10588 8852 10600
rect 7024 10560 8852 10588
rect 1670 10480 1676 10532
rect 1728 10520 1734 10532
rect 5997 10523 6055 10529
rect 5997 10520 6009 10523
rect 1728 10492 6009 10520
rect 1728 10480 1734 10492
rect 5997 10489 6009 10492
rect 6043 10489 6055 10523
rect 7024 10520 7052 10560
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 8956 10588 8984 10628
rect 9214 10616 9220 10668
rect 9272 10656 9278 10668
rect 9987 10659 10045 10665
rect 9987 10656 9999 10659
rect 9272 10628 9999 10656
rect 9272 10616 9278 10628
rect 9987 10625 9999 10628
rect 10033 10625 10045 10659
rect 9987 10619 10045 10625
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 11514 10656 11520 10668
rect 10652 10628 11520 10656
rect 10652 10616 10658 10628
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 12434 10616 12440 10668
rect 12492 10616 12498 10668
rect 12526 10616 12532 10668
rect 12584 10616 12590 10668
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12768 10628 13001 10656
rect 12768 10616 12774 10628
rect 12989 10625 13001 10628
rect 13035 10656 13047 10659
rect 13262 10656 13268 10668
rect 13035 10628 13268 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 13446 10616 13452 10668
rect 13504 10616 13510 10668
rect 13630 10656 13636 10668
rect 13556 10628 13636 10656
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 8956 10560 9597 10588
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 9674 10548 9680 10600
rect 9732 10548 9738 10600
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 13556 10588 13584 10628
rect 13630 10616 13636 10628
rect 13688 10656 13694 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 13688 10628 14197 10656
rect 13688 10616 13694 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 14274 10616 14280 10668
rect 14332 10656 14338 10668
rect 14461 10659 14519 10665
rect 14461 10656 14473 10659
rect 14332 10628 14473 10656
rect 14332 10616 14338 10628
rect 14461 10625 14473 10628
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 12676 10560 13584 10588
rect 13725 10591 13783 10597
rect 12676 10548 12682 10560
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 14642 10588 14648 10600
rect 13771 10560 14648 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 5997 10483 6055 10489
rect 6380 10492 7052 10520
rect 7285 10523 7343 10529
rect 6380 10464 6408 10492
rect 7285 10489 7297 10523
rect 7331 10489 7343 10523
rect 10502 10520 10508 10532
rect 7285 10483 7343 10489
rect 7484 10492 10508 10520
rect 2774 10412 2780 10464
rect 2832 10412 2838 10464
rect 3418 10412 3424 10464
rect 3476 10452 3482 10464
rect 5442 10452 5448 10464
rect 3476 10424 5448 10452
rect 3476 10412 3482 10424
rect 5442 10412 5448 10424
rect 5500 10452 5506 10464
rect 6362 10452 6368 10464
rect 5500 10424 6368 10452
rect 5500 10412 5506 10424
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 7300 10452 7328 10483
rect 7484 10461 7512 10492
rect 10502 10480 10508 10492
rect 10560 10480 10566 10532
rect 12526 10480 12532 10532
rect 12584 10480 12590 10532
rect 6788 10424 7328 10452
rect 7469 10455 7527 10461
rect 6788 10412 6794 10424
rect 7469 10421 7481 10455
rect 7515 10421 7527 10455
rect 7469 10415 7527 10421
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 11514 10452 11520 10464
rect 8536 10424 11520 10452
rect 8536 10412 8542 10424
rect 11514 10412 11520 10424
rect 11572 10452 11578 10464
rect 11793 10455 11851 10461
rect 11793 10452 11805 10455
rect 11572 10424 11805 10452
rect 11572 10412 11578 10424
rect 11793 10421 11805 10424
rect 11839 10452 11851 10455
rect 12434 10452 12440 10464
rect 11839 10424 12440 10452
rect 11839 10421 11851 10424
rect 11793 10415 11851 10421
rect 12434 10412 12440 10424
rect 12492 10452 12498 10464
rect 13740 10452 13768 10551
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 12492 10424 13768 10452
rect 14001 10455 14059 10461
rect 12492 10412 12498 10424
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 15010 10452 15016 10464
rect 14047 10424 15016 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 1104 10362 14812 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 14812 10362
rect 1104 10288 14812 10310
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2958 10248 2964 10260
rect 2280 10220 2964 10248
rect 2280 10208 2286 10220
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 3234 10208 3240 10260
rect 3292 10248 3298 10260
rect 4154 10248 4160 10260
rect 3292 10220 4160 10248
rect 3292 10208 3298 10220
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 5684 10220 6592 10248
rect 5684 10208 5690 10220
rect 3326 10140 3332 10192
rect 3384 10180 3390 10192
rect 4522 10180 4528 10192
rect 3384 10152 4528 10180
rect 3384 10140 3390 10152
rect 4522 10140 4528 10152
rect 4580 10140 4586 10192
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 6086 10180 6092 10192
rect 5408 10152 6092 10180
rect 5408 10140 5414 10152
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 5534 10112 5540 10124
rect 3936 10084 5540 10112
rect 3936 10072 3942 10084
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 6564 10121 6592 10220
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 10413 10251 10471 10257
rect 10413 10248 10425 10251
rect 6972 10220 10425 10248
rect 6972 10208 6978 10220
rect 10413 10217 10425 10220
rect 10459 10217 10471 10251
rect 10413 10211 10471 10217
rect 10502 10208 10508 10260
rect 10560 10248 10566 10260
rect 10560 10220 12848 10248
rect 10560 10208 10566 10220
rect 9490 10140 9496 10192
rect 9548 10180 9554 10192
rect 9548 10152 11652 10180
rect 9548 10140 9554 10152
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 8018 10112 8024 10124
rect 6871 10084 8024 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8478 10072 8484 10124
rect 8536 10112 8542 10124
rect 11054 10112 11060 10124
rect 8536 10084 11060 10112
rect 8536 10072 8542 10084
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 5258 10044 5264 10056
rect 4212 10016 5264 10044
rect 4212 10004 4218 10016
rect 5258 10004 5264 10016
rect 5316 10044 5322 10056
rect 6270 10044 6276 10056
rect 5316 10016 6276 10044
rect 5316 10004 5322 10016
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9692 10016 9965 10044
rect 3142 9936 3148 9988
rect 3200 9976 3206 9988
rect 6546 9976 6552 9988
rect 3200 9948 6552 9976
rect 3200 9936 3206 9948
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 8386 9976 8392 9988
rect 8050 9948 8392 9976
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 9692 9920 9720 10016
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 10226 10004 10232 10056
rect 10284 10004 10290 10056
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10044 10563 10047
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10551 10016 10977 10044
rect 10551 10013 10563 10016
rect 10505 10007 10563 10013
rect 10965 10013 10977 10016
rect 11011 10044 11023 10047
rect 11514 10044 11520 10056
rect 11011 10016 11520 10044
rect 11011 10013 11023 10016
rect 10965 10007 11023 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11624 10044 11652 10152
rect 11698 10140 11704 10192
rect 11756 10180 11762 10192
rect 12618 10180 12624 10192
rect 11756 10152 12624 10180
rect 11756 10140 11762 10152
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 12820 10180 12848 10220
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 13044 10220 13308 10248
rect 13044 10208 13050 10220
rect 12820 10152 13216 10180
rect 12986 10072 12992 10124
rect 13044 10072 13050 10124
rect 12069 10047 12127 10053
rect 12069 10044 12081 10047
rect 11624 10016 12081 10044
rect 12069 10013 12081 10016
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12618 10044 12624 10056
rect 12483 10016 12624 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10686 9976 10692 9988
rect 10100 9948 10692 9976
rect 10100 9936 10106 9948
rect 10686 9936 10692 9948
rect 10744 9936 10750 9988
rect 11054 9936 11060 9988
rect 11112 9976 11118 9988
rect 11238 9976 11244 9988
rect 11112 9948 11244 9976
rect 11112 9936 11118 9948
rect 11238 9936 11244 9948
rect 11296 9936 11302 9988
rect 12084 9976 12112 10007
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 13188 10053 13216 10152
rect 13280 10112 13308 10220
rect 13354 10208 13360 10260
rect 13412 10208 13418 10260
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13633 10251 13691 10257
rect 13633 10248 13645 10251
rect 13504 10220 13645 10248
rect 13504 10208 13510 10220
rect 13633 10217 13645 10220
rect 13679 10217 13691 10251
rect 13633 10211 13691 10217
rect 13354 10112 13360 10124
rect 13280 10084 13360 10112
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 12728 9976 12756 10007
rect 12084 9948 12756 9976
rect 12897 9979 12955 9985
rect 12897 9945 12909 9979
rect 12943 9976 12955 9979
rect 13446 9976 13452 9988
rect 12943 9948 13452 9976
rect 12943 9945 12955 9948
rect 12897 9939 12955 9945
rect 13446 9936 13452 9948
rect 13504 9976 13510 9988
rect 13814 9976 13820 9988
rect 13504 9948 13820 9976
rect 13504 9936 13510 9948
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 5534 9908 5540 9920
rect 2832 9880 5540 9908
rect 2832 9868 2838 9880
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5902 9868 5908 9920
rect 5960 9908 5966 9920
rect 6730 9908 6736 9920
rect 5960 9880 6736 9908
rect 5960 9868 5966 9880
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 6822 9868 6828 9920
rect 6880 9908 6886 9920
rect 8202 9908 8208 9920
rect 6880 9880 8208 9908
rect 6880 9868 6886 9880
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 9214 9908 9220 9920
rect 8343 9880 9220 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 9674 9868 9680 9920
rect 9732 9868 9738 9920
rect 9858 9868 9864 9920
rect 9916 9868 9922 9920
rect 10597 9911 10655 9917
rect 10597 9877 10609 9911
rect 10643 9908 10655 9911
rect 11698 9908 11704 9920
rect 10643 9880 11704 9908
rect 10643 9877 10655 9880
rect 10597 9871 10655 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 11790 9868 11796 9920
rect 11848 9908 11854 9920
rect 12253 9911 12311 9917
rect 12253 9908 12265 9911
rect 11848 9880 12265 9908
rect 11848 9868 11854 9880
rect 12253 9877 12265 9880
rect 12299 9877 12311 9911
rect 12253 9871 12311 9877
rect 12621 9911 12679 9917
rect 12621 9877 12633 9911
rect 12667 9908 12679 9911
rect 13078 9908 13084 9920
rect 12667 9880 13084 9908
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 14458 9868 14464 9920
rect 14516 9868 14522 9920
rect 1104 9818 14812 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 14812 9818
rect 1104 9744 14812 9766
rect 3697 9707 3755 9713
rect 3697 9673 3709 9707
rect 3743 9704 3755 9707
rect 4246 9704 4252 9716
rect 3743 9676 4252 9704
rect 3743 9673 3755 9676
rect 3697 9667 3755 9673
rect 4246 9664 4252 9676
rect 4304 9704 4310 9716
rect 4430 9704 4436 9716
rect 4304 9676 4436 9704
rect 4304 9664 4310 9676
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 5350 9704 5356 9716
rect 4540 9676 5356 9704
rect 3050 9636 3056 9648
rect 2700 9608 3056 9636
rect 842 9528 848 9580
rect 900 9568 906 9580
rect 1486 9568 1492 9580
rect 900 9540 1492 9568
rect 900 9528 906 9540
rect 1486 9528 1492 9540
rect 1544 9528 1550 9580
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 2222 9500 2228 9512
rect 1360 9472 2228 9500
rect 1360 9460 1366 9472
rect 2222 9460 2228 9472
rect 2280 9500 2286 9512
rect 2317 9503 2375 9509
rect 2317 9500 2329 9503
rect 2280 9472 2329 9500
rect 2280 9460 2286 9472
rect 2317 9469 2329 9472
rect 2363 9500 2375 9503
rect 2363 9472 2544 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 1486 9392 1492 9444
rect 1544 9432 1550 9444
rect 2409 9435 2467 9441
rect 2409 9432 2421 9435
rect 1544 9404 2421 9432
rect 1544 9392 1550 9404
rect 2409 9401 2421 9404
rect 2455 9401 2467 9435
rect 2516 9432 2544 9472
rect 2590 9460 2596 9512
rect 2648 9500 2654 9512
rect 2700 9509 2728 9608
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 4540 9636 4568 9676
rect 5350 9664 5356 9676
rect 5408 9704 5414 9716
rect 5626 9704 5632 9716
rect 5408 9676 5632 9704
rect 5408 9664 5414 9676
rect 5626 9664 5632 9676
rect 5684 9664 5690 9716
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6454 9704 6460 9716
rect 6144 9676 6460 9704
rect 6144 9664 6150 9676
rect 6454 9664 6460 9676
rect 6512 9704 6518 9716
rect 6549 9707 6607 9713
rect 6549 9704 6561 9707
rect 6512 9676 6561 9704
rect 6512 9664 6518 9676
rect 6549 9673 6561 9676
rect 6595 9673 6607 9707
rect 6549 9667 6607 9673
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 6788 9676 7328 9704
rect 6788 9664 6794 9676
rect 6178 9636 6184 9648
rect 4448 9608 4568 9636
rect 5934 9608 6184 9636
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 2961 9571 3019 9577
rect 2961 9568 2973 9571
rect 2832 9540 2973 9568
rect 2832 9528 2838 9540
rect 2961 9537 2973 9540
rect 3007 9537 3019 9571
rect 2961 9531 3019 9537
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9568 3203 9571
rect 3326 9568 3332 9580
rect 3191 9540 3332 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2648 9472 2697 9500
rect 2648 9460 2654 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2976 9500 3004 9531
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 3476 9540 3525 9568
rect 3476 9528 3482 9540
rect 3513 9537 3525 9540
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 3660 9540 3801 9568
rect 3660 9528 3666 9540
rect 3789 9537 3801 9540
rect 3835 9568 3847 9571
rect 4154 9568 4160 9580
rect 3835 9540 4160 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4448 9577 4476 9608
rect 6178 9596 6184 9608
rect 6236 9596 6242 9648
rect 6362 9596 6368 9648
rect 6420 9596 6426 9648
rect 7300 9636 7328 9676
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 13998 9704 14004 9716
rect 8076 9676 14004 9704
rect 8076 9664 8082 9676
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 8113 9639 8171 9645
rect 8113 9636 8125 9639
rect 7300 9608 7604 9636
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4062 9500 4068 9512
rect 2976 9472 4068 9500
rect 2685 9463 2743 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 2866 9432 2872 9444
rect 2516 9404 2872 9432
rect 2409 9395 2467 9401
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9364 2835 9367
rect 3050 9364 3056 9376
rect 2823 9336 3056 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3326 9324 3332 9376
rect 3384 9324 3390 9376
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 4120 9336 4169 9364
rect 4120 9324 4126 9336
rect 4157 9333 4169 9336
rect 4203 9333 4215 9367
rect 4356 9364 4384 9531
rect 5994 9528 6000 9580
rect 6052 9568 6058 9580
rect 6270 9568 6276 9580
rect 6052 9540 6276 9568
rect 6052 9528 6058 9540
rect 6270 9528 6276 9540
rect 6328 9568 6334 9580
rect 7576 9577 7604 9608
rect 7668 9608 8125 9636
rect 7668 9580 7696 9608
rect 8113 9605 8125 9608
rect 8159 9605 8171 9639
rect 8113 9599 8171 9605
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 9401 9639 9459 9645
rect 9401 9636 9413 9639
rect 8996 9608 9413 9636
rect 8996 9596 9002 9608
rect 9401 9605 9413 9608
rect 9447 9605 9459 9639
rect 9401 9599 9459 9605
rect 9766 9596 9772 9648
rect 9824 9636 9830 9648
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9824 9608 9873 9636
rect 9824 9596 9830 9608
rect 9861 9605 9873 9608
rect 9907 9605 9919 9639
rect 9861 9599 9919 9605
rect 10318 9596 10324 9648
rect 10376 9596 10382 9648
rect 12066 9596 12072 9648
rect 12124 9636 12130 9648
rect 12621 9639 12679 9645
rect 12621 9636 12633 9639
rect 12124 9608 12633 9636
rect 12124 9596 12130 9608
rect 12621 9605 12633 9608
rect 12667 9605 12679 9639
rect 12621 9599 12679 9605
rect 13909 9639 13967 9645
rect 13909 9605 13921 9639
rect 13955 9636 13967 9639
rect 14274 9636 14280 9648
rect 13955 9608 14280 9636
rect 13955 9605 13967 9608
rect 13909 9599 13967 9605
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 6641 9571 6699 9577
rect 7469 9574 7527 9577
rect 6641 9568 6653 9571
rect 6328 9540 6653 9568
rect 6328 9528 6334 9540
rect 6641 9537 6653 9540
rect 6687 9568 6699 9571
rect 7392 9571 7527 9574
rect 7392 9568 7481 9571
rect 6687 9546 7481 9568
rect 6687 9540 7420 9546
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7469 9537 7481 9546
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7650 9528 7656 9580
rect 7708 9528 7714 9580
rect 8018 9568 8024 9580
rect 7760 9540 8024 9568
rect 4696 9503 4754 9509
rect 4696 9500 4708 9503
rect 4448 9472 4708 9500
rect 4448 9444 4476 9472
rect 4696 9469 4708 9472
rect 4742 9469 4754 9503
rect 4696 9463 4754 9469
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5902 9500 5908 9512
rect 5500 9472 5908 9500
rect 5500 9460 5506 9472
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 6512 9472 7389 9500
rect 6512 9460 6518 9472
rect 7377 9469 7389 9472
rect 7423 9500 7435 9503
rect 7760 9500 7788 9540
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 9033 9571 9091 9577
rect 9033 9568 9045 9571
rect 8266 9540 9045 9568
rect 8266 9512 8294 9540
rect 9033 9537 9045 9540
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 7423 9472 7788 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 7834 9460 7840 9512
rect 7892 9460 7898 9512
rect 8110 9500 8116 9512
rect 8036 9472 8116 9500
rect 4430 9392 4436 9444
rect 4488 9392 4494 9444
rect 8036 9432 8064 9472
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8202 9460 8208 9512
rect 8260 9472 8294 9512
rect 9232 9500 9260 9531
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9364 9540 9597 9568
rect 9364 9528 9370 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11572 9540 11989 9568
rect 11572 9528 11578 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 11977 9531 12035 9537
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12535 9571 12593 9577
rect 12535 9568 12547 9571
rect 12492 9540 12547 9568
rect 12492 9528 12498 9540
rect 12535 9537 12547 9540
rect 12581 9537 12593 9571
rect 12535 9531 12593 9537
rect 12710 9528 12716 9580
rect 12768 9528 12774 9580
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 12860 9540 13676 9568
rect 12860 9528 12866 9540
rect 11238 9500 11244 9512
rect 9232 9472 11244 9500
rect 8260 9460 8266 9472
rect 11238 9460 11244 9472
rect 11296 9500 11302 9512
rect 11609 9503 11667 9509
rect 11296 9472 11376 9500
rect 11296 9460 11302 9472
rect 9306 9432 9312 9444
rect 7760 9404 8064 9432
rect 8128 9404 9312 9432
rect 7760 9376 7788 9404
rect 5074 9364 5080 9376
rect 4356 9336 5080 9364
rect 4157 9327 4215 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 6178 9324 6184 9376
rect 6236 9324 6242 9376
rect 6917 9367 6975 9373
rect 6917 9333 6929 9367
rect 6963 9364 6975 9367
rect 7282 9364 7288 9376
rect 6963 9336 7288 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7742 9324 7748 9376
rect 7800 9324 7806 9376
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8128 9364 8156 9404
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 11348 9441 11376 9472
rect 11609 9469 11621 9503
rect 11655 9500 11667 9503
rect 13648 9500 13676 9540
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14369 9571 14427 9577
rect 14369 9568 14381 9571
rect 13780 9540 14381 9568
rect 13780 9528 13786 9540
rect 14369 9537 14381 9540
rect 14415 9568 14427 9571
rect 15286 9568 15292 9580
rect 14415 9540 15292 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 14182 9500 14188 9512
rect 11655 9472 13584 9500
rect 13648 9472 14188 9500
rect 11655 9469 11667 9472
rect 11609 9463 11667 9469
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9432 11391 9435
rect 12802 9432 12808 9444
rect 11379 9404 12808 9432
rect 11379 9401 11391 9404
rect 11333 9395 11391 9401
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 8076 9336 8156 9364
rect 8076 9324 8082 9336
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 8628 9336 8861 9364
rect 8628 9324 8634 9336
rect 8849 9333 8861 9336
rect 8895 9333 8907 9367
rect 8849 9327 8907 9333
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 10226 9364 10232 9376
rect 8996 9336 10232 9364
rect 8996 9324 9002 9336
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 12066 9364 12072 9376
rect 10376 9336 12072 9364
rect 10376 9324 10382 9336
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12710 9364 12716 9376
rect 12483 9336 12716 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12710 9324 12716 9336
rect 12768 9364 12774 9376
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 12768 9336 13001 9364
rect 12768 9324 12774 9336
rect 12989 9333 13001 9336
rect 13035 9364 13047 9367
rect 13262 9364 13268 9376
rect 13035 9336 13268 9364
rect 13035 9333 13047 9336
rect 12989 9327 13047 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 13412 9336 13461 9364
rect 13412 9324 13418 9336
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 13556 9364 13584 9472
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 13814 9364 13820 9376
rect 13556 9336 13820 9364
rect 13449 9327 13507 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 1104 9274 14812 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 14812 9274
rect 1104 9200 14812 9222
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2774 9160 2780 9172
rect 2280 9132 2780 9160
rect 2280 9120 2286 9132
rect 2774 9120 2780 9132
rect 2832 9120 2838 9172
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3970 9160 3976 9172
rect 3476 9132 3976 9160
rect 3476 9120 3482 9132
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 5718 9160 5724 9172
rect 5408 9132 5724 9160
rect 5408 9120 5414 9132
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 5905 9163 5963 9169
rect 5905 9129 5917 9163
rect 5951 9160 5963 9163
rect 10134 9160 10140 9172
rect 5951 9132 10140 9160
rect 5951 9129 5963 9132
rect 5905 9123 5963 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 10284 9132 13001 9160
rect 10284 9120 10290 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 4430 9092 4436 9104
rect 2455 9064 4436 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 5644 9064 5948 9092
rect 5445 9027 5503 9033
rect 5445 8993 5457 9027
rect 5491 9024 5503 9027
rect 5644 9024 5672 9064
rect 5920 9036 5948 9064
rect 7282 9052 7288 9104
rect 7340 9092 7346 9104
rect 8018 9092 8024 9104
rect 7340 9064 8024 9092
rect 7340 9052 7346 9064
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 9122 9092 9128 9104
rect 8904 9064 9128 9092
rect 8904 9052 8910 9064
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 9309 9095 9367 9101
rect 9309 9061 9321 9095
rect 9355 9061 9367 9095
rect 9309 9055 9367 9061
rect 5491 8996 5672 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 5718 8984 5724 9036
rect 5776 8984 5782 9036
rect 5902 8984 5908 9036
rect 5960 8984 5966 9036
rect 7466 9024 7472 9036
rect 6840 8996 7472 9024
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 4154 8956 4160 8968
rect 2271 8928 4160 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 5736 8928 5825 8956
rect 5736 8900 5764 8928
rect 5813 8925 5825 8928
rect 5859 8956 5871 8959
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 5859 8928 6377 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 6365 8925 6377 8928
rect 6411 8956 6423 8959
rect 6840 8956 6868 8996
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 8202 9024 8208 9036
rect 7800 8996 8208 9024
rect 7800 8984 7806 8996
rect 8202 8984 8208 8996
rect 8260 9024 8266 9036
rect 8570 9024 8576 9036
rect 8260 8996 8576 9024
rect 8260 8984 8266 8996
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 8662 8984 8668 9036
rect 8720 9024 8726 9036
rect 9324 9024 9352 9055
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 11701 9095 11759 9101
rect 11701 9092 11713 9095
rect 10744 9064 11713 9092
rect 10744 9052 10750 9064
rect 11701 9061 11713 9064
rect 11747 9092 11759 9095
rect 12434 9092 12440 9104
rect 11747 9064 12440 9092
rect 11747 9061 11759 9064
rect 11701 9055 11759 9061
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 8720 8996 8984 9024
rect 9324 8996 12434 9024
rect 8720 8984 8726 8996
rect 8956 8968 8984 8996
rect 6411 8928 6868 8956
rect 6411 8925 6423 8928
rect 6365 8919 6423 8925
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 8754 8956 8760 8968
rect 6972 8928 8760 8956
rect 6972 8916 6978 8928
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 4982 8848 4988 8900
rect 5040 8848 5046 8900
rect 5718 8848 5724 8900
rect 5776 8848 5782 8900
rect 6270 8848 6276 8900
rect 6328 8888 6334 8900
rect 7009 8891 7067 8897
rect 7009 8888 7021 8891
rect 6328 8860 7021 8888
rect 6328 8848 6334 8860
rect 7009 8857 7021 8860
rect 7055 8857 7067 8891
rect 7009 8851 7067 8857
rect 7834 8848 7840 8900
rect 7892 8888 7898 8900
rect 8570 8888 8576 8900
rect 7892 8860 8576 8888
rect 7892 8848 7898 8860
rect 8570 8848 8576 8860
rect 8628 8848 8634 8900
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 9416 8888 9444 8919
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11572 8928 11621 8956
rect 11572 8916 11578 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11793 8959 11851 8965
rect 11793 8925 11805 8959
rect 11839 8956 11851 8959
rect 11882 8956 11888 8968
rect 11839 8928 11888 8956
rect 11839 8925 11851 8928
rect 11793 8919 11851 8925
rect 11882 8916 11888 8928
rect 11940 8956 11946 8968
rect 12250 8956 12256 8968
rect 11940 8928 12256 8956
rect 11940 8916 11946 8928
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 8720 8860 9444 8888
rect 8720 8848 8726 8860
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 3142 8820 3148 8832
rect 2648 8792 3148 8820
rect 2648 8780 2654 8792
rect 3142 8780 3148 8792
rect 3200 8820 3206 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 3200 8792 3433 8820
rect 3200 8780 3206 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3973 8823 4031 8829
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 4430 8820 4436 8832
rect 4019 8792 4436 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 7650 8820 7656 8832
rect 4764 8792 7656 8820
rect 4764 8780 4770 8792
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8297 8823 8355 8829
rect 8297 8820 8309 8823
rect 8260 8792 8309 8820
rect 8260 8780 8266 8792
rect 8297 8789 8309 8792
rect 8343 8789 8355 8823
rect 9416 8820 9444 8860
rect 9674 8848 9680 8900
rect 9732 8848 9738 8900
rect 10134 8848 10140 8900
rect 10192 8848 10198 8900
rect 12406 8888 12434 8996
rect 13004 8956 13032 9123
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 13004 8928 13185 8956
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13446 8956 13452 8968
rect 13403 8928 13452 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13446 8916 13452 8928
rect 13504 8956 13510 8968
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 13504 8928 13645 8956
rect 13504 8916 13510 8928
rect 13633 8925 13645 8928
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 12986 8888 12992 8900
rect 12406 8860 12992 8888
rect 12986 8848 12992 8860
rect 13044 8848 13050 8900
rect 9766 8820 9772 8832
rect 9416 8792 9772 8820
rect 8297 8783 8355 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 13265 8823 13323 8829
rect 13265 8789 13277 8823
rect 13311 8820 13323 8823
rect 13538 8820 13544 8832
rect 13311 8792 13544 8820
rect 13311 8789 13323 8792
rect 13265 8783 13323 8789
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 14458 8780 14464 8832
rect 14516 8780 14522 8832
rect 1104 8730 14812 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 14812 8730
rect 1104 8656 14812 8678
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5902 8616 5908 8628
rect 5592 8588 5908 8616
rect 5592 8576 5598 8588
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 9674 8616 9680 8628
rect 6052 8588 9680 8616
rect 6052 8576 6058 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10870 8616 10876 8628
rect 10520 8588 10876 8616
rect 2314 8508 2320 8560
rect 2372 8548 2378 8560
rect 2372 8520 4278 8548
rect 2372 8508 2378 8520
rect 6086 8508 6092 8560
rect 6144 8548 6150 8560
rect 8018 8548 8024 8560
rect 6144 8520 8024 8548
rect 6144 8508 6150 8520
rect 8018 8508 8024 8520
rect 8076 8508 8082 8560
rect 9030 8548 9036 8560
rect 8266 8520 9036 8548
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 5994 8480 6000 8492
rect 5767 8452 6000 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 3050 8372 3056 8424
rect 3108 8412 3114 8424
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 3108 8384 3525 8412
rect 3108 8372 3114 8384
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 3513 8375 3571 8381
rect 3786 8372 3792 8424
rect 3844 8372 3850 8424
rect 5166 8372 5172 8424
rect 5224 8412 5230 8424
rect 5534 8412 5540 8424
rect 5224 8384 5540 8412
rect 5224 8372 5230 8384
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 6656 8412 6684 8443
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 8266 8480 8294 8520
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 10520 8548 10548 8588
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 11020 8588 11253 8616
rect 11020 8576 11026 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 11241 8579 11299 8585
rect 10166 8520 10548 8548
rect 6788 8452 8294 8480
rect 6788 8440 6794 8452
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 10226 8440 10232 8492
rect 10284 8480 10290 8492
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 10284 8452 10517 8480
rect 10284 8440 10290 8452
rect 10505 8449 10517 8452
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 11256 8480 11284 8579
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11664 8588 12081 8616
rect 11664 8576 11670 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 12069 8579 12127 8585
rect 12342 8576 12348 8628
rect 12400 8616 12406 8628
rect 13722 8616 13728 8628
rect 12400 8588 13728 8616
rect 12400 8576 12406 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 13906 8576 13912 8628
rect 13964 8576 13970 8628
rect 14090 8576 14096 8628
rect 14148 8576 14154 8628
rect 15194 8616 15200 8628
rect 14384 8588 15200 8616
rect 11330 8508 11336 8560
rect 11388 8548 11394 8560
rect 11388 8520 12296 8548
rect 11388 8508 11394 8520
rect 12268 8489 12296 8520
rect 12434 8508 12440 8560
rect 12492 8548 12498 8560
rect 14245 8551 14303 8557
rect 14245 8548 14257 8551
rect 12492 8520 14257 8548
rect 12492 8508 12498 8520
rect 14245 8517 14257 8520
rect 14291 8517 14303 8551
rect 14245 8511 14303 8517
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11256 8452 11529 8480
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 13906 8440 13912 8492
rect 13964 8480 13970 8492
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 13964 8452 14013 8480
rect 13964 8440 13970 8452
rect 14001 8449 14013 8452
rect 14047 8480 14059 8483
rect 14384 8480 14412 8588
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 14461 8551 14519 8557
rect 14461 8517 14473 8551
rect 14507 8517 14519 8551
rect 14461 8511 14519 8517
rect 14047 8452 14412 8480
rect 14047 8449 14059 8452
rect 14001 8443 14059 8449
rect 7926 8412 7932 8424
rect 6656 8384 7932 8412
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8680 8384 8953 8412
rect 8680 8356 8708 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 10410 8372 10416 8424
rect 10468 8372 10474 8424
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 11146 8412 11152 8424
rect 10836 8384 11152 8412
rect 10836 8372 10842 8384
rect 11146 8372 11152 8384
rect 11204 8372 11210 8424
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 11974 8412 11980 8424
rect 11839 8384 11980 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 11974 8372 11980 8384
rect 12032 8412 12038 8424
rect 12032 8384 12388 8412
rect 12032 8372 12038 8384
rect 5258 8304 5264 8356
rect 5316 8304 5322 8356
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 6457 8347 6515 8353
rect 6457 8344 6469 8347
rect 5500 8316 6469 8344
rect 5500 8304 5506 8316
rect 6457 8313 6469 8316
rect 6503 8344 6515 8347
rect 7558 8344 7564 8356
rect 6503 8316 7564 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 8662 8304 8668 8356
rect 8720 8304 8726 8356
rect 9950 8304 9956 8356
rect 10008 8344 10014 8356
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 10008 8316 10885 8344
rect 10008 8304 10014 8316
rect 10873 8313 10885 8316
rect 10919 8313 10931 8347
rect 10873 8307 10931 8313
rect 1854 8236 1860 8288
rect 1912 8276 1918 8288
rect 2222 8276 2228 8288
rect 1912 8248 2228 8276
rect 1912 8236 1918 8248
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 3421 8279 3479 8285
rect 3421 8245 3433 8279
rect 3467 8276 3479 8279
rect 4430 8276 4436 8288
rect 3467 8248 4436 8276
rect 3467 8245 3479 8248
rect 3421 8239 3479 8245
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5718 8276 5724 8288
rect 4948 8248 5724 8276
rect 4948 8236 4954 8248
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 6089 8279 6147 8285
rect 6089 8245 6101 8279
rect 6135 8276 6147 8279
rect 7190 8276 7196 8288
rect 6135 8248 7196 8276
rect 6135 8245 6147 8248
rect 6089 8239 6147 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 10226 8276 10232 8288
rect 9088 8248 10232 8276
rect 9088 8236 9094 8248
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 12360 8276 12388 8384
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 12492 8384 13369 8412
rect 12492 8372 12498 8384
rect 13357 8381 13369 8384
rect 13403 8412 13415 8415
rect 14476 8412 14504 8511
rect 13403 8384 14504 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 13446 8344 13452 8356
rect 12584 8316 13452 8344
rect 12584 8304 12590 8316
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 13725 8279 13783 8285
rect 13725 8276 13737 8279
rect 12360 8248 13737 8276
rect 13725 8245 13737 8248
rect 13771 8276 13783 8279
rect 13906 8276 13912 8288
rect 13771 8248 13912 8276
rect 13771 8245 13783 8248
rect 13725 8239 13783 8245
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 14277 8279 14335 8285
rect 14277 8245 14289 8279
rect 14323 8276 14335 8279
rect 14734 8276 14740 8288
rect 14323 8248 14740 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 1104 8186 14812 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 14812 8186
rect 1104 8112 14812 8134
rect 4522 8032 4528 8084
rect 4580 8032 4586 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 6917 8075 6975 8081
rect 5132 8044 6776 8072
rect 5132 8032 5138 8044
rect 6638 8004 6644 8016
rect 4816 7976 6644 8004
rect 3528 7908 4200 7936
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2222 7868 2228 7880
rect 1912 7840 2228 7868
rect 1912 7828 1918 7840
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2314 7828 2320 7880
rect 2372 7868 2378 7880
rect 2409 7871 2467 7877
rect 2409 7868 2421 7871
rect 2372 7840 2421 7868
rect 2372 7828 2378 7840
rect 2409 7837 2421 7840
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7769 3295 7803
rect 3237 7763 3295 7769
rect 2314 7692 2320 7744
rect 2372 7692 2378 7744
rect 3252 7732 3280 7763
rect 3528 7732 3556 7908
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 3752 7840 3893 7868
rect 3752 7828 3758 7840
rect 3881 7837 3893 7840
rect 3927 7837 3939 7871
rect 3881 7831 3939 7837
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4172 7877 4200 7908
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 4028 7840 4077 7868
rect 4028 7828 4034 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4339 7871 4397 7877
rect 4339 7837 4351 7871
rect 4385 7868 4397 7871
rect 4430 7868 4436 7880
rect 4385 7840 4436 7868
rect 4385 7837 4397 7840
rect 4339 7831 4397 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 4816 7877 4844 7976
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 6748 8004 6776 8044
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 9582 8072 9588 8084
rect 6963 8044 9588 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 10042 8072 10048 8084
rect 9824 8044 10048 8072
rect 9824 8032 9830 8044
rect 10042 8032 10048 8044
rect 10100 8072 10106 8084
rect 10689 8075 10747 8081
rect 10689 8072 10701 8075
rect 10100 8044 10701 8072
rect 10100 8032 10106 8044
rect 10689 8041 10701 8044
rect 10735 8072 10747 8075
rect 11057 8075 11115 8081
rect 11057 8072 11069 8075
rect 10735 8044 11069 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 11057 8041 11069 8044
rect 11103 8041 11115 8075
rect 11057 8035 11115 8041
rect 9030 8004 9036 8016
rect 6748 7976 9036 8004
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9122 7964 9128 8016
rect 9180 8004 9186 8016
rect 10873 8007 10931 8013
rect 10873 8004 10885 8007
rect 9180 7976 10885 8004
rect 9180 7964 9186 7976
rect 10873 7973 10885 7976
rect 10919 7973 10931 8007
rect 11072 8004 11100 8035
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 14274 8072 14280 8084
rect 11940 8044 14280 8072
rect 11940 8032 11946 8044
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 12434 8004 12440 8016
rect 11072 7976 12440 8004
rect 10873 7967 10931 7973
rect 12434 7964 12440 7976
rect 12492 7964 12498 8016
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 5224 7908 5457 7936
rect 5224 7896 5230 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 6086 7936 6092 7948
rect 5776 7908 6092 7936
rect 5776 7896 5782 7908
rect 6086 7896 6092 7908
rect 6144 7936 6150 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 6144 7908 6285 7936
rect 6144 7896 6150 7908
rect 6273 7905 6285 7908
rect 6319 7936 6331 7939
rect 10042 7936 10048 7948
rect 6319 7908 10048 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4580 7840 4813 7868
rect 4580 7828 4586 7840
rect 4801 7837 4813 7840
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 5074 7828 5080 7880
rect 5132 7828 5138 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5350 7868 5356 7880
rect 5307 7840 5356 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7868 5595 7871
rect 6178 7868 6184 7880
rect 5583 7840 6184 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6472 7840 6745 7868
rect 6472 7812 6500 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7098 7868 7104 7880
rect 6963 7840 7104 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7098 7828 7104 7840
rect 7156 7868 7162 7880
rect 7558 7868 7564 7880
rect 7156 7840 7564 7868
rect 7156 7828 7162 7840
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 9582 7868 9588 7880
rect 7892 7840 9588 7868
rect 7892 7828 7898 7840
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 10192 7840 11437 7868
rect 10192 7828 10198 7840
rect 11425 7837 11437 7840
rect 11471 7868 11483 7871
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11471 7840 12081 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 3605 7803 3663 7809
rect 3605 7769 3617 7803
rect 3651 7800 3663 7803
rect 4617 7803 4675 7809
rect 4617 7800 4629 7803
rect 3651 7772 4629 7800
rect 3651 7769 3663 7772
rect 3605 7763 3663 7769
rect 4617 7769 4629 7772
rect 4663 7800 4675 7803
rect 4706 7800 4712 7812
rect 4663 7772 4712 7800
rect 4663 7769 4675 7772
rect 4617 7763 4675 7769
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 4985 7803 5043 7809
rect 4985 7769 4997 7803
rect 5031 7769 5043 7803
rect 5994 7800 6000 7812
rect 4985 7763 5043 7769
rect 5184 7772 6000 7800
rect 3694 7732 3700 7744
rect 3252 7704 3700 7732
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 3970 7692 3976 7744
rect 4028 7692 4034 7744
rect 5000 7732 5028 7763
rect 5184 7732 5212 7772
rect 5994 7760 6000 7772
rect 6052 7760 6058 7812
rect 6454 7760 6460 7812
rect 6512 7760 6518 7812
rect 6638 7760 6644 7812
rect 6696 7800 6702 7812
rect 13446 7800 13452 7812
rect 6696 7772 13452 7800
rect 6696 7760 6702 7772
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 5000 7704 5212 7732
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7732 5319 7735
rect 5350 7732 5356 7744
rect 5307 7704 5356 7732
rect 5307 7701 5319 7704
rect 5261 7695 5319 7701
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 6178 7732 6184 7744
rect 5500 7704 6184 7732
rect 5500 7692 5506 7704
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6472 7732 6500 7760
rect 7193 7735 7251 7741
rect 7193 7732 7205 7735
rect 6472 7704 7205 7732
rect 7193 7701 7205 7704
rect 7239 7732 7251 7735
rect 10502 7732 10508 7744
rect 7239 7704 10508 7732
rect 7239 7701 7251 7704
rect 7193 7695 7251 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 11020 7704 11069 7732
rect 11020 7692 11026 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 11701 7735 11759 7741
rect 11701 7732 11713 7735
rect 11204 7704 11713 7732
rect 11204 7692 11210 7704
rect 11701 7701 11713 7704
rect 11747 7732 11759 7735
rect 11882 7732 11888 7744
rect 11747 7704 11888 7732
rect 11747 7701 11759 7704
rect 11701 7695 11759 7701
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 12434 7692 12440 7744
rect 12492 7732 12498 7744
rect 12618 7732 12624 7744
rect 12492 7704 12624 7732
rect 12492 7692 12498 7704
rect 12618 7692 12624 7704
rect 12676 7732 12682 7744
rect 13817 7735 13875 7741
rect 13817 7732 13829 7735
rect 12676 7704 13829 7732
rect 12676 7692 12682 7704
rect 13817 7701 13829 7704
rect 13863 7701 13875 7735
rect 13817 7695 13875 7701
rect 14458 7692 14464 7744
rect 14516 7692 14522 7744
rect 1104 7642 14812 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 14812 7642
rect 1104 7568 14812 7590
rect 842 7488 848 7540
rect 900 7528 906 7540
rect 2409 7531 2467 7537
rect 2409 7528 2421 7531
rect 900 7500 2421 7528
rect 900 7488 906 7500
rect 2409 7497 2421 7500
rect 2455 7497 2467 7531
rect 2409 7491 2467 7497
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 2958 7528 2964 7540
rect 2648 7500 2964 7528
rect 2648 7488 2654 7500
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 4062 7488 4068 7540
rect 4120 7488 4126 7540
rect 4338 7488 4344 7540
rect 4396 7488 4402 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 6454 7528 6460 7540
rect 5500 7500 6460 7528
rect 5500 7488 5506 7500
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6546 7488 6552 7540
rect 6604 7488 6610 7540
rect 6730 7488 6736 7540
rect 6788 7488 6794 7540
rect 6822 7488 6828 7540
rect 6880 7488 6886 7540
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 7374 7528 7380 7540
rect 7331 7500 7380 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10594 7528 10600 7540
rect 10100 7500 10600 7528
rect 10100 7488 10106 7500
rect 1762 7460 1768 7472
rect 1412 7432 1768 7460
rect 658 7352 664 7404
rect 716 7392 722 7404
rect 842 7392 848 7404
rect 716 7364 848 7392
rect 716 7352 722 7364
rect 842 7352 848 7364
rect 900 7352 906 7404
rect 1412 7401 1440 7432
rect 1762 7420 1768 7432
rect 1820 7420 1826 7472
rect 3418 7420 3424 7472
rect 3476 7420 3482 7472
rect 3881 7463 3939 7469
rect 3881 7429 3893 7463
rect 3927 7460 3939 7463
rect 4080 7460 4108 7488
rect 3927 7432 4108 7460
rect 4356 7460 4384 7488
rect 4525 7463 4583 7469
rect 4525 7460 4537 7463
rect 4356 7432 4537 7460
rect 3927 7429 3939 7432
rect 3881 7423 3939 7429
rect 4525 7429 4537 7432
rect 4571 7429 4583 7463
rect 5902 7460 5908 7472
rect 5750 7432 5908 7460
rect 4525 7423 4583 7429
rect 5902 7420 5908 7432
rect 5960 7420 5966 7472
rect 6564 7460 6592 7488
rect 7653 7463 7711 7469
rect 7653 7460 7665 7463
rect 6564 7432 6868 7460
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 2222 7392 2228 7404
rect 1627 7364 2228 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 2498 7284 2504 7336
rect 2556 7324 2562 7336
rect 2682 7324 2688 7336
rect 2556 7296 2688 7324
rect 2556 7284 2562 7296
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4249 7327 4307 7333
rect 4249 7324 4261 7327
rect 4212 7296 4261 7324
rect 4212 7284 4218 7296
rect 4249 7293 4261 7296
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 6380 7324 6408 7355
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6840 7401 6868 7432
rect 7116 7432 7665 7460
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6512 7364 6561 7392
rect 6512 7352 6518 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 7116 7392 7144 7432
rect 7653 7429 7665 7432
rect 7699 7460 7711 7463
rect 10134 7460 10140 7472
rect 7699 7432 10140 7460
rect 7699 7429 7711 7432
rect 7653 7423 7711 7429
rect 10134 7420 10140 7432
rect 10192 7420 10198 7472
rect 10336 7469 10364 7500
rect 10594 7488 10600 7500
rect 10652 7528 10658 7540
rect 10652 7500 13124 7528
rect 10652 7488 10658 7500
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7429 10379 7463
rect 10321 7423 10379 7429
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 10781 7463 10839 7469
rect 10781 7460 10793 7463
rect 10560 7432 10793 7460
rect 10560 7420 10566 7432
rect 10781 7429 10793 7432
rect 10827 7429 10839 7463
rect 10781 7423 10839 7429
rect 11790 7420 11796 7472
rect 11848 7420 11854 7472
rect 6825 7355 6883 7361
rect 6932 7364 7144 7392
rect 6932 7324 6960 7364
rect 7190 7352 7196 7404
rect 7248 7352 7254 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 8021 7395 8079 7401
rect 7423 7364 7457 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 8021 7361 8033 7395
rect 8067 7392 8079 7395
rect 9858 7392 9864 7404
rect 8067 7364 9864 7392
rect 8067 7361 8079 7364
rect 8021 7355 8079 7361
rect 4672 7296 6960 7324
rect 4672 7284 4678 7296
rect 7098 7284 7104 7336
rect 7156 7324 7162 7336
rect 7392 7324 7420 7355
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 10100 7364 10241 7392
rect 10100 7352 10106 7364
rect 10229 7361 10241 7364
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 11146 7352 11152 7404
rect 11204 7352 11210 7404
rect 11238 7352 11244 7404
rect 11296 7392 11302 7404
rect 11333 7395 11391 7401
rect 11333 7392 11345 7395
rect 11296 7364 11345 7392
rect 11296 7352 11302 7364
rect 11333 7361 11345 7364
rect 11379 7361 11391 7395
rect 11333 7355 11391 7361
rect 12894 7352 12900 7404
rect 12952 7352 12958 7404
rect 13096 7392 13124 7500
rect 13446 7488 13452 7540
rect 13504 7488 13510 7540
rect 13906 7488 13912 7540
rect 13964 7488 13970 7540
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 14369 7531 14427 7537
rect 14369 7528 14381 7531
rect 14240 7500 14381 7528
rect 14240 7488 14246 7500
rect 14369 7497 14381 7500
rect 14415 7497 14427 7531
rect 14369 7491 14427 7497
rect 13924 7460 13952 7488
rect 13556 7432 14412 7460
rect 13446 7392 13452 7404
rect 13096 7364 13452 7392
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13556 7401 13584 7432
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13964 7364 14013 7392
rect 13964 7352 13970 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 7466 7324 7472 7336
rect 7156 7296 7472 7324
rect 7156 7284 7162 7296
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 11422 7284 11428 7336
rect 11480 7324 11486 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 11480 7296 11529 7324
rect 11480 7284 11486 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 11790 7284 11796 7336
rect 11848 7324 11854 7336
rect 12342 7324 12348 7336
rect 11848 7296 12348 7324
rect 11848 7284 11854 7296
rect 12342 7284 12348 7296
rect 12400 7324 12406 7336
rect 14292 7324 14320 7355
rect 12400 7296 14320 7324
rect 12400 7284 12406 7296
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 6086 7256 6092 7268
rect 5592 7228 6092 7256
rect 5592 7216 5598 7228
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 6917 7259 6975 7265
rect 6917 7225 6929 7259
rect 6963 7256 6975 7259
rect 7282 7256 7288 7268
rect 6963 7228 7288 7256
rect 6963 7225 6975 7228
rect 6917 7219 6975 7225
rect 7282 7216 7288 7228
rect 7340 7216 7346 7268
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 7929 7259 7987 7265
rect 7929 7256 7941 7259
rect 7432 7228 7941 7256
rect 7432 7216 7438 7228
rect 7929 7225 7941 7228
rect 7975 7225 7987 7259
rect 7929 7219 7987 7225
rect 12802 7216 12808 7268
rect 12860 7256 12866 7268
rect 13265 7259 13323 7265
rect 13265 7256 13277 7259
rect 12860 7228 13277 7256
rect 12860 7216 12866 7228
rect 13265 7225 13277 7228
rect 13311 7256 13323 7259
rect 13630 7256 13636 7268
rect 13311 7228 13636 7256
rect 13311 7225 13323 7228
rect 13265 7219 13323 7225
rect 13630 7216 13636 7228
rect 13688 7216 13694 7268
rect 13909 7259 13967 7265
rect 13909 7225 13921 7259
rect 13955 7256 13967 7259
rect 14384 7256 14412 7432
rect 14642 7256 14648 7268
rect 13955 7228 14648 7256
rect 13955 7225 13967 7228
rect 13909 7219 13967 7225
rect 14642 7216 14648 7228
rect 14700 7216 14706 7268
rect 1489 7191 1547 7197
rect 1489 7157 1501 7191
rect 1535 7188 1547 7191
rect 2314 7188 2320 7200
rect 1535 7160 2320 7188
rect 1535 7157 1547 7160
rect 1489 7151 1547 7157
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 5552 7188 5580 7216
rect 3752 7160 5580 7188
rect 5997 7191 6055 7197
rect 3752 7148 3758 7160
rect 5997 7157 6009 7191
rect 6043 7188 6055 7191
rect 8478 7188 8484 7200
rect 6043 7160 8484 7188
rect 6043 7157 6055 7160
rect 5997 7151 6055 7157
rect 8478 7148 8484 7160
rect 8536 7188 8542 7200
rect 8662 7188 8668 7200
rect 8536 7160 8668 7188
rect 8536 7148 8542 7160
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10229 7191 10287 7197
rect 10229 7188 10241 7191
rect 10192 7160 10241 7188
rect 10192 7148 10198 7160
rect 10229 7157 10241 7160
rect 10275 7157 10287 7191
rect 10229 7151 10287 7157
rect 11241 7191 11299 7197
rect 11241 7157 11253 7191
rect 11287 7188 11299 7191
rect 12250 7188 12256 7200
rect 11287 7160 12256 7188
rect 11287 7157 11299 7160
rect 11241 7151 11299 7157
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 14182 7148 14188 7200
rect 14240 7148 14246 7200
rect 1104 7098 14812 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 14812 7098
rect 1104 7024 14812 7046
rect 2869 6987 2927 6993
rect 2869 6953 2881 6987
rect 2915 6984 2927 6987
rect 2958 6984 2964 6996
rect 2915 6956 2964 6984
rect 2915 6953 2927 6956
rect 2869 6947 2927 6953
rect 2958 6944 2964 6956
rect 3016 6984 3022 6996
rect 4890 6984 4896 6996
rect 3016 6956 4896 6984
rect 3016 6944 3022 6956
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5077 6987 5135 6993
rect 5077 6984 5089 6987
rect 5040 6956 5089 6984
rect 5040 6944 5046 6956
rect 5077 6953 5089 6956
rect 5123 6953 5135 6987
rect 5077 6947 5135 6953
rect 750 6876 756 6928
rect 808 6916 814 6928
rect 808 6888 3188 6916
rect 808 6876 814 6888
rect 3050 6808 3056 6860
rect 3108 6808 3114 6860
rect 3160 6848 3188 6888
rect 4709 6851 4767 6857
rect 4709 6848 4721 6851
rect 3160 6820 4721 6848
rect 4709 6817 4721 6820
rect 4755 6817 4767 6851
rect 5092 6848 5120 6947
rect 6454 6944 6460 6996
rect 6512 6984 6518 6996
rect 9490 6984 9496 6996
rect 6512 6956 9496 6984
rect 6512 6944 6518 6956
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9640 6944 9674 6984
rect 11422 6944 11428 6996
rect 11480 6944 11486 6996
rect 12424 6987 12482 6993
rect 12424 6953 12436 6987
rect 12470 6984 12482 6987
rect 14458 6984 14464 6996
rect 12470 6956 14464 6984
rect 12470 6953 12482 6956
rect 12424 6947 12482 6953
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 5534 6876 5540 6928
rect 5592 6916 5598 6928
rect 5592 6888 6056 6916
rect 5592 6876 5598 6888
rect 5442 6848 5448 6860
rect 5092 6820 5448 6848
rect 4709 6811 4767 6817
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 6028 6848 6056 6888
rect 6086 6876 6092 6928
rect 6144 6916 6150 6928
rect 8018 6916 8024 6928
rect 6144 6888 8024 6916
rect 6144 6876 6150 6888
rect 8018 6876 8024 6888
rect 8076 6876 8082 6928
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 8260 6888 9536 6916
rect 8260 6876 8266 6888
rect 5500 6820 5948 6848
rect 6028 6820 6500 6848
rect 5500 6808 5506 6820
rect 2958 6740 2964 6792
rect 3016 6740 3022 6792
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3660 6752 3801 6780
rect 3660 6740 3666 6752
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3936 6752 4169 6780
rect 3936 6740 3942 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4246 6740 4252 6792
rect 4304 6789 4310 6792
rect 4304 6783 4332 6789
rect 4320 6749 4332 6783
rect 4304 6743 4332 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4304 6740 4310 6743
rect 4632 6712 4660 6743
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4948 6752 5273 6780
rect 4948 6740 4954 6752
rect 5261 6749 5273 6752
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5920 6789 5948 6820
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6472 6780 6500 6820
rect 9122 6808 9128 6860
rect 9180 6808 9186 6860
rect 6472 6752 8708 6780
rect 6454 6712 6460 6724
rect 3620 6684 6460 6712
rect 3620 6653 3648 6684
rect 3896 6656 3924 6684
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 7745 6715 7803 6721
rect 7745 6681 7757 6715
rect 7791 6712 7803 6715
rect 8202 6712 8208 6724
rect 7791 6684 8208 6712
rect 7791 6681 7803 6684
rect 7745 6675 7803 6681
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 8680 6712 8708 6752
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 8812 6752 9229 6780
rect 8812 6740 8818 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9122 6712 9128 6724
rect 8680 6684 9128 6712
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 9508 6712 9536 6888
rect 9646 6848 9674 6944
rect 11882 6848 11888 6860
rect 9646 6820 11888 6848
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 13909 6851 13967 6857
rect 12492 6820 13676 6848
rect 12492 6808 12498 6820
rect 11422 6740 11428 6792
rect 11480 6780 11486 6792
rect 12158 6780 12164 6792
rect 11480 6752 12164 6780
rect 11480 6740 11486 6752
rect 12158 6740 12164 6752
rect 12216 6740 12222 6792
rect 13648 6780 13676 6820
rect 13909 6817 13921 6851
rect 13955 6848 13967 6851
rect 15102 6848 15108 6860
rect 13955 6820 15108 6848
rect 13955 6817 13967 6820
rect 13909 6811 13967 6817
rect 15102 6808 15108 6820
rect 15160 6808 15166 6860
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13648 6752 14105 6780
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 10137 6715 10195 6721
rect 10137 6712 10149 6715
rect 9508 6684 10149 6712
rect 10137 6681 10149 6684
rect 10183 6681 10195 6715
rect 10137 6675 10195 6681
rect 11698 6672 11704 6724
rect 11756 6712 11762 6724
rect 11756 6684 12926 6712
rect 11756 6672 11762 6684
rect 3605 6647 3663 6653
rect 3605 6613 3617 6647
rect 3651 6613 3663 6647
rect 3605 6607 3663 6613
rect 3878 6604 3884 6656
rect 3936 6604 3942 6656
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6644 4123 6647
rect 4338 6644 4344 6656
rect 4111 6616 4344 6644
rect 4111 6613 4123 6616
rect 4065 6607 4123 6613
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 4430 6604 4436 6656
rect 4488 6604 4494 6656
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 4706 6644 4712 6656
rect 4580 6616 4712 6644
rect 4580 6604 4586 6616
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 5442 6604 5448 6656
rect 5500 6604 5506 6656
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 5626 6644 5632 6656
rect 5583 6616 5632 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7926 6644 7932 6656
rect 7340 6616 7932 6644
rect 7340 6604 7346 6616
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 9582 6604 9588 6656
rect 9640 6604 9646 6656
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 14185 6647 14243 6653
rect 14185 6644 14197 6647
rect 10928 6616 14197 6644
rect 10928 6604 10934 6616
rect 14185 6613 14197 6616
rect 14231 6613 14243 6647
rect 14185 6607 14243 6613
rect 1104 6554 14812 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 14812 6554
rect 1104 6480 14812 6502
rect 3513 6443 3571 6449
rect 3513 6409 3525 6443
rect 3559 6440 3571 6443
rect 3602 6440 3608 6452
rect 3559 6412 3608 6440
rect 3559 6409 3571 6412
rect 3513 6403 3571 6409
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4212 6412 5580 6440
rect 4212 6400 4218 6412
rect 3878 6332 3884 6384
rect 3936 6372 3942 6384
rect 5077 6375 5135 6381
rect 5077 6372 5089 6375
rect 3936 6344 5089 6372
rect 3936 6332 3942 6344
rect 5077 6341 5089 6344
rect 5123 6341 5135 6375
rect 5077 6335 5135 6341
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 4304 6276 4353 6304
rect 4304 6264 4310 6276
rect 4341 6273 4353 6276
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 5258 6304 5264 6316
rect 4764 6276 5264 6304
rect 4764 6264 4770 6276
rect 5258 6264 5264 6276
rect 5316 6304 5322 6316
rect 5552 6313 5580 6412
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 6013 6443 6071 6449
rect 6013 6440 6025 6443
rect 5684 6412 6025 6440
rect 5684 6400 5690 6412
rect 6013 6409 6025 6412
rect 6059 6409 6071 6443
rect 6013 6403 6071 6409
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 6880 6412 10364 6440
rect 6880 6400 6886 6412
rect 5718 6332 5724 6384
rect 5776 6372 5782 6384
rect 5813 6375 5871 6381
rect 5813 6372 5825 6375
rect 5776 6344 5825 6372
rect 5776 6332 5782 6344
rect 5813 6341 5825 6344
rect 5859 6372 5871 6375
rect 5902 6372 5908 6384
rect 5859 6344 5908 6372
rect 5859 6341 5871 6344
rect 5813 6335 5871 6341
rect 5902 6332 5908 6344
rect 5960 6332 5966 6384
rect 6028 6344 6868 6372
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 5316 6276 5457 6304
rect 5316 6264 5322 6276
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5626 6304 5632 6316
rect 5583 6276 5632 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 6028 6304 6056 6344
rect 5828 6276 6056 6304
rect 4522 6196 4528 6248
rect 4580 6236 4586 6248
rect 4801 6239 4859 6245
rect 4801 6236 4813 6239
rect 4580 6208 4813 6236
rect 4580 6196 4586 6208
rect 4801 6205 4813 6208
rect 4847 6236 4859 6239
rect 5828 6236 5856 6276
rect 6454 6264 6460 6316
rect 6512 6264 6518 6316
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 4847 6208 5856 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 6748 6236 6776 6267
rect 6840 6248 6868 6344
rect 7466 6332 7472 6384
rect 7524 6372 7530 6384
rect 7561 6375 7619 6381
rect 7561 6372 7573 6375
rect 7524 6344 7573 6372
rect 7524 6332 7530 6344
rect 7561 6341 7573 6344
rect 7607 6341 7619 6375
rect 7561 6335 7619 6341
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 8754 6372 8760 6384
rect 7708 6344 8760 6372
rect 7708 6332 7714 6344
rect 8754 6332 8760 6344
rect 8812 6372 8818 6384
rect 9582 6372 9588 6384
rect 8812 6344 9588 6372
rect 8812 6332 8818 6344
rect 9582 6332 9588 6344
rect 9640 6332 9646 6384
rect 10226 6332 10232 6384
rect 10284 6332 10290 6384
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7098 6304 7104 6316
rect 6963 6276 7104 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 10336 6313 10364 6412
rect 11790 6400 11796 6452
rect 11848 6440 11854 6452
rect 11977 6443 12035 6449
rect 11977 6440 11989 6443
rect 11848 6412 11989 6440
rect 11848 6400 11854 6412
rect 11977 6409 11989 6412
rect 12023 6409 12035 6443
rect 11977 6403 12035 6409
rect 13446 6400 13452 6452
rect 13504 6440 13510 6452
rect 13504 6412 14320 6440
rect 13504 6400 13510 6412
rect 10410 6332 10416 6384
rect 10468 6372 10474 6384
rect 10689 6375 10747 6381
rect 10689 6372 10701 6375
rect 10468 6344 10701 6372
rect 10468 6332 10474 6344
rect 10689 6341 10701 6344
rect 10735 6341 10747 6375
rect 12526 6372 12532 6384
rect 10689 6335 10747 6341
rect 10796 6344 12532 6372
rect 10796 6313 10824 6344
rect 12526 6332 12532 6344
rect 12584 6332 12590 6384
rect 14292 6381 14320 6412
rect 14277 6375 14335 6381
rect 14277 6341 14289 6375
rect 14323 6372 14335 6375
rect 15286 6372 15292 6384
rect 14323 6344 15292 6372
rect 14323 6341 14335 6344
rect 14277 6335 14335 6341
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 10321 6307 10379 6313
rect 7432 6276 10272 6304
rect 7432 6264 7438 6276
rect 5960 6208 6776 6236
rect 5960 6196 5966 6208
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6880 6208 7205 6236
rect 6880 6196 6886 6208
rect 7193 6205 7205 6208
rect 7239 6236 7251 6239
rect 7745 6239 7803 6245
rect 7239 6208 7512 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 6181 6171 6239 6177
rect 4120 6140 6132 6168
rect 4120 6128 4126 6140
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 5353 6103 5411 6109
rect 5353 6100 5365 6103
rect 4580 6072 5365 6100
rect 4580 6060 4586 6072
rect 5353 6069 5365 6072
rect 5399 6069 5411 6103
rect 5353 6063 5411 6069
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 5902 6100 5908 6112
rect 5500 6072 5908 6100
rect 5500 6060 5506 6072
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 5994 6060 6000 6112
rect 6052 6060 6058 6112
rect 6104 6100 6132 6140
rect 6181 6137 6193 6171
rect 6227 6168 6239 6171
rect 7374 6168 7380 6180
rect 6227 6140 7380 6168
rect 6227 6137 6239 6140
rect 6181 6131 6239 6137
rect 7374 6128 7380 6140
rect 7432 6128 7438 6180
rect 7484 6168 7512 6208
rect 7745 6205 7757 6239
rect 7791 6236 7803 6239
rect 7834 6236 7840 6248
rect 7791 6208 7840 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 8202 6196 8208 6248
rect 8260 6236 8266 6248
rect 8386 6236 8392 6248
rect 8260 6208 8392 6236
rect 8260 6196 8266 6208
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 8478 6196 8484 6248
rect 8536 6196 8542 6248
rect 10244 6236 10272 6276
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 10870 6304 10876 6316
rect 10827 6276 10876 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6304 11851 6307
rect 11882 6304 11888 6316
rect 11839 6276 11888 6304
rect 11839 6273 11851 6276
rect 11793 6267 11851 6273
rect 11348 6236 11376 6267
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 12216 6276 12265 6304
rect 12216 6264 12222 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 13630 6264 13636 6316
rect 13688 6264 13694 6316
rect 10244 6208 11376 6236
rect 11609 6239 11667 6245
rect 11609 6205 11621 6239
rect 11655 6236 11667 6239
rect 11698 6236 11704 6248
rect 11655 6208 11704 6236
rect 11655 6205 11667 6208
rect 11609 6199 11667 6205
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6236 12587 6239
rect 12575 6208 13676 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 13648 6180 13676 6208
rect 10410 6168 10416 6180
rect 7484 6140 10416 6168
rect 10410 6128 10416 6140
rect 10468 6128 10474 6180
rect 10505 6171 10563 6177
rect 10505 6137 10517 6171
rect 10551 6168 10563 6171
rect 10551 6140 12112 6168
rect 10551 6137 10563 6140
rect 10505 6131 10563 6137
rect 6362 6100 6368 6112
rect 6104 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6546 6060 6552 6112
rect 6604 6060 6610 6112
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 7834 6100 7840 6112
rect 7248 6072 7840 6100
rect 7248 6060 7254 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 8018 6060 8024 6112
rect 8076 6060 8082 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 10284 6072 11161 6100
rect 10284 6060 10290 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 12084 6100 12112 6140
rect 13630 6128 13636 6180
rect 13688 6128 13694 6180
rect 14274 6100 14280 6112
rect 12084 6072 14280 6100
rect 11149 6063 11207 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 1104 6010 14812 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 14812 6010
rect 1104 5936 14812 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 3234 5896 3240 5908
rect 2823 5868 3240 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4062 5896 4068 5908
rect 4019 5868 4068 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4154 5856 4160 5908
rect 4212 5856 4218 5908
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 5074 5896 5080 5908
rect 4571 5868 5080 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5626 5856 5632 5908
rect 5684 5896 5690 5908
rect 6178 5896 6184 5908
rect 5684 5868 6184 5896
rect 5684 5856 5690 5868
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 7285 5899 7343 5905
rect 7285 5865 7297 5899
rect 7331 5896 7343 5899
rect 8294 5896 8300 5908
rect 7331 5868 8300 5896
rect 7331 5865 7343 5868
rect 7285 5859 7343 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 8846 5896 8852 5908
rect 8720 5868 8852 5896
rect 8720 5856 8726 5868
rect 8846 5856 8852 5868
rect 8904 5896 8910 5908
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 8904 5868 9229 5896
rect 8904 5856 8910 5868
rect 9217 5865 9229 5868
rect 9263 5896 9275 5899
rect 10318 5896 10324 5908
rect 9263 5868 10324 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 10870 5856 10876 5908
rect 10928 5856 10934 5908
rect 11698 5896 11704 5908
rect 11348 5868 11704 5896
rect 1857 5831 1915 5837
rect 1857 5797 1869 5831
rect 1903 5828 1915 5831
rect 3694 5828 3700 5840
rect 1903 5800 3700 5828
rect 1903 5797 1915 5800
rect 1857 5791 1915 5797
rect 3694 5788 3700 5800
rect 3752 5788 3758 5840
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 4341 5831 4399 5837
rect 4341 5828 4353 5831
rect 3844 5800 4353 5828
rect 3844 5788 3850 5800
rect 4341 5797 4353 5800
rect 4387 5797 4399 5831
rect 4341 5791 4399 5797
rect 4985 5831 5043 5837
rect 4985 5797 4997 5831
rect 5031 5828 5043 5831
rect 5031 5800 5212 5828
rect 5031 5797 5043 5800
rect 4985 5791 5043 5797
rect 3326 5720 3332 5772
rect 3384 5720 3390 5772
rect 4522 5720 4528 5772
rect 4580 5760 4586 5772
rect 4580 5732 4660 5760
rect 4580 5720 4586 5732
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1673 5695 1731 5701
rect 1673 5692 1685 5695
rect 1544 5664 1685 5692
rect 1544 5652 1550 5664
rect 1673 5661 1685 5664
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1688 5624 1716 5655
rect 2958 5652 2964 5704
rect 3016 5652 3022 5704
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5692 3111 5695
rect 3602 5692 3608 5704
rect 3099 5664 3608 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 4062 5692 4068 5704
rect 3712 5664 4068 5692
rect 2225 5627 2283 5633
rect 2225 5624 2237 5627
rect 1688 5596 2237 5624
rect 2225 5593 2237 5596
rect 2271 5624 2283 5627
rect 3712 5624 3740 5664
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4430 5652 4436 5704
rect 4488 5652 4494 5704
rect 4632 5701 4660 5732
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4893 5695 4951 5701
rect 4893 5694 4905 5695
rect 4816 5692 4905 5694
rect 4617 5655 4675 5661
rect 4724 5666 4905 5692
rect 4724 5664 4844 5666
rect 2271 5596 3740 5624
rect 3789 5627 3847 5633
rect 2271 5593 2283 5596
rect 2225 5587 2283 5593
rect 3789 5593 3801 5627
rect 3835 5624 3847 5627
rect 3878 5624 3884 5636
rect 3835 5596 3884 5624
rect 3835 5593 3847 5596
rect 3789 5587 3847 5593
rect 3878 5584 3884 5596
rect 3936 5584 3942 5636
rect 4522 5584 4528 5636
rect 4580 5624 4586 5636
rect 4724 5624 4752 5664
rect 4893 5661 4905 5666
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5184 5692 5212 5800
rect 6730 5788 6736 5840
rect 6788 5828 6794 5840
rect 7745 5831 7803 5837
rect 7745 5828 7757 5831
rect 6788 5800 7757 5828
rect 6788 5788 6794 5800
rect 7745 5797 7757 5800
rect 7791 5797 7803 5831
rect 7745 5791 7803 5797
rect 8389 5831 8447 5837
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 11146 5828 11152 5840
rect 8435 5800 11152 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 11146 5788 11152 5800
rect 11204 5788 11210 5840
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 5626 5760 5632 5772
rect 5307 5732 5632 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 5626 5720 5632 5732
rect 5684 5720 5690 5772
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 9950 5760 9956 5772
rect 5960 5732 9956 5760
rect 5960 5720 5966 5732
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 10410 5720 10416 5772
rect 10468 5760 10474 5772
rect 11348 5760 11376 5868
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 14277 5899 14335 5905
rect 14277 5896 14289 5899
rect 13412 5868 14289 5896
rect 13412 5856 13418 5868
rect 14277 5865 14289 5868
rect 14323 5865 14335 5899
rect 14277 5859 14335 5865
rect 11514 5788 11520 5840
rect 11572 5828 11578 5840
rect 11572 5800 12020 5828
rect 11572 5788 11578 5800
rect 10468 5732 11376 5760
rect 10468 5720 10474 5732
rect 11422 5720 11428 5772
rect 11480 5760 11486 5772
rect 11882 5760 11888 5772
rect 11480 5732 11888 5760
rect 11480 5720 11486 5732
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 11992 5760 12020 5800
rect 14090 5788 14096 5840
rect 14148 5788 14154 5840
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 11992 5732 12173 5760
rect 12161 5729 12173 5732
rect 12207 5729 12219 5763
rect 12161 5723 12219 5729
rect 13909 5763 13967 5769
rect 13909 5729 13921 5763
rect 13955 5760 13967 5763
rect 14182 5760 14188 5772
rect 13955 5732 14188 5760
rect 13955 5729 13967 5732
rect 13909 5723 13967 5729
rect 14182 5720 14188 5732
rect 14240 5760 14246 5772
rect 14918 5760 14924 5772
rect 14240 5732 14924 5760
rect 14240 5720 14246 5732
rect 14918 5720 14924 5732
rect 14976 5720 14982 5772
rect 5184 5664 5304 5692
rect 5077 5655 5135 5661
rect 4580 5596 4752 5624
rect 4801 5627 4859 5633
rect 4580 5584 4586 5596
rect 4801 5593 4813 5627
rect 4847 5624 4859 5627
rect 4982 5624 4988 5636
rect 4847 5596 4988 5624
rect 4847 5593 4859 5596
rect 4801 5587 4859 5593
rect 4982 5584 4988 5596
rect 5040 5584 5046 5636
rect 5092 5624 5120 5655
rect 5166 5624 5172 5636
rect 5092 5596 5172 5624
rect 5166 5584 5172 5596
rect 5224 5584 5230 5636
rect 5276 5624 5304 5664
rect 6638 5652 6644 5704
rect 6696 5652 6702 5704
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 7558 5692 7564 5704
rect 7423 5664 7564 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7834 5692 7840 5704
rect 7668 5664 7840 5692
rect 5442 5624 5448 5636
rect 5276 5596 5448 5624
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 5537 5627 5595 5633
rect 5537 5593 5549 5627
rect 5583 5593 5595 5627
rect 7668 5624 7696 5664
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8076 5664 8248 5692
rect 8076 5652 8082 5664
rect 5537 5587 5595 5593
rect 6840 5596 7696 5624
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 3602 5556 3608 5568
rect 3191 5528 3608 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 3999 5559 4057 5565
rect 3999 5525 4011 5559
rect 4045 5556 4057 5559
rect 4154 5556 4160 5568
rect 4045 5528 4160 5556
rect 4045 5525 4057 5528
rect 3999 5519 4057 5525
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 5552 5556 5580 5587
rect 6840 5556 6868 5596
rect 7742 5584 7748 5636
rect 7800 5584 7806 5636
rect 7852 5624 7880 5652
rect 8113 5627 8171 5633
rect 8113 5624 8125 5627
rect 7852 5596 8125 5624
rect 8113 5593 8125 5596
rect 8159 5593 8171 5627
rect 8220 5624 8248 5664
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8665 5695 8723 5701
rect 8665 5692 8677 5695
rect 8444 5664 8677 5692
rect 8444 5652 8450 5664
rect 8665 5661 8677 5664
rect 8711 5661 8723 5695
rect 8665 5655 8723 5661
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 9364 5664 11621 5692
rect 9364 5652 9370 5664
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 11790 5652 11796 5704
rect 11848 5652 11854 5704
rect 9122 5624 9128 5636
rect 8220 5596 9128 5624
rect 8113 5587 8171 5593
rect 9122 5584 9128 5596
rect 9180 5584 9186 5636
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 14245 5627 14303 5633
rect 14245 5624 14257 5627
rect 9732 5596 12650 5624
rect 14016 5596 14257 5624
rect 9732 5584 9738 5596
rect 4488 5528 6868 5556
rect 7009 5559 7067 5565
rect 4488 5516 4494 5528
rect 7009 5525 7021 5559
rect 7055 5556 7067 5559
rect 7374 5556 7380 5568
rect 7055 5528 7380 5556
rect 7055 5525 7067 5528
rect 7009 5519 7067 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 7760 5556 7788 5584
rect 7524 5528 7788 5556
rect 7929 5559 7987 5565
rect 7524 5516 7530 5528
rect 7929 5525 7941 5559
rect 7975 5556 7987 5559
rect 8478 5556 8484 5568
rect 7975 5528 8484 5556
rect 7975 5525 7987 5528
rect 7929 5519 7987 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 9364 5528 9505 5556
rect 9364 5516 9370 5528
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 9493 5519 9551 5525
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 10318 5556 10324 5568
rect 9824 5528 10324 5556
rect 9824 5516 9830 5528
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 11425 5559 11483 5565
rect 11425 5556 11437 5559
rect 10468 5528 11437 5556
rect 10468 5516 10474 5528
rect 11425 5525 11437 5528
rect 11471 5525 11483 5559
rect 11425 5519 11483 5525
rect 11606 5516 11612 5568
rect 11664 5516 11670 5568
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 14016 5556 14044 5596
rect 14245 5593 14257 5596
rect 14291 5593 14303 5627
rect 14245 5587 14303 5593
rect 14461 5627 14519 5633
rect 14461 5593 14473 5627
rect 14507 5593 14519 5627
rect 14461 5587 14519 5593
rect 11756 5528 14044 5556
rect 11756 5516 11762 5528
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 14476 5556 14504 5587
rect 14148 5528 14504 5556
rect 14148 5516 14154 5528
rect 1104 5466 14812 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 14812 5466
rect 1104 5392 14812 5414
rect 3234 5312 3240 5364
rect 3292 5312 3298 5364
rect 3602 5312 3608 5364
rect 3660 5312 3666 5364
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4341 5355 4399 5361
rect 4341 5352 4353 5355
rect 4212 5324 4353 5352
rect 4212 5312 4218 5324
rect 4341 5321 4353 5324
rect 4387 5352 4399 5355
rect 4614 5352 4620 5364
rect 4387 5324 4620 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4982 5312 4988 5364
rect 5040 5352 5046 5364
rect 5040 5324 5304 5352
rect 5040 5312 5046 5324
rect 3418 5244 3424 5296
rect 3476 5284 3482 5296
rect 5077 5287 5135 5293
rect 5077 5284 5089 5287
rect 3476 5256 5089 5284
rect 3476 5244 3482 5256
rect 5077 5253 5089 5256
rect 5123 5284 5135 5287
rect 5166 5284 5172 5296
rect 5123 5256 5172 5284
rect 5123 5253 5135 5256
rect 5077 5247 5135 5253
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 5276 5293 5304 5324
rect 5350 5312 5356 5364
rect 5408 5352 5414 5364
rect 5461 5355 5519 5361
rect 5461 5352 5473 5355
rect 5408 5324 5473 5352
rect 5408 5312 5414 5324
rect 5461 5321 5473 5324
rect 5507 5321 5519 5355
rect 5461 5315 5519 5321
rect 6178 5312 6184 5364
rect 6236 5352 6242 5364
rect 9858 5352 9864 5364
rect 6236 5324 8800 5352
rect 6236 5312 6242 5324
rect 5261 5287 5319 5293
rect 5261 5253 5273 5287
rect 5307 5253 5319 5287
rect 5261 5247 5319 5253
rect 5718 5244 5724 5296
rect 5776 5284 5782 5296
rect 5813 5287 5871 5293
rect 5813 5284 5825 5287
rect 5776 5256 5825 5284
rect 5776 5244 5782 5256
rect 5813 5253 5825 5256
rect 5859 5253 5871 5287
rect 5813 5247 5871 5253
rect 6029 5287 6087 5293
rect 6029 5253 6041 5287
rect 6075 5284 6087 5287
rect 6454 5284 6460 5296
rect 6075 5256 6460 5284
rect 6075 5253 6087 5256
rect 6029 5247 6087 5253
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 6733 5287 6791 5293
rect 6733 5253 6745 5287
rect 6779 5284 6791 5287
rect 7190 5284 7196 5296
rect 6779 5256 7196 5284
rect 6779 5253 6791 5256
rect 6733 5247 6791 5253
rect 7190 5244 7196 5256
rect 7248 5244 7254 5296
rect 8018 5244 8024 5296
rect 8076 5244 8082 5296
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 4246 5216 4252 5228
rect 3384 5188 4252 5216
rect 3384 5176 3390 5188
rect 4246 5176 4252 5188
rect 4304 5216 4310 5228
rect 5736 5216 5764 5244
rect 8772 5225 8800 5324
rect 9600 5324 9864 5352
rect 4304 5188 5764 5216
rect 6549 5219 6607 5225
rect 4304 5176 4310 5188
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 8757 5219 8815 5225
rect 6595 5188 7328 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 4522 5108 4528 5160
rect 4580 5148 4586 5160
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 4580 5120 4813 5148
rect 4580 5108 4586 5120
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 6365 5151 6423 5157
rect 4801 5111 4859 5117
rect 5552 5120 6316 5148
rect 4338 5040 4344 5092
rect 4396 5080 4402 5092
rect 5552 5080 5580 5120
rect 4396 5052 5580 5080
rect 5629 5083 5687 5089
rect 4396 5040 4402 5052
rect 5629 5049 5641 5083
rect 5675 5080 5687 5083
rect 5810 5080 5816 5092
rect 5675 5052 5816 5080
rect 5675 5049 5687 5052
rect 5629 5043 5687 5049
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 6178 5040 6184 5092
rect 6236 5040 6242 5092
rect 6288 5080 6316 5120
rect 6365 5117 6377 5151
rect 6411 5148 6423 5151
rect 6730 5148 6736 5160
rect 6411 5120 6736 5148
rect 6411 5117 6423 5120
rect 6365 5111 6423 5117
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 7300 5148 7328 5188
rect 8757 5185 8769 5219
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 9306 5176 9312 5228
rect 9364 5176 9370 5228
rect 9490 5176 9496 5228
rect 9548 5176 9554 5228
rect 9600 5225 9628 5324
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 14182 5352 14188 5364
rect 12492 5324 14188 5352
rect 12492 5312 12498 5324
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 11790 5244 11796 5296
rect 11848 5244 11854 5296
rect 11974 5244 11980 5296
rect 12032 5244 12038 5296
rect 12713 5287 12771 5293
rect 12713 5253 12725 5287
rect 12759 5284 12771 5287
rect 12986 5284 12992 5296
rect 12759 5256 12992 5284
rect 12759 5253 12771 5256
rect 12713 5247 12771 5253
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 14274 5244 14280 5296
rect 14332 5284 14338 5296
rect 14461 5287 14519 5293
rect 14461 5284 14473 5287
rect 14332 5256 14473 5284
rect 14332 5244 14338 5256
rect 14461 5253 14473 5256
rect 14507 5253 14519 5287
rect 14461 5247 14519 5253
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 11808 5216 11836 5244
rect 9585 5179 9643 5185
rect 8386 5148 8392 5160
rect 7300 5120 8392 5148
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8481 5151 8539 5157
rect 8481 5117 8493 5151
rect 8527 5148 8539 5151
rect 8527 5120 9352 5148
rect 8527 5117 8539 5120
rect 8481 5111 8539 5117
rect 7009 5083 7067 5089
rect 7009 5080 7021 5083
rect 6288 5052 7021 5080
rect 7009 5049 7021 5052
rect 7055 5049 7067 5083
rect 7009 5043 7067 5049
rect 8846 5040 8852 5092
rect 8904 5080 8910 5092
rect 9324 5080 9352 5120
rect 9858 5108 9864 5160
rect 9916 5108 9922 5160
rect 10980 5080 11008 5202
rect 11072 5188 11836 5216
rect 11072 5160 11100 5188
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 11940 5188 12449 5216
rect 11940 5176 11946 5188
rect 12437 5185 12449 5188
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 13814 5176 13820 5228
rect 13872 5176 13878 5228
rect 11054 5108 11060 5160
rect 11112 5108 11118 5160
rect 11330 5108 11336 5160
rect 11388 5108 11394 5160
rect 13078 5148 13084 5160
rect 12544 5120 13084 5148
rect 12544 5080 12572 5120
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 8904 5052 9260 5080
rect 9324 5052 9720 5080
rect 10980 5052 12572 5080
rect 8904 5040 8910 5052
rect 5445 5015 5503 5021
rect 5445 4981 5457 5015
rect 5491 5012 5503 5015
rect 5902 5012 5908 5024
rect 5491 4984 5908 5012
rect 5491 4981 5503 4984
rect 5445 4975 5503 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 5994 4972 6000 5024
rect 6052 4972 6058 5024
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 6822 5012 6828 5024
rect 6420 4984 6828 5012
rect 6420 4972 6426 4984
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 9125 5015 9183 5021
rect 9125 5012 9137 5015
rect 7432 4984 9137 5012
rect 7432 4972 7438 4984
rect 9125 4981 9137 4984
rect 9171 4981 9183 5015
rect 9232 5012 9260 5052
rect 9309 5015 9367 5021
rect 9309 5012 9321 5015
rect 9232 4984 9321 5012
rect 9125 4975 9183 4981
rect 9309 4981 9321 4984
rect 9355 5012 9367 5015
rect 9398 5012 9404 5024
rect 9355 4984 9404 5012
rect 9355 4981 9367 4984
rect 9309 4975 9367 4981
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 9692 5012 9720 5052
rect 10226 5012 10232 5024
rect 9692 4984 10232 5012
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 11609 5015 11667 5021
rect 11609 5012 11621 5015
rect 10928 4984 11621 5012
rect 10928 4972 10934 4984
rect 11609 4981 11621 4984
rect 11655 4981 11667 5015
rect 11609 4975 11667 4981
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 11848 4984 12265 5012
rect 11848 4972 11854 4984
rect 12253 4981 12265 4984
rect 12299 5012 12311 5015
rect 13262 5012 13268 5024
rect 12299 4984 13268 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 1104 4922 14812 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 14812 4922
rect 1104 4848 14812 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 1949 4811 2007 4817
rect 1949 4808 1961 4811
rect 1360 4780 1961 4808
rect 1360 4768 1366 4780
rect 1949 4777 1961 4780
rect 1995 4777 2007 4811
rect 3513 4811 3571 4817
rect 3513 4808 3525 4811
rect 1949 4771 2007 4777
rect 2240 4780 3525 4808
rect 1026 4700 1032 4752
rect 1084 4740 1090 4752
rect 2240 4740 2268 4780
rect 3513 4777 3525 4780
rect 3559 4777 3571 4811
rect 3513 4771 3571 4777
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 7374 4808 7380 4820
rect 5684 4780 7380 4808
rect 5684 4768 5690 4780
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7837 4811 7895 4817
rect 7837 4777 7849 4811
rect 7883 4808 7895 4811
rect 7926 4808 7932 4820
rect 7883 4780 7932 4808
rect 7883 4777 7895 4780
rect 7837 4771 7895 4777
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8021 4811 8079 4817
rect 8021 4777 8033 4811
rect 8067 4777 8079 4811
rect 8021 4771 8079 4777
rect 8389 4811 8447 4817
rect 8389 4777 8401 4811
rect 8435 4808 8447 4811
rect 9674 4808 9680 4820
rect 8435 4780 9680 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 1084 4712 2268 4740
rect 2317 4743 2375 4749
rect 1084 4700 1090 4712
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 2498 4740 2504 4752
rect 2363 4712 2504 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 2498 4700 2504 4712
rect 2556 4700 2562 4752
rect 2869 4743 2927 4749
rect 2869 4709 2881 4743
rect 2915 4740 2927 4743
rect 3234 4740 3240 4752
rect 2915 4712 3240 4740
rect 2915 4709 2927 4712
rect 2869 4703 2927 4709
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 5350 4700 5356 4752
rect 5408 4700 5414 4752
rect 8036 4740 8064 4771
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9824 4780 9965 4808
rect 9824 4768 9830 4780
rect 9953 4777 9965 4780
rect 9999 4808 10011 4811
rect 10778 4808 10784 4820
rect 9999 4780 10784 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11149 4811 11207 4817
rect 11149 4777 11161 4811
rect 11195 4808 11207 4811
rect 13354 4808 13360 4820
rect 11195 4780 13360 4808
rect 11195 4777 11207 4780
rect 11149 4771 11207 4777
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 14090 4808 14096 4820
rect 13679 4780 14096 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 14458 4768 14464 4820
rect 14516 4768 14522 4820
rect 8662 4740 8668 4752
rect 5460 4712 5948 4740
rect 8036 4712 8668 4740
rect 2406 4672 2412 4684
rect 2148 4644 2412 4672
rect 1762 4564 1768 4616
rect 1820 4564 1826 4616
rect 1854 4564 1860 4616
rect 1912 4604 1918 4616
rect 2148 4613 2176 4644
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 5460 4672 5488 4712
rect 2700 4644 5488 4672
rect 2700 4613 2728 4644
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 5920 4672 5948 4712
rect 8662 4700 8668 4712
rect 8720 4700 8726 4752
rect 8941 4743 8999 4749
rect 8941 4709 8953 4743
rect 8987 4740 8999 4743
rect 13998 4740 14004 4752
rect 8987 4712 14004 4740
rect 8987 4709 8999 4712
rect 8941 4703 8999 4709
rect 13998 4700 14004 4712
rect 14056 4700 14062 4752
rect 6730 4672 6736 4684
rect 5592 4644 5856 4672
rect 5920 4644 6736 4672
rect 5592 4632 5598 4644
rect 5828 4616 5856 4644
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7561 4675 7619 4681
rect 7561 4672 7573 4675
rect 6880 4644 7573 4672
rect 6880 4632 6886 4644
rect 7561 4641 7573 4644
rect 7607 4672 7619 4675
rect 8846 4672 8852 4684
rect 7607 4644 8852 4672
rect 7607 4641 7619 4644
rect 7561 4635 7619 4641
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 9766 4672 9772 4684
rect 9324 4644 9772 4672
rect 1949 4607 2007 4613
rect 1949 4604 1961 4607
rect 1912 4576 1961 4604
rect 1912 4564 1918 4576
rect 1949 4573 1961 4576
rect 1995 4573 2007 4607
rect 1949 4567 2007 4573
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4573 2743 4607
rect 2685 4567 2743 4573
rect 842 4496 848 4548
rect 900 4536 906 4548
rect 2332 4536 2360 4567
rect 3234 4564 3240 4616
rect 3292 4564 3298 4616
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 5169 4607 5227 4613
rect 3651 4576 4108 4604
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 2958 4536 2964 4548
rect 900 4508 2964 4536
rect 900 4496 906 4508
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 1673 4471 1731 4477
rect 1673 4437 1685 4471
rect 1719 4468 1731 4471
rect 1762 4468 1768 4480
rect 1719 4440 1768 4468
rect 1719 4437 1731 4440
rect 1673 4431 1731 4437
rect 1762 4428 1768 4440
rect 1820 4468 1826 4480
rect 2498 4468 2504 4480
rect 1820 4440 2504 4468
rect 1820 4428 1826 4440
rect 2498 4428 2504 4440
rect 2556 4428 2562 4480
rect 3053 4471 3111 4477
rect 3053 4437 3065 4471
rect 3099 4468 3111 4471
rect 3326 4468 3332 4480
rect 3099 4440 3332 4468
rect 3099 4437 3111 4440
rect 3053 4431 3111 4437
rect 3326 4428 3332 4440
rect 3384 4428 3390 4480
rect 4080 4477 4108 4576
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5626 4604 5632 4616
rect 5215 4576 5632 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 5810 4564 5816 4616
rect 5868 4564 5874 4616
rect 8297 4607 8355 4613
rect 8297 4573 8309 4607
rect 8343 4604 8355 4607
rect 8386 4604 8392 4616
rect 8343 4576 8392 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 9324 4613 9352 4644
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 11054 4672 11060 4684
rect 10152 4644 11060 4672
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 6089 4539 6147 4545
rect 6089 4536 6101 4539
rect 5500 4508 6101 4536
rect 5500 4496 5506 4508
rect 6089 4505 6101 4508
rect 6135 4505 6147 4539
rect 6089 4499 6147 4505
rect 6546 4496 6552 4548
rect 6604 4496 6610 4548
rect 8205 4539 8263 4545
rect 8205 4505 8217 4539
rect 8251 4536 8263 4539
rect 8938 4536 8944 4548
rect 8251 4508 8944 4536
rect 8251 4505 8263 4508
rect 8205 4499 8263 4505
rect 8938 4496 8944 4508
rect 8996 4496 9002 4548
rect 9416 4536 9444 4567
rect 9582 4564 9588 4616
rect 9640 4564 9646 4616
rect 9766 4536 9772 4548
rect 9416 4508 9772 4536
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 4065 4471 4123 4477
rect 4065 4437 4077 4471
rect 4111 4468 4123 4471
rect 4154 4468 4160 4480
rect 4111 4440 4160 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 4982 4428 4988 4480
rect 5040 4468 5046 4480
rect 5721 4471 5779 4477
rect 5721 4468 5733 4471
rect 5040 4440 5733 4468
rect 5040 4428 5046 4440
rect 5721 4437 5733 4440
rect 5767 4468 5779 4471
rect 5994 4468 6000 4480
rect 5767 4440 6000 4468
rect 5767 4437 5779 4440
rect 5721 4431 5779 4437
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 8005 4471 8063 4477
rect 8005 4437 8017 4471
rect 8051 4468 8063 4471
rect 8478 4468 8484 4480
rect 8051 4440 8484 4468
rect 8051 4437 8063 4440
rect 8005 4431 8063 4437
rect 8478 4428 8484 4440
rect 8536 4428 8542 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 10152 4468 10180 4644
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 12158 4672 12164 4684
rect 11296 4644 11744 4672
rect 11296 4632 11302 4644
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 10744 4576 11008 4604
rect 10744 4564 10750 4576
rect 10781 4539 10839 4545
rect 10781 4505 10793 4539
rect 10827 4536 10839 4539
rect 10870 4536 10876 4548
rect 10827 4508 10876 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 8720 4440 10180 4468
rect 8720 4428 8726 4440
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10597 4471 10655 4477
rect 10597 4468 10609 4471
rect 10284 4440 10609 4468
rect 10284 4428 10290 4440
rect 10597 4437 10609 4440
rect 10643 4468 10655 4471
rect 10796 4468 10824 4499
rect 10870 4496 10876 4508
rect 10928 4496 10934 4548
rect 10980 4545 11008 4576
rect 11514 4564 11520 4616
rect 11572 4613 11578 4616
rect 11716 4613 11744 4644
rect 11808 4644 12164 4672
rect 11808 4613 11836 4644
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12345 4675 12403 4681
rect 12345 4641 12357 4675
rect 12391 4672 12403 4675
rect 13446 4672 13452 4684
rect 12391 4644 13452 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 11572 4607 11621 4613
rect 11572 4573 11575 4607
rect 11609 4573 11621 4607
rect 11572 4567 11621 4573
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 11572 4564 11578 4567
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 11977 4607 12035 4613
rect 11977 4604 11989 4607
rect 11940 4576 11989 4604
rect 11940 4564 11946 4576
rect 11977 4573 11989 4576
rect 12023 4604 12035 4607
rect 12250 4604 12256 4616
rect 12023 4576 12256 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 12250 4564 12256 4576
rect 12308 4564 12314 4616
rect 10965 4539 11023 4545
rect 10965 4505 10977 4539
rect 11011 4505 11023 4539
rect 10965 4499 11023 4505
rect 10643 4440 10824 4468
rect 10980 4468 11008 4499
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 11333 4539 11391 4545
rect 11333 4536 11345 4539
rect 11112 4508 11345 4536
rect 11112 4496 11118 4508
rect 11333 4505 11345 4508
rect 11379 4505 11391 4539
rect 11333 4499 11391 4505
rect 12360 4468 12388 4635
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 12529 4607 12587 4613
rect 12529 4601 12541 4607
rect 10980 4440 12388 4468
rect 12452 4573 12541 4601
rect 12575 4573 12587 4607
rect 12452 4468 12480 4573
rect 12529 4567 12587 4573
rect 12621 4607 12679 4613
rect 12621 4573 12633 4607
rect 12667 4573 12679 4607
rect 12621 4567 12679 4573
rect 12636 4536 12664 4567
rect 12894 4564 12900 4616
rect 12952 4604 12958 4616
rect 13725 4607 13783 4613
rect 13725 4604 13737 4607
rect 12952 4576 13737 4604
rect 12952 4564 12958 4576
rect 13725 4573 13737 4576
rect 13771 4573 13783 4607
rect 13725 4567 13783 4573
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14826 4604 14832 4616
rect 14323 4576 14832 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14826 4564 14832 4576
rect 14884 4564 14890 4616
rect 13262 4536 13268 4548
rect 12636 4508 13268 4536
rect 13262 4496 13268 4508
rect 13320 4496 13326 4548
rect 13081 4471 13139 4477
rect 13081 4468 13093 4471
rect 12452 4440 13093 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 13081 4437 13093 4440
rect 13127 4468 13139 4471
rect 13170 4468 13176 4480
rect 13127 4440 13176 4468
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 13906 4428 13912 4480
rect 13964 4428 13970 4480
rect 1104 4378 14812 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 14812 4378
rect 1104 4304 14812 4326
rect 2958 4224 2964 4276
rect 3016 4224 3022 4276
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 3421 4267 3479 4273
rect 3421 4264 3433 4267
rect 3292 4236 3433 4264
rect 3292 4224 3298 4236
rect 3421 4233 3433 4236
rect 3467 4264 3479 4267
rect 4982 4264 4988 4276
rect 3467 4236 4988 4264
rect 3467 4233 3479 4236
rect 3421 4227 3479 4233
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 10686 4264 10692 4276
rect 5224 4236 10692 4264
rect 5224 4224 5230 4236
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 11606 4224 11612 4276
rect 11664 4264 11670 4276
rect 11790 4264 11796 4276
rect 11664 4236 11796 4264
rect 11664 4224 11670 4236
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 12434 4264 12440 4276
rect 12176 4236 12440 4264
rect 2590 4156 2596 4208
rect 2648 4196 2654 4208
rect 8389 4199 8447 4205
rect 8389 4196 8401 4199
rect 2648 4168 8401 4196
rect 2648 4156 2654 4168
rect 8389 4165 8401 4168
rect 8435 4196 8447 4199
rect 8478 4196 8484 4208
rect 8435 4168 8484 4196
rect 8435 4165 8447 4168
rect 8389 4159 8447 4165
rect 8478 4156 8484 4168
rect 8536 4196 8542 4208
rect 12176 4196 12204 4236
rect 12434 4224 12440 4236
rect 12492 4224 12498 4276
rect 13906 4224 13912 4276
rect 13964 4224 13970 4276
rect 8536 4168 12204 4196
rect 8536 4156 8542 4168
rect 12250 4156 12256 4208
rect 12308 4196 12314 4208
rect 12805 4199 12863 4205
rect 12805 4196 12817 4199
rect 12308 4168 12817 4196
rect 12308 4156 12314 4168
rect 12805 4165 12817 4168
rect 12851 4196 12863 4199
rect 14182 4196 14188 4208
rect 12851 4168 14188 4196
rect 12851 4165 12863 4168
rect 12805 4159 12863 4165
rect 14182 4156 14188 4168
rect 14240 4156 14246 4208
rect 14642 4196 14648 4208
rect 14292 4168 14648 4196
rect 2501 4131 2559 4137
rect 2501 4097 2513 4131
rect 2547 4128 2559 4131
rect 6822 4128 6828 4140
rect 2547 4100 6828 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 9306 4128 9312 4140
rect 6963 4100 9312 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 3050 4020 3056 4072
rect 3108 4060 3114 4072
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 3108 4032 6101 4060
rect 3108 4020 3114 4032
rect 6089 4029 6101 4032
rect 6135 4060 6147 4063
rect 6932 4060 6960 4091
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9640 4100 11284 4128
rect 9640 4088 9646 4100
rect 6135 4032 6960 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 7006 4020 7012 4072
rect 7064 4020 7070 4072
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8444 4032 9137 4060
rect 8444 4020 8450 4032
rect 9125 4029 9137 4032
rect 9171 4060 9183 4063
rect 10870 4060 10876 4072
rect 9171 4032 10876 4060
rect 9171 4029 9183 4032
rect 9125 4023 9183 4029
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 1578 3952 1584 4004
rect 1636 3992 1642 4004
rect 2685 3995 2743 4001
rect 2685 3992 2697 3995
rect 1636 3964 2697 3992
rect 1636 3952 1642 3964
rect 2685 3961 2697 3964
rect 2731 3961 2743 3995
rect 2685 3955 2743 3961
rect 5718 3952 5724 4004
rect 5776 3952 5782 4004
rect 6546 3952 6552 4004
rect 6604 3952 6610 4004
rect 7745 3995 7803 4001
rect 7745 3961 7757 3995
rect 7791 3992 7803 3995
rect 9398 3992 9404 4004
rect 7791 3964 9404 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 9582 3952 9588 4004
rect 9640 3952 9646 4004
rect 11256 4001 11284 4100
rect 11422 4088 11428 4140
rect 11480 4128 11486 4140
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 11480 4100 11805 4128
rect 11480 4088 11486 4100
rect 11793 4097 11805 4100
rect 11839 4128 11851 4131
rect 11977 4131 12035 4137
rect 11977 4128 11989 4131
rect 11839 4100 11989 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 11977 4097 11989 4100
rect 12023 4097 12035 4131
rect 11977 4091 12035 4097
rect 13354 4088 13360 4140
rect 13412 4128 13418 4140
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13412 4100 13737 4128
rect 13412 4088 13418 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11532 4032 12173 4060
rect 11241 3995 11299 4001
rect 11241 3961 11253 3995
rect 11287 3992 11299 3995
rect 11422 3992 11428 4004
rect 11287 3964 11428 3992
rect 11287 3961 11299 3964
rect 11241 3955 11299 3961
rect 11422 3952 11428 3964
rect 11480 3952 11486 4004
rect 5736 3924 5764 3952
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 5736 3896 8769 3924
rect 8757 3893 8769 3896
rect 8803 3924 8815 3927
rect 9600 3924 9628 3952
rect 8803 3896 9628 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 11532 3924 11560 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 12176 3992 12204 4023
rect 13170 4020 13176 4072
rect 13228 4060 13234 4072
rect 14016 4060 14044 4091
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 14292 4137 14320 4168
rect 14642 4156 14648 4168
rect 14700 4156 14706 4208
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 14148 4100 14289 4128
rect 14148 4088 14154 4100
rect 14277 4097 14289 4100
rect 14323 4097 14335 4131
rect 14277 4091 14335 4097
rect 14366 4088 14372 4140
rect 14424 4088 14430 4140
rect 13228 4032 14044 4060
rect 13228 4020 13234 4032
rect 13188 3992 13216 4020
rect 12176 3964 13216 3992
rect 13446 3952 13452 4004
rect 13504 3952 13510 4004
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14093 3995 14151 4001
rect 14093 3992 14105 3995
rect 13872 3964 14105 3992
rect 13872 3952 13878 3964
rect 14093 3961 14105 3964
rect 14139 3961 14151 3995
rect 14093 3955 14151 3961
rect 9732 3896 11560 3924
rect 9732 3884 9738 3896
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 13170 3924 13176 3936
rect 12584 3896 13176 3924
rect 12584 3884 12590 3896
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 1104 3834 14812 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 14812 3834
rect 1104 3760 14812 3782
rect 1394 3680 1400 3732
rect 1452 3720 1458 3732
rect 1489 3723 1547 3729
rect 1489 3720 1501 3723
rect 1452 3692 1501 3720
rect 1452 3680 1458 3692
rect 1489 3689 1501 3692
rect 1535 3689 1547 3723
rect 1489 3683 1547 3689
rect 2501 3723 2559 3729
rect 2501 3689 2513 3723
rect 2547 3720 2559 3723
rect 2590 3720 2596 3732
rect 2547 3692 2596 3720
rect 2547 3689 2559 3692
rect 2501 3683 2559 3689
rect 2516 3584 2544 3683
rect 2590 3680 2596 3692
rect 2648 3680 2654 3732
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 4856 3692 6837 3720
rect 4856 3680 4862 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 8938 3720 8944 3732
rect 7708 3692 8944 3720
rect 7708 3680 7714 3692
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9858 3720 9864 3732
rect 9539 3692 9864 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9858 3680 9864 3692
rect 9916 3720 9922 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 9916 3692 10057 3720
rect 9916 3680 9922 3692
rect 10045 3689 10057 3692
rect 10091 3720 10103 3723
rect 10318 3720 10324 3732
rect 10091 3692 10324 3720
rect 10091 3689 10103 3692
rect 10045 3683 10103 3689
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 11701 3723 11759 3729
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 13725 3723 13783 3729
rect 11747 3692 13676 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 4614 3612 4620 3664
rect 4672 3652 4678 3664
rect 4672 3624 7328 3652
rect 4672 3612 4678 3624
rect 1504 3556 2544 3584
rect 1504 3525 1532 3556
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 7300 3584 7328 3624
rect 7374 3612 7380 3664
rect 7432 3652 7438 3664
rect 8573 3655 8631 3661
rect 8573 3652 8585 3655
rect 7432 3624 8585 3652
rect 7432 3612 7438 3624
rect 8573 3621 8585 3624
rect 8619 3621 8631 3655
rect 8573 3615 8631 3621
rect 9677 3655 9735 3661
rect 9677 3621 9689 3655
rect 9723 3652 9735 3655
rect 12986 3652 12992 3664
rect 9723 3624 12992 3652
rect 9723 3621 9735 3624
rect 9677 3615 9735 3621
rect 12986 3612 12992 3624
rect 13044 3612 13050 3664
rect 9122 3584 9128 3596
rect 5316 3556 7144 3584
rect 7300 3556 9128 3584
rect 5316 3544 5322 3556
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3516 1823 3519
rect 1854 3516 1860 3528
rect 1811 3488 1860 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 4430 3476 4436 3528
rect 4488 3516 4494 3528
rect 7116 3525 7144 3556
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 4488 3488 6929 3516
rect 4488 3476 4494 3488
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3516 7343 3519
rect 7466 3516 7472 3528
rect 7331 3488 7472 3516
rect 7331 3485 7343 3488
rect 7285 3479 7343 3485
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 6733 3451 6791 3457
rect 6733 3448 6745 3451
rect 6696 3420 6745 3448
rect 6696 3408 6702 3420
rect 6733 3417 6745 3420
rect 6779 3448 6791 3451
rect 7024 3448 7052 3479
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 7616 3488 8033 3516
rect 7616 3476 7622 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 7374 3448 7380 3460
rect 6779 3420 7380 3448
rect 6779 3417 6791 3420
rect 6733 3411 6791 3417
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 8036 3448 8064 3479
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8312 3525 8340 3556
rect 9122 3544 9128 3556
rect 9180 3544 9186 3596
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 12434 3584 12440 3596
rect 9272 3556 12440 3584
rect 9272 3544 9278 3556
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 13446 3584 13452 3596
rect 12544 3556 13452 3584
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 8168 3488 8217 3516
rect 8168 3476 8174 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8570 3516 8576 3528
rect 8435 3488 8576 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 10134 3516 10140 3528
rect 9324 3488 10140 3516
rect 8662 3448 8668 3460
rect 8036 3420 8668 3448
rect 8662 3408 8668 3420
rect 8720 3408 8726 3460
rect 9324 3457 9352 3488
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 12544 3516 12572 3556
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 13648 3584 13676 3692
rect 13725 3689 13737 3723
rect 13771 3720 13783 3723
rect 14274 3720 14280 3732
rect 13771 3692 14280 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 14090 3612 14096 3664
rect 14148 3612 14154 3664
rect 15654 3584 15660 3596
rect 13648 3556 15660 3584
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 12986 3516 12992 3528
rect 10928 3488 12572 3516
rect 12636 3488 12992 3516
rect 10928 3476 10934 3488
rect 9309 3451 9367 3457
rect 9309 3417 9321 3451
rect 9355 3417 9367 3451
rect 9309 3411 9367 3417
rect 9525 3451 9583 3457
rect 9525 3417 9537 3451
rect 9571 3448 9583 3451
rect 11054 3448 11060 3460
rect 9571 3420 11060 3448
rect 9571 3417 9583 3420
rect 9525 3411 9583 3417
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 11790 3448 11796 3460
rect 11480 3420 11796 3448
rect 11480 3408 11486 3420
rect 11790 3408 11796 3420
rect 11848 3448 11854 3460
rect 11885 3451 11943 3457
rect 11885 3448 11897 3451
rect 11848 3420 11897 3448
rect 11848 3408 11854 3420
rect 11885 3417 11897 3420
rect 11931 3417 11943 3451
rect 11885 3411 11943 3417
rect 1673 3383 1731 3389
rect 1673 3349 1685 3383
rect 1719 3380 1731 3383
rect 2133 3383 2191 3389
rect 2133 3380 2145 3383
rect 1719 3352 2145 3380
rect 1719 3349 1731 3352
rect 1673 3343 1731 3349
rect 2133 3349 2145 3352
rect 2179 3380 2191 3383
rect 7650 3380 7656 3392
rect 2179 3352 7656 3380
rect 2179 3349 2191 3352
rect 2133 3343 2191 3349
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 9214 3380 9220 3392
rect 8812 3352 9220 3380
rect 8812 3340 8818 3352
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 10134 3340 10140 3392
rect 10192 3380 10198 3392
rect 11238 3380 11244 3392
rect 10192 3352 11244 3380
rect 10192 3340 10198 3352
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11514 3340 11520 3392
rect 11572 3340 11578 3392
rect 11685 3383 11743 3389
rect 11685 3349 11697 3383
rect 11731 3380 11743 3383
rect 12342 3380 12348 3392
rect 11731 3352 12348 3380
rect 11731 3349 11743 3352
rect 11685 3343 11743 3349
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 12636 3380 12664 3488
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13078 3476 13084 3528
rect 13136 3476 13142 3528
rect 14182 3476 14188 3528
rect 14240 3476 14246 3528
rect 14200 3448 14228 3476
rect 14461 3451 14519 3457
rect 14461 3448 14473 3451
rect 14200 3420 14473 3448
rect 14461 3417 14473 3420
rect 14507 3417 14519 3451
rect 14461 3411 14519 3417
rect 12483 3352 12664 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 12710 3340 12716 3392
rect 12768 3380 12774 3392
rect 12805 3383 12863 3389
rect 12805 3380 12817 3383
rect 12768 3352 12817 3380
rect 12768 3340 12774 3352
rect 12805 3349 12817 3352
rect 12851 3349 12863 3383
rect 12805 3343 12863 3349
rect 14261 3383 14319 3389
rect 14261 3349 14273 3383
rect 14307 3380 14319 3383
rect 14734 3380 14740 3392
rect 14307 3352 14740 3380
rect 14307 3349 14319 3352
rect 14261 3343 14319 3349
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 1104 3290 14812 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 14812 3290
rect 1104 3216 14812 3238
rect 3142 3136 3148 3188
rect 3200 3136 3206 3188
rect 3786 3176 3792 3188
rect 3252 3148 3792 3176
rect 3252 3108 3280 3148
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8570 3176 8576 3188
rect 7883 3148 8576 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8846 3136 8852 3188
rect 8904 3136 8910 3188
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 9180 3148 9505 3176
rect 9180 3136 9186 3148
rect 9493 3145 9505 3148
rect 9539 3145 9551 3179
rect 9493 3139 9551 3145
rect 9858 3136 9864 3188
rect 9916 3136 9922 3188
rect 10597 3179 10655 3185
rect 10597 3145 10609 3179
rect 10643 3176 10655 3179
rect 10962 3176 10968 3188
rect 10643 3148 10968 3176
rect 10643 3145 10655 3148
rect 10597 3139 10655 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11790 3176 11796 3188
rect 11072 3148 11796 3176
rect 3160 3080 3280 3108
rect 3421 3111 3479 3117
rect 3160 3049 3188 3080
rect 3421 3077 3433 3111
rect 3467 3108 3479 3111
rect 4430 3108 4436 3120
rect 3467 3080 4436 3108
rect 3467 3077 3479 3080
rect 3421 3071 3479 3077
rect 4430 3068 4436 3080
rect 4488 3068 4494 3120
rect 8665 3111 8723 3117
rect 8665 3077 8677 3111
rect 8711 3108 8723 3111
rect 8754 3108 8760 3120
rect 8711 3080 8760 3108
rect 8711 3077 8723 3080
rect 8665 3071 8723 3077
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 9140 3108 9168 3136
rect 8956 3080 9168 3108
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 3510 3040 3516 3052
rect 3283 3012 3516 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 5994 3000 6000 3052
rect 6052 3040 6058 3052
rect 8956 3049 8984 3080
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 11072 3108 11100 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 12434 3176 12440 3188
rect 11931 3148 12440 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12434 3136 12440 3148
rect 12492 3176 12498 3188
rect 12492 3148 14412 3176
rect 12492 3136 12498 3148
rect 9272 3080 11100 3108
rect 9272 3068 9278 3080
rect 11146 3068 11152 3120
rect 11204 3108 11210 3120
rect 12253 3111 12311 3117
rect 12253 3108 12265 3111
rect 11204 3080 12265 3108
rect 11204 3068 11210 3080
rect 12253 3077 12265 3080
rect 12299 3077 12311 3111
rect 12253 3071 12311 3077
rect 13262 3068 13268 3120
rect 13320 3068 13326 3120
rect 13722 3068 13728 3120
rect 13780 3108 13786 3120
rect 14277 3111 14335 3117
rect 14277 3108 14289 3111
rect 13780 3080 14289 3108
rect 13780 3068 13786 3080
rect 14277 3077 14289 3080
rect 14323 3077 14335 3111
rect 14277 3071 14335 3077
rect 8941 3043 8999 3049
rect 6052 3012 8892 3040
rect 6052 3000 6058 3012
rect 8864 2972 8892 3012
rect 8941 3009 8953 3043
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9858 3040 9864 3052
rect 9079 3012 9864 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9048 2972 9076 3003
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10134 3000 10140 3052
rect 10192 3000 10198 3052
rect 10412 3043 10470 3049
rect 10412 3009 10424 3043
rect 10458 3038 10470 3043
rect 10502 3038 10508 3052
rect 10458 3010 10508 3038
rect 10458 3009 10470 3010
rect 10412 3003 10470 3009
rect 10502 3000 10508 3010
rect 10560 3040 10566 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10560 3012 10885 3040
rect 10560 3000 10566 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11756 3012 11989 3040
rect 11756 3000 11762 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 13817 3043 13875 3049
rect 13817 3009 13829 3043
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3040 14243 3043
rect 14384 3040 14412 3148
rect 14231 3012 14412 3040
rect 14231 3009 14243 3012
rect 14185 3003 14243 3009
rect 8864 2944 9076 2972
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 10100 2944 10241 2972
rect 10100 2932 10106 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 10229 2935 10287 2941
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2972 10379 2975
rect 10778 2972 10784 2984
rect 10367 2944 10784 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 10778 2932 10784 2944
rect 10836 2972 10842 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 10836 2944 11253 2972
rect 10836 2932 10842 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 13832 2972 13860 3003
rect 12400 2944 13860 2972
rect 14016 2972 14044 3003
rect 14550 2972 14556 2984
rect 14016 2944 14556 2972
rect 12400 2932 12406 2944
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8665 2907 8723 2913
rect 8665 2904 8677 2907
rect 8352 2876 8677 2904
rect 8352 2864 8358 2876
rect 8665 2873 8677 2876
rect 8711 2873 8723 2907
rect 8665 2867 8723 2873
rect 8754 2864 8760 2916
rect 8812 2904 8818 2916
rect 9125 2907 9183 2913
rect 9125 2904 9137 2907
rect 8812 2876 9137 2904
rect 8812 2864 8818 2876
rect 9125 2873 9137 2876
rect 9171 2904 9183 2907
rect 14093 2907 14151 2913
rect 14093 2904 14105 2907
rect 9171 2876 11008 2904
rect 9171 2873 9183 2876
rect 9125 2867 9183 2873
rect 3786 2796 3792 2848
rect 3844 2836 3850 2848
rect 10226 2836 10232 2848
rect 3844 2808 10232 2836
rect 3844 2796 3850 2808
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 10980 2836 11008 2876
rect 13280 2876 14105 2904
rect 13280 2836 13308 2876
rect 14093 2873 14105 2876
rect 14139 2873 14151 2907
rect 14093 2867 14151 2873
rect 10980 2808 13308 2836
rect 13354 2796 13360 2848
rect 13412 2836 13418 2848
rect 13725 2839 13783 2845
rect 13725 2836 13737 2839
rect 13412 2808 13737 2836
rect 13412 2796 13418 2808
rect 13725 2805 13737 2808
rect 13771 2805 13783 2839
rect 13725 2799 13783 2805
rect 1104 2746 14812 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 14812 2746
rect 1104 2672 14812 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 6270 2632 6276 2644
rect 1627 2604 6276 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 6270 2592 6276 2604
rect 6328 2632 6334 2644
rect 6328 2604 6592 2632
rect 6328 2592 6334 2604
rect 4062 2524 4068 2576
rect 4120 2564 4126 2576
rect 6564 2564 6592 2604
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9217 2635 9275 2641
rect 9217 2632 9229 2635
rect 9088 2604 9229 2632
rect 9088 2592 9094 2604
rect 9217 2601 9229 2604
rect 9263 2601 9275 2635
rect 12897 2635 12955 2641
rect 12897 2632 12909 2635
rect 9217 2595 9275 2601
rect 9876 2604 12909 2632
rect 9674 2564 9680 2576
rect 4120 2536 5948 2564
rect 6564 2536 9680 2564
rect 4120 2524 4126 2536
rect 1670 2456 1676 2508
rect 1728 2496 1734 2508
rect 3053 2499 3111 2505
rect 3053 2496 3065 2499
rect 1728 2468 3065 2496
rect 1728 2456 1734 2468
rect 3053 2465 3065 2468
rect 3099 2465 3111 2499
rect 3053 2459 3111 2465
rect 3329 2499 3387 2505
rect 3329 2465 3341 2499
rect 3375 2496 3387 2499
rect 5810 2496 5816 2508
rect 3375 2468 5816 2496
rect 3375 2465 3387 2468
rect 3329 2459 3387 2465
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 5920 2496 5948 2536
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 9876 2496 9904 2604
rect 12897 2601 12909 2604
rect 12943 2632 12955 2635
rect 12943 2604 13492 2632
rect 12943 2601 12955 2604
rect 12897 2595 12955 2601
rect 11514 2524 11520 2576
rect 11572 2524 11578 2576
rect 11790 2524 11796 2576
rect 11848 2564 11854 2576
rect 13354 2564 13360 2576
rect 11848 2536 13360 2564
rect 11848 2524 11854 2536
rect 13354 2524 13360 2536
rect 13412 2524 13418 2576
rect 5920 2468 9904 2496
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10008 2468 10701 2496
rect 10008 2456 10014 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 13262 2456 13268 2508
rect 13320 2456 13326 2508
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 8018 2428 8024 2440
rect 4212 2400 8024 2428
rect 4212 2388 4218 2400
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 9033 2431 9091 2437
rect 9033 2428 9045 2431
rect 8168 2400 9045 2428
rect 8168 2388 8174 2400
rect 9033 2397 9045 2400
rect 9079 2397 9091 2431
rect 9033 2391 9091 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9398 2388 9404 2440
rect 9456 2388 9462 2440
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 9600 2400 11069 2428
rect 2498 2320 2504 2372
rect 2556 2320 2562 2372
rect 7374 2320 7380 2372
rect 7432 2360 7438 2372
rect 8757 2363 8815 2369
rect 8757 2360 8769 2363
rect 7432 2332 8769 2360
rect 7432 2320 7438 2332
rect 8757 2329 8769 2332
rect 8803 2360 8815 2363
rect 9493 2363 9551 2369
rect 9493 2360 9505 2363
rect 8803 2332 9505 2360
rect 8803 2329 8815 2332
rect 8757 2323 8815 2329
rect 9493 2329 9505 2332
rect 9539 2329 9551 2363
rect 9493 2323 9551 2329
rect 9600 2304 9628 2400
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 13464 2437 13492 2604
rect 13630 2592 13636 2644
rect 13688 2632 13694 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 13688 2604 14289 2632
rect 13688 2592 13694 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 14277 2595 14335 2601
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11756 2400 11989 2428
rect 11756 2388 11762 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 13725 2431 13783 2437
rect 13725 2428 13737 2431
rect 13596 2400 13737 2428
rect 13596 2388 13602 2400
rect 13725 2397 13737 2400
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 9815 2332 10548 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 9582 2252 9588 2304
rect 9640 2252 9646 2304
rect 10134 2252 10140 2304
rect 10192 2252 10198 2304
rect 10520 2292 10548 2332
rect 10870 2320 10876 2372
rect 10928 2320 10934 2372
rect 10962 2320 10968 2372
rect 11020 2320 11026 2372
rect 14476 2360 14504 2391
rect 12544 2332 14504 2360
rect 10980 2292 11008 2320
rect 12544 2304 12572 2332
rect 10520 2264 11008 2292
rect 11238 2252 11244 2304
rect 11296 2252 11302 2304
rect 12526 2252 12532 2304
rect 12584 2252 12590 2304
rect 13630 2252 13636 2304
rect 13688 2252 13694 2304
rect 13906 2252 13912 2304
rect 13964 2252 13970 2304
rect 1104 2202 14812 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 14812 2202
rect 1104 2128 14812 2150
rect 1210 2048 1216 2100
rect 1268 2088 1274 2100
rect 12526 2088 12532 2100
rect 1268 2060 12532 2088
rect 1268 2048 1274 2060
rect 12526 2048 12532 2060
rect 12584 2048 12590 2100
rect 8018 1980 8024 2032
rect 8076 2020 8082 2032
rect 9122 2020 9128 2032
rect 8076 1992 9128 2020
rect 8076 1980 8082 1992
rect 9122 1980 9128 1992
rect 9180 2020 9186 2032
rect 10134 2020 10140 2032
rect 9180 1992 10140 2020
rect 9180 1980 9186 1992
rect 10134 1980 10140 1992
rect 10192 2020 10198 2032
rect 13170 2020 13176 2032
rect 10192 1992 13176 2020
rect 10192 1980 10198 1992
rect 13170 1980 13176 1992
rect 13228 1980 13234 2032
rect 4706 1844 4712 1896
rect 4764 1884 4770 1896
rect 9582 1884 9588 1896
rect 4764 1856 9588 1884
rect 4764 1844 4770 1856
rect 9582 1844 9588 1856
rect 9640 1844 9646 1896
rect 6730 1640 6736 1692
rect 6788 1680 6794 1692
rect 11238 1680 11244 1692
rect 6788 1652 11244 1680
rect 6788 1640 6794 1652
rect 11238 1640 11244 1652
rect 11296 1640 11302 1692
<< via1 >>
rect 6644 15920 6696 15972
rect 14740 15920 14792 15972
rect 664 15852 716 15904
rect 9680 15852 9732 15904
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 14556 15648 14608 15700
rect 14372 15580 14424 15632
rect 8208 15512 8260 15564
rect 10600 15512 10652 15564
rect 13728 15512 13780 15564
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 4896 15444 4948 15496
rect 8944 15444 8996 15496
rect 9128 15444 9180 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 6000 15376 6052 15428
rect 10140 15376 10192 15428
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 15292 15376 15344 15428
rect 2412 15351 2464 15360
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 3240 15308 3292 15360
rect 5080 15308 5132 15360
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 6828 15308 6880 15317
rect 12440 15351 12492 15360
rect 12440 15317 12449 15351
rect 12449 15317 12483 15351
rect 12483 15317 12492 15351
rect 12440 15308 12492 15317
rect 13176 15308 13228 15360
rect 13912 15351 13964 15360
rect 13912 15317 13921 15351
rect 13921 15317 13955 15351
rect 13955 15317 13964 15351
rect 13912 15308 13964 15317
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 2412 15104 2464 15156
rect 3884 15104 3936 15156
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 6552 15104 6604 15156
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 4344 15036 4396 15088
rect 6920 15036 6972 15088
rect 8116 15104 8168 15156
rect 10784 15104 10836 15156
rect 14280 15104 14332 15156
rect 14924 15104 14976 15156
rect 5356 14968 5408 15020
rect 5908 14968 5960 15020
rect 3240 14900 3292 14952
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 4528 14943 4580 14952
rect 4528 14909 4537 14943
rect 4537 14909 4571 14943
rect 4571 14909 4580 14943
rect 4528 14900 4580 14909
rect 3148 14832 3200 14884
rect 5172 14832 5224 14884
rect 5724 14832 5776 14884
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 7288 15036 7340 15088
rect 10692 15036 10744 15088
rect 10876 15036 10928 15088
rect 10508 14968 10560 15020
rect 10968 14968 11020 15020
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 8484 14900 8536 14952
rect 14464 15011 14516 15020
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 1492 14764 1544 14816
rect 1860 14764 1912 14816
rect 3240 14764 3292 14816
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 5632 14807 5684 14816
rect 5632 14773 5641 14807
rect 5641 14773 5675 14807
rect 5675 14773 5684 14807
rect 5632 14764 5684 14773
rect 7104 14764 7156 14816
rect 8392 14764 8444 14816
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 10416 14764 10468 14816
rect 11060 14832 11112 14884
rect 12348 14832 12400 14884
rect 12532 14832 12584 14884
rect 11520 14764 11572 14816
rect 11612 14807 11664 14816
rect 11612 14773 11621 14807
rect 11621 14773 11655 14807
rect 11655 14773 11664 14807
rect 11612 14764 11664 14773
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 940 14492 992 14544
rect 4712 14560 4764 14612
rect 5264 14560 5316 14612
rect 1952 14424 2004 14476
rect 4344 14492 4396 14544
rect 7472 14560 7524 14612
rect 10784 14560 10836 14612
rect 8300 14492 8352 14544
rect 3792 14424 3844 14476
rect 5724 14467 5776 14476
rect 5724 14433 5733 14467
rect 5733 14433 5767 14467
rect 5767 14433 5776 14467
rect 5724 14424 5776 14433
rect 12348 14492 12400 14544
rect 4160 14356 4212 14408
rect 1860 14288 1912 14340
rect 1768 14263 1820 14272
rect 1768 14229 1777 14263
rect 1777 14229 1811 14263
rect 1811 14229 1820 14263
rect 1768 14220 1820 14229
rect 2964 14220 3016 14272
rect 4436 14220 4488 14272
rect 4620 14220 4672 14272
rect 5264 14220 5316 14272
rect 13268 14424 13320 14476
rect 6552 14356 6604 14408
rect 8760 14356 8812 14408
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 10968 14356 11020 14408
rect 12348 14356 12400 14408
rect 9220 14331 9272 14340
rect 9220 14297 9229 14331
rect 9229 14297 9263 14331
rect 9263 14297 9272 14331
rect 9220 14288 9272 14297
rect 13912 14288 13964 14340
rect 6092 14220 6144 14272
rect 9864 14220 9916 14272
rect 9956 14220 10008 14272
rect 10876 14220 10928 14272
rect 13544 14220 13596 14272
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14464 14220 14516 14229
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 2780 13948 2832 14000
rect 3608 13948 3660 14000
rect 4160 14016 4212 14068
rect 6828 14016 6880 14068
rect 4620 13948 4672 14000
rect 4804 13948 4856 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 4344 13923 4396 13932
rect 4344 13889 4353 13923
rect 4353 13889 4387 13923
rect 4387 13889 4396 13923
rect 4344 13880 4396 13889
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 4712 13880 4764 13932
rect 5724 13880 5776 13932
rect 8484 14059 8536 14068
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 11336 14016 11388 14068
rect 12532 14016 12584 14068
rect 9036 13948 9088 14000
rect 9588 13948 9640 14000
rect 9680 13948 9732 14000
rect 9864 13880 9916 13932
rect 12348 13880 12400 13932
rect 13544 13948 13596 14000
rect 13820 13948 13872 14000
rect 14004 13991 14056 14000
rect 14004 13957 14013 13991
rect 14013 13957 14047 13991
rect 14047 13957 14056 13991
rect 14004 13948 14056 13957
rect 1768 13812 1820 13864
rect 3516 13812 3568 13864
rect 5356 13812 5408 13864
rect 6736 13812 6788 13864
rect 8300 13812 8352 13864
rect 9312 13812 9364 13864
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 13452 13923 13504 13932
rect 13452 13889 13461 13923
rect 13461 13889 13495 13923
rect 13495 13889 13504 13923
rect 13452 13880 13504 13889
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 6000 13787 6052 13796
rect 6000 13753 6009 13787
rect 6009 13753 6043 13787
rect 6043 13753 6052 13787
rect 6000 13744 6052 13753
rect 8024 13744 8076 13796
rect 1676 13676 1728 13728
rect 2136 13676 2188 13728
rect 3976 13676 4028 13728
rect 4620 13676 4672 13728
rect 5356 13676 5408 13728
rect 5448 13676 5500 13728
rect 7564 13676 7616 13728
rect 8300 13719 8352 13728
rect 8300 13685 8309 13719
rect 8309 13685 8343 13719
rect 8343 13685 8352 13719
rect 8300 13676 8352 13685
rect 9404 13676 9456 13728
rect 11152 13676 11204 13728
rect 11796 13676 11848 13728
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 15660 13812 15712 13864
rect 13544 13676 13596 13728
rect 14096 13676 14148 13728
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 4068 13515 4120 13524
rect 4068 13481 4077 13515
rect 4077 13481 4111 13515
rect 4111 13481 4120 13515
rect 4068 13472 4120 13481
rect 4620 13472 4672 13524
rect 6460 13472 6512 13524
rect 5540 13404 5592 13456
rect 3516 13336 3568 13388
rect 8116 13404 8168 13456
rect 8208 13404 8260 13456
rect 8484 13404 8536 13456
rect 9036 13472 9088 13524
rect 9772 13404 9824 13456
rect 11152 13404 11204 13456
rect 1124 13200 1176 13252
rect 2872 13268 2924 13320
rect 3608 13311 3660 13320
rect 3608 13277 3617 13311
rect 3617 13277 3651 13311
rect 3651 13277 3660 13311
rect 3608 13268 3660 13277
rect 8576 13336 8628 13388
rect 8944 13336 8996 13388
rect 5448 13268 5500 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 7380 13268 7432 13320
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 9404 13268 9456 13320
rect 11428 13268 11480 13320
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 1308 13132 1360 13184
rect 4344 13243 4396 13252
rect 4344 13209 4353 13243
rect 4353 13209 4387 13243
rect 4387 13209 4396 13243
rect 4344 13200 4396 13209
rect 5264 13200 5316 13252
rect 5356 13200 5408 13252
rect 8300 13200 8352 13252
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 4252 13132 4304 13141
rect 4712 13132 4764 13184
rect 6736 13132 6788 13184
rect 9036 13132 9088 13184
rect 9864 13132 9916 13184
rect 10784 13243 10836 13252
rect 10784 13209 10793 13243
rect 10793 13209 10827 13243
rect 10827 13209 10836 13243
rect 10784 13200 10836 13209
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 14648 13268 14700 13320
rect 11428 13175 11480 13184
rect 11428 13141 11437 13175
rect 11437 13141 11471 13175
rect 11471 13141 11480 13175
rect 11428 13132 11480 13141
rect 12256 13200 12308 13252
rect 12348 13243 12400 13252
rect 12348 13209 12357 13243
rect 12357 13209 12391 13243
rect 12391 13209 12400 13243
rect 12348 13200 12400 13209
rect 12440 13200 12492 13252
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 3056 12928 3108 12980
rect 3516 12928 3568 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 13268 12928 13320 12980
rect 14096 12971 14148 12980
rect 14096 12937 14105 12971
rect 14105 12937 14139 12971
rect 14139 12937 14148 12971
rect 14096 12928 14148 12937
rect 2412 12860 2464 12912
rect 2504 12792 2556 12844
rect 1216 12724 1268 12776
rect 3148 12724 3200 12776
rect 6276 12860 6328 12912
rect 5724 12792 5776 12844
rect 6000 12835 6052 12844
rect 6000 12801 6009 12835
rect 6009 12801 6043 12835
rect 6043 12801 6052 12835
rect 6000 12792 6052 12801
rect 6184 12835 6236 12844
rect 6184 12801 6193 12835
rect 6193 12801 6227 12835
rect 6227 12801 6236 12835
rect 6184 12792 6236 12801
rect 6460 12792 6512 12844
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 8300 12860 8352 12912
rect 9220 12860 9272 12912
rect 12348 12860 12400 12912
rect 8760 12835 8812 12844
rect 8760 12801 8767 12835
rect 8767 12801 8801 12835
rect 8801 12801 8812 12835
rect 8760 12792 8812 12801
rect 9128 12792 9180 12844
rect 4252 12724 4304 12776
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 4896 12656 4948 12708
rect 6000 12656 6052 12708
rect 6644 12656 6696 12708
rect 6736 12656 6788 12708
rect 7564 12656 7616 12708
rect 8208 12588 8260 12640
rect 9312 12724 9364 12776
rect 11152 12724 11204 12776
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 14096 12792 14148 12844
rect 9496 12656 9548 12708
rect 9588 12656 9640 12708
rect 11704 12656 11756 12708
rect 12256 12699 12308 12708
rect 12256 12665 12265 12699
rect 12265 12665 12299 12699
rect 12299 12665 12308 12699
rect 12256 12656 12308 12665
rect 9128 12588 9180 12640
rect 9312 12588 9364 12640
rect 11244 12588 11296 12640
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 14832 12588 14884 12640
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 3424 12384 3476 12436
rect 4528 12384 4580 12436
rect 5448 12384 5500 12436
rect 8392 12384 8444 12436
rect 9588 12384 9640 12436
rect 10876 12384 10928 12436
rect 8116 12316 8168 12368
rect 8300 12316 8352 12368
rect 8852 12316 8904 12368
rect 10140 12316 10192 12368
rect 11980 12384 12032 12436
rect 13268 12427 13320 12436
rect 13268 12393 13277 12427
rect 13277 12393 13311 12427
rect 13311 12393 13320 12427
rect 13268 12384 13320 12393
rect 15016 12316 15068 12368
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 4528 12248 4580 12300
rect 5632 12248 5684 12300
rect 6736 12248 6788 12300
rect 6552 12180 6604 12232
rect 8392 12180 8444 12232
rect 9680 12248 9732 12300
rect 10324 12180 10376 12232
rect 10968 12180 11020 12232
rect 11520 12180 11572 12232
rect 12532 12180 12584 12232
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 4712 12112 4764 12164
rect 6092 12155 6144 12164
rect 6092 12121 6101 12155
rect 6101 12121 6135 12155
rect 6135 12121 6144 12155
rect 6092 12112 6144 12121
rect 6920 12112 6972 12164
rect 7748 12112 7800 12164
rect 8208 12155 8260 12164
rect 8208 12121 8217 12155
rect 8217 12121 8251 12155
rect 8251 12121 8260 12155
rect 8208 12112 8260 12121
rect 8576 12112 8628 12164
rect 9312 12112 9364 12164
rect 3608 12044 3660 12096
rect 10876 12112 10928 12164
rect 13268 12180 13320 12232
rect 13452 12155 13504 12164
rect 13452 12121 13461 12155
rect 13461 12121 13495 12155
rect 13495 12121 13504 12155
rect 13452 12112 13504 12121
rect 10140 12044 10192 12096
rect 10508 12044 10560 12096
rect 10968 12044 11020 12096
rect 11796 12087 11848 12096
rect 11796 12053 11805 12087
rect 11805 12053 11839 12087
rect 11839 12053 11848 12087
rect 11796 12044 11848 12053
rect 12992 12044 13044 12096
rect 13544 12044 13596 12096
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 2964 11840 3016 11892
rect 8392 11840 8444 11892
rect 8576 11840 8628 11892
rect 11520 11840 11572 11892
rect 4712 11815 4764 11824
rect 4712 11781 4721 11815
rect 4721 11781 4755 11815
rect 4755 11781 4764 11815
rect 4712 11772 4764 11781
rect 4896 11772 4948 11824
rect 5172 11815 5224 11824
rect 5172 11781 5181 11815
rect 5181 11781 5215 11815
rect 5215 11781 5224 11815
rect 5172 11772 5224 11781
rect 5632 11772 5684 11824
rect 9680 11772 9732 11824
rect 10048 11772 10100 11824
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 13452 11840 13504 11892
rect 14924 11840 14976 11892
rect 15200 11840 15252 11892
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 3424 11704 3476 11756
rect 3608 11704 3660 11756
rect 4252 11704 4304 11756
rect 5448 11704 5500 11756
rect 4712 11636 4764 11688
rect 5540 11636 5592 11688
rect 4068 11568 4120 11620
rect 6276 11704 6328 11756
rect 6644 11704 6696 11756
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 8300 11704 8352 11756
rect 11520 11704 11572 11756
rect 11704 11747 11756 11756
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 13820 11772 13872 11824
rect 14280 11704 14332 11756
rect 7748 11636 7800 11688
rect 8576 11636 8628 11688
rect 8760 11679 8812 11688
rect 8760 11645 8778 11679
rect 8778 11645 8812 11679
rect 8760 11636 8812 11645
rect 8852 11679 8904 11688
rect 8852 11645 8861 11679
rect 8861 11645 8895 11679
rect 8895 11645 8904 11679
rect 8852 11636 8904 11645
rect 2964 11500 3016 11552
rect 3424 11543 3476 11552
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 3424 11500 3476 11509
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 5540 11500 5592 11552
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 6552 11500 6604 11552
rect 8300 11500 8352 11552
rect 8576 11543 8628 11552
rect 8576 11509 8585 11543
rect 8585 11509 8619 11543
rect 8619 11509 8628 11543
rect 8576 11500 8628 11509
rect 8852 11500 8904 11552
rect 9312 11679 9364 11688
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 9312 11636 9364 11645
rect 9588 11679 9640 11688
rect 9588 11645 9597 11679
rect 9597 11645 9631 11679
rect 9631 11645 9640 11679
rect 9588 11636 9640 11645
rect 11428 11568 11480 11620
rect 10692 11500 10744 11552
rect 13452 11568 13504 11620
rect 12900 11500 12952 11552
rect 13268 11500 13320 11552
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 1492 11296 1544 11348
rect 2596 11296 2648 11348
rect 2780 11296 2832 11348
rect 3608 11296 3660 11348
rect 3148 11160 3200 11212
rect 3700 11160 3752 11212
rect 5172 11296 5224 11348
rect 5540 11296 5592 11348
rect 7012 11296 7064 11348
rect 3976 11271 4028 11280
rect 3976 11237 3985 11271
rect 3985 11237 4019 11271
rect 4019 11237 4028 11271
rect 3976 11228 4028 11237
rect 4344 11228 4396 11280
rect 7656 11228 7708 11280
rect 7840 11228 7892 11280
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 1584 11092 1636 11144
rect 4252 11092 4304 11144
rect 4160 11024 4212 11076
rect 4896 11160 4948 11212
rect 5356 11160 5408 11212
rect 6460 11024 6512 11076
rect 7012 11160 7064 11212
rect 7196 11160 7248 11212
rect 8576 11160 8628 11212
rect 7288 11092 7340 11144
rect 8300 11092 8352 11144
rect 9312 11228 9364 11280
rect 11152 11228 11204 11280
rect 12900 11228 12952 11280
rect 13084 11228 13136 11280
rect 11520 11160 11572 11212
rect 12440 11203 12492 11212
rect 12440 11169 12449 11203
rect 12449 11169 12483 11203
rect 12483 11169 12492 11203
rect 12440 11160 12492 11169
rect 12532 11160 12584 11212
rect 12808 11160 12860 11212
rect 10968 11092 11020 11144
rect 12992 11092 13044 11144
rect 4620 10956 4672 11008
rect 4896 10956 4948 11008
rect 6184 10956 6236 11008
rect 6644 10956 6696 11008
rect 7012 11024 7064 11076
rect 7840 11024 7892 11076
rect 8484 11067 8536 11076
rect 8484 11033 8493 11067
rect 8493 11033 8527 11067
rect 8527 11033 8536 11067
rect 8484 11024 8536 11033
rect 12256 11024 12308 11076
rect 12808 11067 12860 11076
rect 12808 11033 12817 11067
rect 12817 11033 12851 11067
rect 12851 11033 12860 11067
rect 12808 11024 12860 11033
rect 13268 11092 13320 11144
rect 13544 11024 13596 11076
rect 13636 11024 13688 11076
rect 13820 11024 13872 11076
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 7104 10956 7156 11008
rect 7288 10956 7340 11008
rect 12992 10956 13044 11008
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 2780 10616 2832 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 4712 10752 4764 10804
rect 5264 10795 5316 10804
rect 5264 10761 5273 10795
rect 5273 10761 5307 10795
rect 5307 10761 5316 10795
rect 5264 10752 5316 10761
rect 6368 10752 6420 10804
rect 6644 10752 6696 10804
rect 7288 10752 7340 10804
rect 7564 10752 7616 10804
rect 9036 10752 9088 10804
rect 10324 10752 10376 10804
rect 12532 10752 12584 10804
rect 13728 10752 13780 10804
rect 5908 10684 5960 10736
rect 6920 10684 6972 10736
rect 4436 10616 4488 10668
rect 5816 10616 5868 10668
rect 6368 10616 6420 10668
rect 6828 10616 6880 10668
rect 9864 10684 9916 10736
rect 10692 10684 10744 10736
rect 12348 10727 12400 10736
rect 12348 10693 12357 10727
rect 12357 10693 12391 10727
rect 12391 10693 12400 10727
rect 12348 10684 12400 10693
rect 7748 10616 7800 10668
rect 4712 10548 4764 10600
rect 4896 10591 4948 10600
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 6276 10548 6328 10600
rect 6736 10548 6788 10600
rect 1676 10480 1728 10532
rect 8852 10548 8904 10600
rect 9220 10616 9272 10668
rect 10600 10616 10652 10668
rect 11520 10616 11572 10668
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 12532 10659 12584 10668
rect 12532 10625 12541 10659
rect 12541 10625 12575 10659
rect 12575 10625 12584 10659
rect 12532 10616 12584 10625
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 13268 10616 13320 10668
rect 13452 10659 13504 10668
rect 13452 10625 13461 10659
rect 13461 10625 13495 10659
rect 13495 10625 13504 10659
rect 13452 10616 13504 10625
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 12624 10548 12676 10600
rect 13636 10616 13688 10668
rect 14280 10616 14332 10668
rect 2780 10455 2832 10464
rect 2780 10421 2789 10455
rect 2789 10421 2823 10455
rect 2823 10421 2832 10455
rect 2780 10412 2832 10421
rect 3424 10412 3476 10464
rect 5448 10412 5500 10464
rect 6368 10412 6420 10464
rect 6736 10412 6788 10464
rect 10508 10480 10560 10532
rect 12532 10523 12584 10532
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 8484 10412 8536 10464
rect 11520 10412 11572 10464
rect 12440 10412 12492 10464
rect 14648 10548 14700 10600
rect 15016 10412 15068 10464
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 2228 10208 2280 10260
rect 2964 10208 3016 10260
rect 3240 10208 3292 10260
rect 4160 10208 4212 10260
rect 5632 10208 5684 10260
rect 3332 10183 3384 10192
rect 3332 10149 3341 10183
rect 3341 10149 3375 10183
rect 3375 10149 3384 10183
rect 3332 10140 3384 10149
rect 4528 10140 4580 10192
rect 5356 10140 5408 10192
rect 6092 10140 6144 10192
rect 3884 10072 3936 10124
rect 5540 10072 5592 10124
rect 6920 10208 6972 10260
rect 10508 10208 10560 10260
rect 9496 10140 9548 10192
rect 8024 10072 8076 10124
rect 8484 10072 8536 10124
rect 11060 10072 11112 10124
rect 4160 10004 4212 10056
rect 5264 10004 5316 10056
rect 6276 10004 6328 10056
rect 3148 9936 3200 9988
rect 6552 9936 6604 9988
rect 8392 9936 8444 9988
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 11520 10004 11572 10056
rect 11704 10140 11756 10192
rect 12624 10140 12676 10192
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 10048 9936 10100 9988
rect 10692 9936 10744 9988
rect 11060 9936 11112 9988
rect 11244 9936 11296 9988
rect 12624 10004 12676 10056
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13452 10208 13504 10260
rect 13360 10072 13412 10124
rect 13452 9936 13504 9988
rect 13820 9936 13872 9988
rect 2780 9868 2832 9920
rect 5540 9868 5592 9920
rect 5908 9868 5960 9920
rect 6736 9868 6788 9920
rect 6828 9868 6880 9920
rect 8208 9868 8260 9920
rect 9220 9868 9272 9920
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 9864 9911 9916 9920
rect 9864 9877 9873 9911
rect 9873 9877 9907 9911
rect 9907 9877 9916 9911
rect 9864 9868 9916 9877
rect 11704 9868 11756 9920
rect 11796 9868 11848 9920
rect 13084 9868 13136 9920
rect 14464 9911 14516 9920
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 4252 9664 4304 9716
rect 4436 9664 4488 9716
rect 848 9528 900 9580
rect 1492 9528 1544 9580
rect 1308 9460 1360 9512
rect 2228 9460 2280 9512
rect 1492 9392 1544 9444
rect 2596 9460 2648 9512
rect 3056 9596 3108 9648
rect 5356 9664 5408 9716
rect 5632 9664 5684 9716
rect 6092 9664 6144 9716
rect 6460 9664 6512 9716
rect 6736 9707 6788 9716
rect 6736 9673 6745 9707
rect 6745 9673 6779 9707
rect 6779 9673 6788 9707
rect 6736 9664 6788 9673
rect 2780 9528 2832 9580
rect 3332 9528 3384 9580
rect 3424 9528 3476 9580
rect 3608 9528 3660 9580
rect 4160 9528 4212 9580
rect 6184 9596 6236 9648
rect 6368 9639 6420 9648
rect 6368 9605 6377 9639
rect 6377 9605 6411 9639
rect 6411 9605 6420 9639
rect 6368 9596 6420 9605
rect 8024 9664 8076 9716
rect 14004 9664 14056 9716
rect 4068 9460 4120 9512
rect 2872 9435 2924 9444
rect 2872 9401 2881 9435
rect 2881 9401 2915 9435
rect 2915 9401 2924 9435
rect 2872 9392 2924 9401
rect 3056 9324 3108 9376
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 4068 9324 4120 9376
rect 6000 9528 6052 9580
rect 6276 9528 6328 9580
rect 8944 9596 8996 9648
rect 9772 9596 9824 9648
rect 10324 9596 10376 9648
rect 12072 9596 12124 9648
rect 14280 9596 14332 9648
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 5448 9460 5500 9512
rect 5908 9460 5960 9512
rect 6460 9460 6512 9512
rect 8024 9528 8076 9580
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 4436 9392 4488 9444
rect 8116 9460 8168 9512
rect 8208 9460 8260 9512
rect 9312 9528 9364 9580
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 12440 9528 12492 9580
rect 12716 9571 12768 9580
rect 12716 9537 12725 9571
rect 12725 9537 12759 9571
rect 12759 9537 12768 9571
rect 12716 9528 12768 9537
rect 12808 9528 12860 9580
rect 11244 9460 11296 9512
rect 5080 9324 5132 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 7288 9324 7340 9376
rect 7748 9324 7800 9376
rect 8024 9324 8076 9376
rect 9312 9392 9364 9444
rect 13728 9528 13780 9580
rect 15292 9528 15344 9580
rect 12808 9392 12860 9444
rect 8576 9324 8628 9376
rect 8944 9324 8996 9376
rect 10232 9324 10284 9376
rect 10324 9324 10376 9376
rect 12072 9324 12124 9376
rect 12716 9324 12768 9376
rect 13268 9324 13320 9376
rect 13360 9324 13412 9376
rect 14188 9460 14240 9512
rect 13820 9324 13872 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 2228 9120 2280 9172
rect 2780 9120 2832 9172
rect 3424 9120 3476 9172
rect 3976 9120 4028 9172
rect 5356 9120 5408 9172
rect 5724 9120 5776 9172
rect 10140 9120 10192 9172
rect 10232 9120 10284 9172
rect 4436 9052 4488 9104
rect 7288 9052 7340 9104
rect 8024 9052 8076 9104
rect 8852 9052 8904 9104
rect 9128 9052 9180 9104
rect 5724 9027 5776 9036
rect 5724 8993 5733 9027
rect 5733 8993 5767 9027
rect 5767 8993 5776 9027
rect 5724 8984 5776 8993
rect 5908 8984 5960 9036
rect 4160 8916 4212 8968
rect 7472 8984 7524 9036
rect 7748 8984 7800 9036
rect 8208 8984 8260 9036
rect 8576 8984 8628 9036
rect 8668 8984 8720 9036
rect 10692 9052 10744 9104
rect 12440 9052 12492 9104
rect 6920 8916 6972 8968
rect 8760 8916 8812 8968
rect 8944 8916 8996 8968
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 4988 8848 5040 8900
rect 5724 8848 5776 8900
rect 6276 8848 6328 8900
rect 7840 8848 7892 8900
rect 8576 8848 8628 8900
rect 8668 8848 8720 8900
rect 11520 8916 11572 8968
rect 11888 8916 11940 8968
rect 12256 8916 12308 8968
rect 2596 8780 2648 8832
rect 3148 8780 3200 8832
rect 4436 8780 4488 8832
rect 4712 8780 4764 8832
rect 7656 8780 7708 8832
rect 8208 8780 8260 8832
rect 9680 8891 9732 8900
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 10140 8848 10192 8900
rect 13452 8916 13504 8968
rect 12992 8848 13044 8900
rect 9772 8780 9824 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 13544 8780 13596 8832
rect 14464 8823 14516 8832
rect 14464 8789 14473 8823
rect 14473 8789 14507 8823
rect 14507 8789 14516 8823
rect 14464 8780 14516 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 5540 8576 5592 8628
rect 5908 8576 5960 8628
rect 6000 8576 6052 8628
rect 9680 8576 9732 8628
rect 2320 8508 2372 8560
rect 6092 8508 6144 8560
rect 8024 8508 8076 8560
rect 6000 8440 6052 8492
rect 3056 8372 3108 8424
rect 3792 8415 3844 8424
rect 3792 8381 3801 8415
rect 3801 8381 3835 8415
rect 3835 8381 3844 8415
rect 3792 8372 3844 8381
rect 5172 8372 5224 8424
rect 5540 8372 5592 8424
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 6736 8440 6788 8492
rect 9036 8508 9088 8560
rect 10876 8576 10928 8628
rect 10968 8576 11020 8628
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 10232 8440 10284 8492
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 11612 8576 11664 8628
rect 12348 8576 12400 8628
rect 13728 8576 13780 8628
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 14096 8619 14148 8628
rect 14096 8585 14105 8619
rect 14105 8585 14139 8619
rect 14139 8585 14148 8619
rect 14096 8576 14148 8585
rect 11336 8508 11388 8560
rect 12440 8508 12492 8560
rect 13912 8440 13964 8492
rect 15200 8576 15252 8628
rect 7932 8372 7984 8424
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 10784 8372 10836 8424
rect 11152 8372 11204 8424
rect 11980 8372 12032 8424
rect 5264 8347 5316 8356
rect 5264 8313 5273 8347
rect 5273 8313 5307 8347
rect 5307 8313 5316 8347
rect 5264 8304 5316 8313
rect 5448 8304 5500 8356
rect 7564 8304 7616 8356
rect 8668 8304 8720 8356
rect 9956 8304 10008 8356
rect 1860 8236 1912 8288
rect 2228 8236 2280 8288
rect 4436 8236 4488 8288
rect 4896 8236 4948 8288
rect 5724 8236 5776 8288
rect 7196 8236 7248 8288
rect 9036 8236 9088 8288
rect 10232 8236 10284 8288
rect 12440 8372 12492 8424
rect 12532 8304 12584 8356
rect 13452 8304 13504 8356
rect 13912 8236 13964 8288
rect 14740 8236 14792 8288
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 4528 8075 4580 8084
rect 4528 8041 4537 8075
rect 4537 8041 4571 8075
rect 4571 8041 4580 8075
rect 4528 8032 4580 8041
rect 5080 8032 5132 8084
rect 1860 7828 1912 7880
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2320 7828 2372 7880
rect 2320 7735 2372 7744
rect 2320 7701 2329 7735
rect 2329 7701 2363 7735
rect 2363 7701 2372 7735
rect 2320 7692 2372 7701
rect 3700 7828 3752 7880
rect 3976 7828 4028 7880
rect 4436 7828 4488 7880
rect 4528 7828 4580 7880
rect 6644 7964 6696 8016
rect 9588 8032 9640 8084
rect 9772 8032 9824 8084
rect 10048 8032 10100 8084
rect 9036 7964 9088 8016
rect 9128 7964 9180 8016
rect 11888 8032 11940 8084
rect 14280 8032 14332 8084
rect 12440 7964 12492 8016
rect 5172 7896 5224 7948
rect 5724 7896 5776 7948
rect 6092 7896 6144 7948
rect 10048 7896 10100 7948
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 5356 7828 5408 7880
rect 6184 7828 6236 7880
rect 7104 7828 7156 7880
rect 7564 7828 7616 7880
rect 7840 7828 7892 7880
rect 9588 7828 9640 7880
rect 10140 7828 10192 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 4712 7760 4764 7812
rect 3700 7692 3752 7744
rect 3976 7735 4028 7744
rect 3976 7701 3985 7735
rect 3985 7701 4019 7735
rect 4019 7701 4028 7735
rect 3976 7692 4028 7701
rect 6000 7760 6052 7812
rect 6460 7760 6512 7812
rect 6644 7760 6696 7812
rect 13452 7760 13504 7812
rect 5356 7692 5408 7744
rect 5448 7692 5500 7744
rect 6184 7692 6236 7744
rect 10508 7692 10560 7744
rect 10968 7692 11020 7744
rect 11152 7692 11204 7744
rect 11888 7692 11940 7744
rect 12440 7692 12492 7744
rect 12624 7692 12676 7744
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 848 7488 900 7540
rect 2596 7488 2648 7540
rect 2964 7488 3016 7540
rect 4068 7488 4120 7540
rect 4344 7488 4396 7540
rect 5448 7488 5500 7540
rect 6460 7488 6512 7540
rect 6552 7488 6604 7540
rect 6736 7531 6788 7540
rect 6736 7497 6745 7531
rect 6745 7497 6779 7531
rect 6779 7497 6788 7531
rect 6736 7488 6788 7497
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 7380 7488 7432 7540
rect 10048 7531 10100 7540
rect 10048 7497 10057 7531
rect 10057 7497 10091 7531
rect 10091 7497 10100 7531
rect 10048 7488 10100 7497
rect 664 7352 716 7404
rect 848 7352 900 7404
rect 1768 7420 1820 7472
rect 3424 7420 3476 7472
rect 5908 7420 5960 7472
rect 2228 7352 2280 7404
rect 2504 7284 2556 7336
rect 2688 7284 2740 7336
rect 4160 7327 4212 7336
rect 4160 7293 4169 7327
rect 4169 7293 4203 7327
rect 4203 7293 4212 7327
rect 4160 7284 4212 7293
rect 4620 7284 4672 7336
rect 6460 7352 6512 7404
rect 10140 7420 10192 7472
rect 10600 7488 10652 7540
rect 10508 7463 10560 7472
rect 10508 7429 10517 7463
rect 10517 7429 10551 7463
rect 10551 7429 10560 7463
rect 10508 7420 10560 7429
rect 11796 7463 11848 7472
rect 11796 7429 11805 7463
rect 11805 7429 11839 7463
rect 11839 7429 11848 7463
rect 11796 7420 11848 7429
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 9864 7352 9916 7404
rect 10048 7352 10100 7404
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 11244 7352 11296 7404
rect 12900 7352 12952 7404
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 13912 7488 13964 7540
rect 14188 7488 14240 7540
rect 13452 7352 13504 7404
rect 13912 7352 13964 7404
rect 7104 7284 7156 7293
rect 7472 7284 7524 7336
rect 11428 7284 11480 7336
rect 11796 7284 11848 7336
rect 12348 7284 12400 7336
rect 5540 7216 5592 7268
rect 6092 7216 6144 7268
rect 7288 7216 7340 7268
rect 7380 7216 7432 7268
rect 12808 7216 12860 7268
rect 13636 7216 13688 7268
rect 14648 7216 14700 7268
rect 2320 7148 2372 7200
rect 3700 7148 3752 7200
rect 8484 7148 8536 7200
rect 8668 7148 8720 7200
rect 10140 7148 10192 7200
rect 12256 7148 12308 7200
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 2964 6944 3016 6996
rect 4896 6944 4948 6996
rect 4988 6944 5040 6996
rect 756 6876 808 6928
rect 3056 6851 3108 6860
rect 3056 6817 3065 6851
rect 3065 6817 3099 6851
rect 3099 6817 3108 6851
rect 3056 6808 3108 6817
rect 6460 6944 6512 6996
rect 9496 6944 9548 6996
rect 9588 6944 9640 6996
rect 11428 6987 11480 6996
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 14464 6944 14516 6996
rect 5540 6876 5592 6928
rect 5448 6808 5500 6860
rect 6092 6876 6144 6928
rect 8024 6876 8076 6928
rect 8208 6876 8260 6928
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 3608 6740 3660 6792
rect 3884 6740 3936 6792
rect 4252 6783 4304 6792
rect 4252 6749 4286 6783
rect 4286 6749 4304 6783
rect 4252 6740 4304 6749
rect 4896 6740 4948 6792
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 6460 6672 6512 6724
rect 8208 6672 8260 6724
rect 8760 6740 8812 6792
rect 9128 6672 9180 6724
rect 11888 6808 11940 6860
rect 12440 6808 12492 6860
rect 11428 6740 11480 6792
rect 12164 6783 12216 6792
rect 12164 6749 12173 6783
rect 12173 6749 12207 6783
rect 12207 6749 12216 6783
rect 12164 6740 12216 6749
rect 15108 6808 15160 6860
rect 11704 6672 11756 6724
rect 3884 6604 3936 6656
rect 4344 6604 4396 6656
rect 4436 6647 4488 6656
rect 4436 6613 4445 6647
rect 4445 6613 4479 6647
rect 4479 6613 4488 6647
rect 4436 6604 4488 6613
rect 4528 6604 4580 6656
rect 4712 6604 4764 6656
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 5632 6604 5684 6656
rect 7288 6604 7340 6656
rect 7932 6604 7984 6656
rect 9588 6647 9640 6656
rect 9588 6613 9597 6647
rect 9597 6613 9631 6647
rect 9631 6613 9640 6647
rect 9588 6604 9640 6613
rect 10876 6604 10928 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 3608 6400 3660 6452
rect 4160 6400 4212 6452
rect 3884 6332 3936 6384
rect 4252 6264 4304 6316
rect 4712 6264 4764 6316
rect 5264 6264 5316 6316
rect 5632 6400 5684 6452
rect 6828 6400 6880 6452
rect 5724 6332 5776 6384
rect 5908 6332 5960 6384
rect 5632 6264 5684 6316
rect 4528 6196 4580 6248
rect 6460 6307 6512 6316
rect 6460 6273 6469 6307
rect 6469 6273 6503 6307
rect 6503 6273 6512 6307
rect 6460 6264 6512 6273
rect 5908 6196 5960 6248
rect 7472 6332 7524 6384
rect 7656 6332 7708 6384
rect 8760 6375 8812 6384
rect 8760 6341 8769 6375
rect 8769 6341 8803 6375
rect 8803 6341 8812 6375
rect 8760 6332 8812 6341
rect 9588 6332 9640 6384
rect 10232 6375 10284 6384
rect 10232 6341 10241 6375
rect 10241 6341 10275 6375
rect 10275 6341 10284 6375
rect 10232 6332 10284 6341
rect 7104 6264 7156 6316
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7380 6264 7432 6316
rect 11796 6400 11848 6452
rect 13452 6400 13504 6452
rect 10416 6332 10468 6384
rect 12532 6332 12584 6384
rect 15292 6332 15344 6384
rect 6828 6196 6880 6248
rect 4068 6128 4120 6180
rect 4528 6060 4580 6112
rect 5448 6060 5500 6112
rect 5908 6060 5960 6112
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 7380 6128 7432 6180
rect 7840 6196 7892 6248
rect 8208 6196 8260 6248
rect 8392 6196 8444 6248
rect 8484 6239 8536 6248
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 10876 6264 10928 6316
rect 11888 6264 11940 6316
rect 12164 6264 12216 6316
rect 13636 6264 13688 6316
rect 11704 6196 11756 6248
rect 10416 6128 10468 6180
rect 6368 6060 6420 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 7196 6060 7248 6112
rect 7840 6060 7892 6112
rect 8024 6103 8076 6112
rect 8024 6069 8033 6103
rect 8033 6069 8067 6103
rect 8067 6069 8076 6103
rect 8024 6060 8076 6069
rect 10232 6060 10284 6112
rect 13636 6128 13688 6180
rect 14280 6060 14332 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 3240 5856 3292 5908
rect 4068 5856 4120 5908
rect 4160 5899 4212 5908
rect 4160 5865 4169 5899
rect 4169 5865 4203 5899
rect 4203 5865 4212 5899
rect 4160 5856 4212 5865
rect 5080 5856 5132 5908
rect 5632 5856 5684 5908
rect 6184 5856 6236 5908
rect 8300 5856 8352 5908
rect 8668 5856 8720 5908
rect 8852 5856 8904 5908
rect 10324 5856 10376 5908
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 3700 5788 3752 5840
rect 3792 5788 3844 5840
rect 3332 5763 3384 5772
rect 3332 5729 3341 5763
rect 3341 5729 3375 5763
rect 3375 5729 3384 5763
rect 3332 5720 3384 5729
rect 4528 5720 4580 5772
rect 1492 5652 1544 5704
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 3608 5652 3660 5704
rect 4068 5652 4120 5704
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 3884 5584 3936 5636
rect 4528 5584 4580 5636
rect 6736 5788 6788 5840
rect 11152 5788 11204 5840
rect 5632 5720 5684 5772
rect 5908 5720 5960 5772
rect 9956 5720 10008 5772
rect 10416 5720 10468 5772
rect 11704 5856 11756 5908
rect 13360 5856 13412 5908
rect 11520 5788 11572 5840
rect 11428 5720 11480 5772
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 14096 5831 14148 5840
rect 14096 5797 14105 5831
rect 14105 5797 14139 5831
rect 14139 5797 14148 5831
rect 14096 5788 14148 5797
rect 14188 5720 14240 5772
rect 14924 5720 14976 5772
rect 4988 5584 5040 5636
rect 5172 5584 5224 5636
rect 6644 5652 6696 5704
rect 7564 5652 7616 5704
rect 5448 5584 5500 5636
rect 7840 5652 7892 5704
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 3608 5516 3660 5568
rect 4160 5516 4212 5568
rect 4436 5516 4488 5568
rect 7748 5627 7800 5636
rect 7748 5593 7757 5627
rect 7757 5593 7791 5627
rect 7791 5593 7800 5627
rect 7748 5584 7800 5593
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9312 5652 9364 5704
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 9128 5584 9180 5636
rect 9680 5584 9732 5636
rect 7380 5516 7432 5568
rect 7472 5516 7524 5568
rect 8484 5516 8536 5568
rect 9312 5516 9364 5568
rect 9772 5516 9824 5568
rect 10324 5516 10376 5568
rect 10416 5516 10468 5568
rect 11612 5559 11664 5568
rect 11612 5525 11621 5559
rect 11621 5525 11655 5559
rect 11655 5525 11664 5559
rect 11612 5516 11664 5525
rect 11704 5516 11756 5568
rect 14096 5516 14148 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 4160 5312 4212 5364
rect 4620 5312 4672 5364
rect 4988 5312 5040 5364
rect 3424 5244 3476 5296
rect 5172 5244 5224 5296
rect 5356 5312 5408 5364
rect 6184 5312 6236 5364
rect 5724 5244 5776 5296
rect 6460 5244 6512 5296
rect 7196 5244 7248 5296
rect 8024 5244 8076 5296
rect 3332 5176 3384 5228
rect 4252 5176 4304 5228
rect 4528 5108 4580 5160
rect 4344 5040 4396 5092
rect 5816 5040 5868 5092
rect 6184 5083 6236 5092
rect 6184 5049 6193 5083
rect 6193 5049 6227 5083
rect 6227 5049 6236 5083
rect 6184 5040 6236 5049
rect 6736 5108 6788 5160
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 9864 5312 9916 5364
rect 12440 5312 12492 5364
rect 14188 5312 14240 5364
rect 11796 5287 11848 5296
rect 11796 5253 11805 5287
rect 11805 5253 11839 5287
rect 11839 5253 11848 5287
rect 11796 5244 11848 5253
rect 11980 5287 12032 5296
rect 11980 5253 11989 5287
rect 11989 5253 12023 5287
rect 12023 5253 12032 5287
rect 11980 5244 12032 5253
rect 12992 5244 13044 5296
rect 14280 5244 14332 5296
rect 8392 5108 8444 5160
rect 8852 5040 8904 5092
rect 9864 5151 9916 5160
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 11888 5176 11940 5228
rect 13820 5176 13872 5228
rect 11060 5108 11112 5160
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11336 5108 11388 5117
rect 13084 5108 13136 5160
rect 5908 4972 5960 5024
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 6368 4972 6420 5024
rect 6828 4972 6880 5024
rect 7380 4972 7432 5024
rect 9404 4972 9456 5024
rect 10232 4972 10284 5024
rect 10876 4972 10928 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 13268 4972 13320 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 1308 4768 1360 4820
rect 1032 4700 1084 4752
rect 5632 4768 5684 4820
rect 7380 4768 7432 4820
rect 7932 4768 7984 4820
rect 2504 4700 2556 4752
rect 3240 4700 3292 4752
rect 5356 4743 5408 4752
rect 5356 4709 5365 4743
rect 5365 4709 5399 4743
rect 5399 4709 5408 4743
rect 5356 4700 5408 4709
rect 9680 4768 9732 4820
rect 9772 4768 9824 4820
rect 10784 4768 10836 4820
rect 13360 4768 13412 4820
rect 14096 4768 14148 4820
rect 14464 4811 14516 4820
rect 14464 4777 14473 4811
rect 14473 4777 14507 4811
rect 14507 4777 14516 4811
rect 14464 4768 14516 4777
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 1860 4564 1912 4616
rect 2412 4632 2464 4684
rect 5540 4632 5592 4684
rect 8668 4700 8720 4752
rect 14004 4700 14056 4752
rect 6736 4632 6788 4684
rect 6828 4632 6880 4684
rect 8852 4632 8904 4684
rect 848 4496 900 4548
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 2964 4496 3016 4548
rect 1768 4428 1820 4480
rect 2504 4428 2556 4480
rect 3332 4428 3384 4480
rect 5632 4564 5684 4616
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 8392 4564 8444 4616
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9772 4632 9824 4684
rect 5448 4496 5500 4548
rect 6552 4496 6604 4548
rect 8944 4496 8996 4548
rect 9588 4607 9640 4616
rect 9588 4573 9597 4607
rect 9597 4573 9631 4607
rect 9631 4573 9640 4607
rect 9588 4564 9640 4573
rect 9772 4496 9824 4548
rect 4160 4428 4212 4480
rect 4988 4428 5040 4480
rect 6000 4428 6052 4480
rect 8484 4428 8536 4480
rect 8668 4428 8720 4480
rect 11060 4632 11112 4684
rect 11244 4632 11296 4684
rect 10692 4564 10744 4616
rect 10232 4428 10284 4480
rect 10876 4496 10928 4548
rect 11520 4564 11572 4616
rect 12164 4632 12216 4684
rect 11888 4564 11940 4616
rect 12256 4564 12308 4616
rect 11060 4496 11112 4548
rect 13452 4632 13504 4684
rect 12900 4564 12952 4616
rect 14832 4564 14884 4616
rect 13268 4496 13320 4548
rect 13176 4428 13228 4480
rect 13912 4471 13964 4480
rect 13912 4437 13921 4471
rect 13921 4437 13955 4471
rect 13955 4437 13964 4471
rect 13912 4428 13964 4437
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 2964 4267 3016 4276
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 3240 4224 3292 4276
rect 4988 4224 5040 4276
rect 5172 4224 5224 4276
rect 10692 4224 10744 4276
rect 11612 4224 11664 4276
rect 11796 4224 11848 4276
rect 2596 4156 2648 4208
rect 8484 4156 8536 4208
rect 12440 4224 12492 4276
rect 13912 4267 13964 4276
rect 13912 4233 13921 4267
rect 13921 4233 13955 4267
rect 13955 4233 13964 4267
rect 13912 4224 13964 4233
rect 12256 4156 12308 4208
rect 14188 4156 14240 4208
rect 6828 4088 6880 4140
rect 3056 4020 3108 4072
rect 9312 4088 9364 4140
rect 9588 4088 9640 4140
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7012 4020 7064 4029
rect 8392 4020 8444 4072
rect 10876 4020 10928 4072
rect 1584 3952 1636 4004
rect 5724 3995 5776 4004
rect 5724 3961 5733 3995
rect 5733 3961 5767 3995
rect 5767 3961 5776 3995
rect 5724 3952 5776 3961
rect 6552 3995 6604 4004
rect 6552 3961 6561 3995
rect 6561 3961 6595 3995
rect 6595 3961 6604 3995
rect 6552 3952 6604 3961
rect 9404 3952 9456 4004
rect 9588 3952 9640 4004
rect 11428 4088 11480 4140
rect 13360 4088 13412 4140
rect 11428 3952 11480 4004
rect 9680 3884 9732 3936
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 14096 4088 14148 4140
rect 14648 4156 14700 4208
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 13176 4020 13228 4029
rect 13452 3995 13504 4004
rect 13452 3961 13461 3995
rect 13461 3961 13495 3995
rect 13495 3961 13504 3995
rect 13452 3952 13504 3961
rect 13820 3952 13872 4004
rect 12532 3884 12584 3936
rect 13176 3884 13228 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 1400 3680 1452 3732
rect 2596 3680 2648 3732
rect 4804 3680 4856 3732
rect 7656 3723 7708 3732
rect 7656 3689 7665 3723
rect 7665 3689 7699 3723
rect 7699 3689 7708 3723
rect 7656 3680 7708 3689
rect 8944 3680 8996 3732
rect 9864 3680 9916 3732
rect 10324 3680 10376 3732
rect 4620 3612 4672 3664
rect 5264 3544 5316 3596
rect 7380 3612 7432 3664
rect 12992 3612 13044 3664
rect 9128 3587 9180 3596
rect 1860 3476 1912 3528
rect 4436 3476 4488 3528
rect 6644 3408 6696 3460
rect 7472 3476 7524 3528
rect 7564 3476 7616 3528
rect 7380 3408 7432 3460
rect 8116 3476 8168 3528
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9128 3544 9180 3553
rect 9220 3544 9272 3596
rect 12440 3544 12492 3596
rect 8576 3476 8628 3528
rect 8668 3408 8720 3460
rect 10140 3476 10192 3528
rect 10876 3476 10928 3528
rect 13452 3544 13504 3596
rect 14280 3723 14332 3732
rect 14280 3689 14289 3723
rect 14289 3689 14323 3723
rect 14323 3689 14332 3723
rect 14280 3680 14332 3689
rect 14096 3655 14148 3664
rect 14096 3621 14105 3655
rect 14105 3621 14139 3655
rect 14139 3621 14148 3655
rect 14096 3612 14148 3621
rect 15660 3544 15712 3596
rect 12992 3519 13044 3528
rect 11060 3408 11112 3460
rect 11428 3451 11480 3460
rect 11428 3417 11437 3451
rect 11437 3417 11471 3451
rect 11471 3417 11480 3451
rect 11428 3408 11480 3417
rect 11796 3408 11848 3460
rect 7656 3340 7708 3392
rect 8760 3340 8812 3392
rect 9220 3340 9272 3392
rect 10140 3340 10192 3392
rect 11244 3340 11296 3392
rect 11520 3383 11572 3392
rect 11520 3349 11529 3383
rect 11529 3349 11563 3383
rect 11563 3349 11572 3383
rect 11520 3340 11572 3349
rect 12348 3340 12400 3392
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 14188 3476 14240 3528
rect 12716 3340 12768 3392
rect 14740 3340 14792 3392
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 3148 3179 3200 3188
rect 3148 3145 3157 3179
rect 3157 3145 3191 3179
rect 3191 3145 3200 3179
rect 3148 3136 3200 3145
rect 3792 3179 3844 3188
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 8576 3136 8628 3188
rect 8852 3179 8904 3188
rect 8852 3145 8861 3179
rect 8861 3145 8895 3179
rect 8895 3145 8904 3179
rect 8852 3136 8904 3145
rect 9128 3136 9180 3188
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 10968 3136 11020 3188
rect 4436 3068 4488 3120
rect 8760 3068 8812 3120
rect 3516 3000 3568 3052
rect 6000 3000 6052 3052
rect 9220 3068 9272 3120
rect 11796 3136 11848 3188
rect 12440 3136 12492 3188
rect 11152 3068 11204 3120
rect 13268 3068 13320 3120
rect 13728 3068 13780 3120
rect 9864 3000 9916 3052
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10140 3000 10192 3009
rect 10508 3000 10560 3052
rect 11704 3000 11756 3052
rect 10048 2932 10100 2984
rect 10784 2932 10836 2984
rect 12348 2932 12400 2984
rect 14556 2932 14608 2984
rect 8300 2864 8352 2916
rect 8760 2864 8812 2916
rect 3792 2796 3844 2848
rect 10232 2796 10284 2848
rect 13360 2796 13412 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 6276 2592 6328 2644
rect 4068 2524 4120 2576
rect 9036 2592 9088 2644
rect 1676 2456 1728 2508
rect 5816 2456 5868 2508
rect 9680 2524 9732 2576
rect 11520 2567 11572 2576
rect 11520 2533 11529 2567
rect 11529 2533 11563 2567
rect 11563 2533 11572 2567
rect 11520 2524 11572 2533
rect 11796 2524 11848 2576
rect 13360 2524 13412 2576
rect 9956 2456 10008 2508
rect 13268 2499 13320 2508
rect 13268 2465 13277 2499
rect 13277 2465 13311 2499
rect 13311 2465 13320 2499
rect 13268 2456 13320 2465
rect 4160 2388 4212 2440
rect 8024 2388 8076 2440
rect 8116 2388 8168 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 2504 2320 2556 2372
rect 7380 2320 7432 2372
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 13636 2592 13688 2644
rect 11704 2388 11756 2397
rect 13544 2388 13596 2440
rect 9588 2295 9640 2304
rect 9588 2261 9597 2295
rect 9597 2261 9631 2295
rect 9631 2261 9640 2295
rect 9588 2252 9640 2261
rect 10140 2295 10192 2304
rect 10140 2261 10149 2295
rect 10149 2261 10183 2295
rect 10183 2261 10192 2295
rect 10140 2252 10192 2261
rect 10876 2363 10928 2372
rect 10876 2329 10885 2363
rect 10885 2329 10919 2363
rect 10919 2329 10928 2363
rect 10876 2320 10928 2329
rect 10968 2363 11020 2372
rect 10968 2329 10977 2363
rect 10977 2329 11011 2363
rect 11011 2329 11020 2363
rect 10968 2320 11020 2329
rect 11244 2295 11296 2304
rect 11244 2261 11253 2295
rect 11253 2261 11287 2295
rect 11287 2261 11296 2295
rect 11244 2252 11296 2261
rect 12532 2295 12584 2304
rect 12532 2261 12541 2295
rect 12541 2261 12575 2295
rect 12575 2261 12584 2295
rect 12532 2252 12584 2261
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 13912 2295 13964 2304
rect 13912 2261 13921 2295
rect 13921 2261 13955 2295
rect 13955 2261 13964 2295
rect 13912 2252 13964 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 1216 2048 1268 2100
rect 12532 2048 12584 2100
rect 8024 1980 8076 2032
rect 9128 1980 9180 2032
rect 10140 1980 10192 2032
rect 13176 1980 13228 2032
rect 4712 1844 4764 1896
rect 9588 1844 9640 1896
rect 6736 1640 6788 1692
rect 11244 1640 11296 1692
<< metal2 >>
rect 14462 16416 14518 16425
rect 14462 16351 14518 16360
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 664 15904 716 15910
rect 664 15846 716 15852
rect 676 7410 704 15846
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 2318 15600 2374 15609
rect 2318 15535 2374 15544
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1872 14822 1900 14962
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 940 14544 992 14550
rect 940 14486 992 14492
rect 754 10024 810 10033
rect 754 9959 810 9968
rect 664 7404 716 7410
rect 664 7346 716 7352
rect 768 6934 796 9959
rect 848 9580 900 9586
rect 848 9522 900 9528
rect 860 7546 888 9522
rect 848 7540 900 7546
rect 848 7482 900 7488
rect 848 7404 900 7410
rect 848 7346 900 7352
rect 756 6928 808 6934
rect 756 6870 808 6876
rect 860 4554 888 7346
rect 848 4548 900 4554
rect 848 4490 900 4496
rect 952 4185 980 14486
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13433 1440 13874
rect 1398 13424 1454 13433
rect 1398 13359 1454 13368
rect 1124 13252 1176 13258
rect 1124 13194 1176 13200
rect 1030 12336 1086 12345
rect 1030 12271 1086 12280
rect 1044 4758 1072 12271
rect 1032 4752 1084 4758
rect 1032 4694 1084 4700
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1136 3505 1164 13194
rect 1308 13184 1360 13190
rect 1308 13126 1360 13132
rect 1216 12776 1268 12782
rect 1216 12718 1268 12724
rect 1122 3496 1178 3505
rect 1122 3431 1178 3440
rect 1228 2106 1256 12718
rect 1320 9625 1348 13126
rect 1504 11354 1532 14758
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1596 14521 1624 14554
rect 1582 14512 1638 14521
rect 1582 14447 1638 14456
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1780 13977 1808 14214
rect 1766 13968 1822 13977
rect 1766 13903 1822 13912
rect 1768 13864 1820 13870
rect 1766 13832 1768 13841
rect 1820 13832 1822 13841
rect 1766 13767 1822 13776
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1398 11248 1454 11257
rect 1398 11183 1454 11192
rect 1306 9616 1362 9625
rect 1306 9551 1362 9560
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 1320 4826 1348 9454
rect 1308 4820 1360 4826
rect 1308 4762 1360 4768
rect 1412 3738 1440 11183
rect 1504 9586 1532 11290
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1504 5710 1532 9386
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1596 4010 1624 11086
rect 1688 10713 1716 13670
rect 1766 11792 1822 11801
rect 1766 11727 1822 11736
rect 1674 10704 1730 10713
rect 1674 10639 1730 10648
rect 1676 10532 1728 10538
rect 1676 10474 1728 10480
rect 1584 4004 1636 4010
rect 1584 3946 1636 3952
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 1688 2514 1716 10474
rect 1780 7478 1808 11727
rect 1872 8401 1900 14282
rect 1964 13938 1992 14418
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2240 13818 2268 13874
rect 2148 13790 2268 13818
rect 2148 13734 2176 13790
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2240 9518 2268 10202
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 1858 8392 1914 8401
rect 1858 8327 1914 8336
rect 2240 8294 2268 9114
rect 2332 8566 2360 15535
rect 4896 15496 4948 15502
rect 3606 15464 3662 15473
rect 4896 15438 4948 15444
rect 3606 15399 3662 15408
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 2424 15162 2452 15302
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 3252 14958 3280 15302
rect 3240 14952 3292 14958
rect 3292 14900 3464 14906
rect 3240 14894 3464 14900
rect 3148 14884 3200 14890
rect 3252 14878 3464 14894
rect 3148 14826 3200 14832
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 2780 14000 2832 14006
rect 2976 13954 3004 14214
rect 2832 13948 3004 13954
rect 2780 13942 3004 13948
rect 2792 13926 3004 13942
rect 2884 13326 2912 13926
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2424 10810 2452 12854
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2410 10704 2466 10713
rect 2410 10639 2466 10648
rect 2424 10441 2452 10639
rect 2410 10432 2466 10441
rect 2410 10367 2466 10376
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 2228 8288 2280 8294
rect 2424 8242 2452 10367
rect 2228 8230 2280 8236
rect 1872 7886 1900 8230
rect 2332 8214 2452 8242
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2332 7886 2360 8214
rect 2410 8120 2466 8129
rect 2410 8055 2466 8064
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 1768 7472 1820 7478
rect 1766 7440 1768 7449
rect 1820 7440 1822 7449
rect 2240 7410 2268 7822
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 1766 7375 1822 7384
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2332 7313 2360 7686
rect 1858 7304 1914 7313
rect 1858 7239 1914 7248
rect 2318 7304 2374 7313
rect 2318 7239 2374 7248
rect 1872 4622 1900 7239
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1780 4486 1808 4558
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1872 3534 1900 4558
rect 2332 3890 2360 7142
rect 2424 4690 2452 8055
rect 2516 7342 2544 12786
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2778 11792 2834 11801
rect 2778 11727 2780 11736
rect 2832 11727 2834 11736
rect 2780 11698 2832 11704
rect 2594 11384 2650 11393
rect 2792 11354 2820 11698
rect 2976 11558 3004 11834
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2594 11319 2596 11328
rect 2648 11319 2650 11328
rect 2780 11348 2832 11354
rect 2596 11290 2648 11296
rect 2780 11290 2832 11296
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2792 10470 2820 10610
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 9926 2820 10406
rect 2976 10266 3004 11494
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2962 10160 3018 10169
rect 2962 10095 3018 10104
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 8838 2636 9454
rect 2792 9178 2820 9522
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 9217 2912 9386
rect 2870 9208 2926 9217
rect 2780 9172 2832 9178
rect 2870 9143 2926 9152
rect 2780 9114 2832 9120
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2976 7546 3004 10095
rect 3068 9654 3096 12922
rect 3160 12782 3188 14826
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3160 11218 3188 12718
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 9994 3188 10610
rect 3252 10418 3280 14758
rect 3330 13424 3386 13433
rect 3330 13359 3386 13368
rect 3344 10810 3372 13359
rect 3436 12832 3464 14878
rect 3620 14006 3648 15399
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3528 13394 3556 13806
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3528 13002 3556 13330
rect 3608 13320 3660 13326
rect 3606 13288 3608 13297
rect 3660 13288 3662 13297
rect 3606 13223 3662 13232
rect 3528 12986 3648 13002
rect 3516 12980 3648 12986
rect 3568 12974 3648 12980
rect 3516 12922 3568 12928
rect 3436 12804 3556 12832
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3436 11762 3464 12378
rect 3528 11801 3556 12804
rect 3620 12102 3648 12974
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3514 11792 3570 11801
rect 3424 11756 3476 11762
rect 3514 11727 3570 11736
rect 3608 11756 3660 11762
rect 3424 11698 3476 11704
rect 3608 11698 3660 11704
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3620 11506 3648 11698
rect 3804 11665 3832 14418
rect 3790 11656 3846 11665
rect 3790 11591 3846 11600
rect 3436 11121 3464 11494
rect 3422 11112 3478 11121
rect 3422 11047 3478 11056
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3424 10464 3476 10470
rect 3252 10412 3424 10418
rect 3252 10406 3476 10412
rect 3252 10390 3464 10406
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 8809 3096 9318
rect 3148 8832 3200 8838
rect 3054 8800 3110 8809
rect 3148 8774 3200 8780
rect 3054 8735 3110 8744
rect 3056 8424 3108 8430
rect 3054 8392 3056 8401
rect 3108 8392 3110 8401
rect 3054 8327 3110 8336
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2608 7188 2636 7482
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2516 7160 2636 7188
rect 2516 4758 2544 7160
rect 2700 6914 2728 7278
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2700 6886 2820 6914
rect 2792 6769 2820 6886
rect 2976 6798 3004 6938
rect 3054 6896 3110 6905
rect 3054 6831 3056 6840
rect 3108 6831 3110 6840
rect 3056 6802 3108 6808
rect 2964 6792 3016 6798
rect 2778 6760 2834 6769
rect 2964 6734 3016 6740
rect 2778 6695 2834 6704
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 3160 6066 3188 8774
rect 3068 6038 3188 6066
rect 2962 5808 3018 5817
rect 2962 5743 3018 5752
rect 2976 5710 3004 5743
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2516 4162 2544 4422
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2976 4282 3004 4490
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2596 4208 2648 4214
rect 2516 4156 2596 4162
rect 2516 4150 2648 4156
rect 2516 4134 2636 4150
rect 2410 3904 2466 3913
rect 2332 3862 2410 3890
rect 1950 3836 2258 3845
rect 2410 3839 2466 3848
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2608 3738 2636 4134
rect 3068 4078 3096 6038
rect 3146 5944 3202 5953
rect 3252 5914 3280 10202
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 3344 9586 3372 10134
rect 3436 9586 3464 10390
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 8265 3372 9318
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3330 8256 3386 8265
rect 3330 8191 3386 8200
rect 3436 8106 3464 9114
rect 3344 8078 3464 8106
rect 3344 6610 3372 8078
rect 3422 7984 3478 7993
rect 3422 7919 3478 7928
rect 3436 7478 3464 7919
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3344 6582 3464 6610
rect 3330 6488 3386 6497
rect 3330 6423 3386 6432
rect 3146 5879 3202 5888
rect 3240 5908 3292 5914
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 3160 3194 3188 5879
rect 3240 5850 3292 5856
rect 3344 5778 3372 6423
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3238 5672 3294 5681
rect 3238 5607 3294 5616
rect 3252 5370 3280 5607
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3252 4758 3280 5306
rect 3436 5302 3464 6582
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4282 3280 4558
rect 3344 4486 3372 5170
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3528 3058 3556 11494
rect 3620 11478 3832 11506
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3620 11121 3648 11290
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3606 11112 3662 11121
rect 3606 11047 3662 11056
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3620 6798 3648 9522
rect 3712 7886 3740 11154
rect 3804 8673 3832 11478
rect 3896 11098 3924 15098
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 4252 14952 4304 14958
rect 4250 14920 4252 14929
rect 4304 14920 4306 14929
rect 4250 14855 4306 14864
rect 4356 14550 4384 15030
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4160 14408 4212 14414
rect 4540 14362 4568 14894
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4160 14350 4212 14356
rect 4172 14074 4200 14350
rect 4356 14334 4568 14362
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4356 13938 4384 14334
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13161 4016 13670
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 3974 13152 4030 13161
rect 3974 13087 4030 13096
rect 4080 11626 4108 13466
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12782 4292 13126
rect 4356 13025 4384 13194
rect 4342 13016 4398 13025
rect 4342 12951 4398 12960
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4342 12472 4398 12481
rect 4342 12407 4398 12416
rect 4356 12306 4384 12407
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3974 11384 4030 11393
rect 3974 11319 4030 11328
rect 3988 11286 4016 11319
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3896 11070 4016 11098
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3790 8664 3846 8673
rect 3790 8599 3846 8608
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3712 7206 3740 7686
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3606 6624 3662 6633
rect 3606 6559 3662 6568
rect 3620 6458 3648 6559
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3620 5710 3648 6394
rect 3804 5846 3832 8366
rect 3896 6798 3924 10066
rect 3988 9178 4016 11070
rect 4080 9518 4108 11562
rect 4264 11150 4292 11698
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10266 4200 11018
rect 4264 10985 4292 11086
rect 4250 10976 4306 10985
rect 4250 10911 4306 10920
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9586 4200 9998
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4158 9480 4214 9489
rect 4158 9415 4214 9424
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3974 8256 4030 8265
rect 3974 8191 4030 8200
rect 3988 7886 4016 8191
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6390 3924 6598
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3882 6216 3938 6225
rect 3882 6151 3938 6160
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3620 5370 3648 5510
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3620 3641 3648 5306
rect 3712 5137 3740 5782
rect 3896 5642 3924 6151
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3988 5545 4016 7686
rect 4080 7546 4108 9318
rect 4172 8974 4200 9415
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4158 8392 4214 8401
rect 4158 8327 4214 8336
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4172 7342 4200 8327
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4172 6458 4200 7278
rect 4264 6798 4292 9658
rect 4356 7546 4384 11222
rect 4448 10674 4476 14214
rect 4632 14006 4660 14214
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4724 13938 4752 14554
rect 4804 14000 4856 14006
rect 4802 13968 4804 13977
rect 4856 13968 4858 13977
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4712 13932 4764 13938
rect 4802 13903 4858 13912
rect 4712 13874 4764 13880
rect 4540 13841 4568 13874
rect 4526 13832 4582 13841
rect 4526 13767 4582 13776
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4632 13530 4660 13670
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4526 13016 4582 13025
rect 4526 12951 4582 12960
rect 4540 12442 4568 12951
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4448 9722 4476 10610
rect 4540 10198 4568 12242
rect 4632 11014 4660 13466
rect 4712 13184 4764 13190
rect 4710 13152 4712 13161
rect 4764 13152 4766 13161
rect 4710 13087 4766 13096
rect 4908 12714 4936 15438
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 5092 14249 5120 15302
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 5078 14240 5134 14249
rect 5078 14175 5134 14184
rect 4986 12744 5042 12753
rect 4896 12708 4948 12714
rect 4986 12679 5042 12688
rect 4896 12650 4948 12656
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12170 4752 12582
rect 4908 12434 4936 12650
rect 4816 12406 4936 12434
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4712 11824 4764 11830
rect 4710 11792 4712 11801
rect 4764 11792 4766 11801
rect 4710 11727 4766 11736
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4724 10810 4752 11630
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4724 10441 4752 10542
rect 4710 10432 4766 10441
rect 4710 10367 4766 10376
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4526 9752 4582 9761
rect 4436 9716 4488 9722
rect 4526 9687 4582 9696
rect 4436 9658 4488 9664
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4448 9353 4476 9386
rect 4434 9344 4490 9353
rect 4434 9279 4490 9288
rect 4436 9104 4488 9110
rect 4434 9072 4436 9081
rect 4488 9072 4490 9081
rect 4434 9007 4490 9016
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8294 4476 8774
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4448 7886 4476 8230
rect 4540 8090 4568 9687
rect 4816 9674 4844 12406
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4908 11218 4936 11766
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10606 4936 10950
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4632 9646 4844 9674
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4448 7721 4476 7822
rect 4434 7712 4490 7721
rect 4434 7647 4490 7656
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4252 6792 4304 6798
rect 4540 6746 4568 7822
rect 4632 7342 4660 9646
rect 4908 9602 4936 10542
rect 4724 9574 4936 9602
rect 4724 8838 4752 9574
rect 4802 9344 4858 9353
rect 4802 9279 4858 9288
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4724 7818 4752 8774
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4252 6734 4304 6740
rect 4356 6718 4568 6746
rect 4356 6662 4384 6718
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5914 4108 6122
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4172 5817 4200 5850
rect 4158 5808 4214 5817
rect 4158 5743 4214 5752
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3974 5536 4030 5545
rect 3974 5471 4030 5480
rect 3790 5264 3846 5273
rect 3790 5199 3846 5208
rect 3698 5128 3754 5137
rect 3698 5063 3754 5072
rect 3606 3632 3662 3641
rect 3606 3567 3662 3576
rect 3804 3194 3832 5199
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3804 2854 3832 3130
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 4080 2582 4108 5646
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5370 4200 5510
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4264 5234 4292 6258
rect 4252 5228 4304 5234
rect 4252 5170 4304 5176
rect 4356 5098 4384 6598
rect 4448 6361 4476 6598
rect 4434 6352 4490 6361
rect 4434 6287 4490 6296
rect 4540 6254 4568 6598
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5778 4568 6054
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4448 5574 4476 5646
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4068 2576 4120 2582
rect 4068 2518 4120 2524
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 4172 2446 4200 4422
rect 4448 3534 4476 5510
rect 4540 5273 4568 5578
rect 4632 5370 4660 7278
rect 4724 6662 4752 7754
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4526 5264 4582 5273
rect 4526 5199 4582 5208
rect 4540 5166 4568 5199
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4632 3670 4660 5306
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4448 3126 4476 3470
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 1216 2100 1268 2106
rect 1216 2042 1268 2048
rect 2516 2009 2544 2314
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 2502 2000 2558 2009
rect 2502 1935 2558 1944
rect 4724 1902 4752 6258
rect 4816 3738 4844 9279
rect 5000 8906 5028 12679
rect 5092 10690 5120 14175
rect 5184 11830 5212 14826
rect 5368 14822 5396 14962
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5276 14278 5304 14554
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5368 13870 5396 14758
rect 5356 13864 5408 13870
rect 5644 13841 5672 14758
rect 5736 14482 5764 14826
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5356 13806 5408 13812
rect 5630 13832 5686 13841
rect 5368 13734 5396 13806
rect 5630 13767 5686 13776
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5460 13326 5488 13670
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5184 10985 5212 11290
rect 5170 10976 5226 10985
rect 5170 10911 5226 10920
rect 5276 10810 5304 13194
rect 5368 12345 5396 13194
rect 5552 13172 5580 13398
rect 5460 13144 5580 13172
rect 5460 12442 5488 13144
rect 5736 12850 5764 13874
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5538 12608 5594 12617
rect 5538 12543 5594 12552
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5354 12336 5410 12345
rect 5354 12271 5410 12280
rect 5460 11762 5488 12378
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5552 11694 5580 12543
rect 5736 12356 5764 12786
rect 5736 12328 5856 12356
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5644 11830 5672 12242
rect 5632 11824 5684 11830
rect 5632 11766 5684 11772
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5354 11248 5410 11257
rect 5354 11183 5356 11192
rect 5408 11183 5410 11192
rect 5356 11154 5408 11160
rect 5538 10976 5594 10985
rect 5538 10911 5594 10920
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5092 10662 5212 10690
rect 5078 10432 5134 10441
rect 5078 10367 5134 10376
rect 5092 9382 5120 10367
rect 5184 9674 5212 10662
rect 5276 10062 5304 10746
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5368 10198 5396 10542
rect 5460 10470 5488 10542
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5552 10130 5580 10911
rect 5644 10266 5672 11766
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11393 5764 11494
rect 5722 11384 5778 11393
rect 5722 11319 5778 11328
rect 5828 11268 5856 12328
rect 5736 11240 5856 11268
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5540 9920 5592 9926
rect 5446 9888 5502 9897
rect 5540 9862 5592 9868
rect 5446 9823 5502 9832
rect 5356 9716 5408 9722
rect 5184 9646 5304 9674
rect 5356 9658 5408 9664
rect 5080 9376 5132 9382
rect 5276 9364 5304 9646
rect 5080 9318 5132 9324
rect 5184 9336 5304 9364
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4986 8664 5042 8673
rect 4986 8599 5042 8608
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4908 7002 4936 8230
rect 5000 7993 5028 8599
rect 5184 8430 5212 9336
rect 5368 9178 5396 9658
rect 5460 9602 5488 9823
rect 5451 9574 5488 9602
rect 5451 9518 5479 9574
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5446 8664 5502 8673
rect 5552 8634 5580 9862
rect 5644 9722 5672 10202
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5736 9330 5764 11240
rect 5920 10742 5948 14962
rect 6012 13802 6040 15370
rect 6656 15162 6684 15914
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 15178 6868 15302
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6644 15156 6696 15162
rect 6840 15150 7328 15178
rect 6644 15098 6696 15104
rect 6564 14414 6592 15098
rect 6932 15094 6960 15150
rect 7300 15094 7328 15150
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14822 7144 14962
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6092 14272 6144 14278
rect 6090 14240 6092 14249
rect 6144 14240 6146 14249
rect 6090 14175 6146 14184
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6182 13968 6238 13977
rect 6182 13903 6238 13912
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 6196 12986 6224 13903
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6012 12714 6040 12786
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6196 12209 6224 12786
rect 6182 12200 6238 12209
rect 6092 12164 6144 12170
rect 6182 12135 6238 12144
rect 6092 12106 6144 12112
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5644 9302 5764 9330
rect 5644 8888 5672 9302
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5736 9042 5764 9114
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5724 8900 5776 8906
rect 5644 8860 5724 8888
rect 5724 8842 5776 8848
rect 5630 8664 5686 8673
rect 5446 8599 5502 8608
rect 5540 8628 5592 8634
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5460 8362 5488 8599
rect 5630 8599 5686 8608
rect 5540 8570 5592 8576
rect 5644 8430 5672 8599
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4986 7984 5042 7993
rect 4986 7919 5042 7928
rect 5092 7886 5120 8026
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4986 7576 5042 7585
rect 4986 7511 5042 7520
rect 5000 7002 5028 7511
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4986 6896 5042 6905
rect 4986 6831 5042 6840
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4908 3097 4936 6734
rect 5000 5642 5028 6831
rect 5092 5914 5120 7822
rect 5184 6202 5212 7890
rect 5276 6322 5304 8298
rect 5356 7880 5408 7886
rect 5408 7840 5488 7868
rect 5356 7822 5408 7828
rect 5460 7750 5488 7840
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5184 6174 5304 6202
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 5000 4486 5028 5306
rect 5184 5302 5212 5578
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5000 4282 5028 4422
rect 5184 4282 5212 5238
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5276 3602 5304 6174
rect 5368 6100 5396 7686
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5460 6866 5488 7482
rect 5552 7274 5580 8366
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5540 6928 5592 6934
rect 5644 6914 5672 8366
rect 5736 8294 5764 8842
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5592 6886 5672 6914
rect 5540 6870 5592 6876
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6202 5488 6598
rect 5552 6440 5580 6870
rect 5736 6798 5764 7890
rect 5724 6792 5776 6798
rect 5630 6760 5686 6769
rect 5724 6734 5776 6740
rect 5630 6695 5686 6704
rect 5644 6662 5672 6695
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5632 6452 5684 6458
rect 5552 6412 5632 6440
rect 5632 6394 5684 6400
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5460 6174 5580 6202
rect 5448 6112 5500 6118
rect 5368 6072 5448 6100
rect 5368 5370 5396 6072
rect 5448 6054 5500 6060
rect 5446 5672 5502 5681
rect 5446 5607 5448 5616
rect 5500 5607 5502 5616
rect 5448 5578 5500 5584
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5552 5080 5580 6174
rect 5644 5914 5672 6258
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5644 5778 5672 5850
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5460 5052 5580 5080
rect 5356 4752 5408 4758
rect 5354 4720 5356 4729
rect 5408 4720 5410 4729
rect 5354 4655 5410 4664
rect 5460 4554 5488 5052
rect 5644 5012 5672 5714
rect 5736 5302 5764 6326
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5552 4984 5672 5012
rect 5552 4690 5580 4984
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5644 4622 5672 4762
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5736 4010 5764 5238
rect 5828 5098 5856 10610
rect 5920 9926 5948 10678
rect 6104 10305 6132 12106
rect 6288 11880 6316 12854
rect 6472 12850 6500 13466
rect 6748 13190 6776 13806
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6196 11852 6316 11880
rect 6366 11928 6422 11937
rect 6366 11863 6422 11872
rect 6196 11257 6224 11852
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 6182 11248 6238 11257
rect 6182 11183 6238 11192
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6090 10296 6146 10305
rect 6090 10231 6146 10240
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 6104 9722 6132 10134
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6196 9654 6224 10950
rect 6288 10606 6316 11698
rect 6380 10810 6408 11863
rect 6472 11370 6500 12786
rect 6748 12714 6776 12786
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6552 12232 6604 12238
rect 6656 12209 6684 12650
rect 6748 12617 6776 12650
rect 6734 12608 6790 12617
rect 6734 12543 6790 12552
rect 6734 12472 6790 12481
rect 6734 12407 6790 12416
rect 6840 12424 6868 14010
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 7288 13320 7340 13326
rect 7194 13288 7250 13297
rect 7288 13262 7340 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7194 13223 7250 13232
rect 7208 12730 7236 13223
rect 7300 13161 7328 13262
rect 7286 13152 7342 13161
rect 7286 13087 7342 13096
rect 7208 12702 7328 12730
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 6748 12306 6776 12407
rect 6840 12396 7052 12424
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6552 12174 6604 12180
rect 6642 12200 6698 12209
rect 6564 11558 6592 12174
rect 6642 12135 6698 12144
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11937 6960 12106
rect 6918 11928 6974 11937
rect 6918 11863 6974 11872
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6656 11370 6684 11698
rect 7024 11540 7052 12396
rect 7102 12064 7158 12073
rect 7102 11999 7158 12008
rect 7116 11762 7144 11999
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 6472 11342 6684 11370
rect 6840 11512 7052 11540
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6366 10704 6422 10713
rect 6366 10639 6368 10648
rect 6420 10639 6422 10648
rect 6368 10610 6420 10616
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6288 10169 6316 10542
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6274 10160 6330 10169
rect 6274 10095 6330 10104
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6288 9586 6316 9998
rect 6380 9654 6408 10406
rect 6472 10169 6500 11018
rect 6458 10160 6514 10169
rect 6458 10095 6514 10104
rect 6564 9994 6592 11342
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10810 6684 10950
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6642 10704 6698 10713
rect 6840 10674 6868 11512
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6918 11248 6974 11257
rect 7024 11218 7052 11290
rect 7102 11248 7158 11257
rect 6918 11183 6974 11192
rect 7012 11212 7064 11218
rect 6932 10742 6960 11183
rect 7102 11183 7158 11192
rect 7196 11212 7248 11218
rect 7012 11154 7064 11160
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10849 7052 11018
rect 7116 11014 7144 11183
rect 7196 11154 7248 11160
rect 7104 11008 7156 11014
rect 7208 10985 7236 11154
rect 7300 11150 7328 12702
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7288 11008 7340 11014
rect 7104 10950 7156 10956
rect 7194 10976 7250 10985
rect 7288 10950 7340 10956
rect 7194 10911 7250 10920
rect 7010 10840 7066 10849
rect 7300 10810 7328 10950
rect 7392 10849 7420 13262
rect 7484 13025 7512 14554
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 8128 14113 8156 15098
rect 8114 14104 8170 14113
rect 8114 14039 8170 14048
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7576 13326 7604 13670
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7470 13016 7526 13025
rect 7610 13019 7918 13028
rect 8036 12968 8064 13738
rect 8220 13462 8248 15506
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8312 13870 8340 14486
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 7470 12951 7526 12960
rect 7484 11257 7512 12951
rect 7760 12940 8064 12968
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 12481 7604 12650
rect 7562 12472 7618 12481
rect 7562 12407 7618 12416
rect 7760 12170 7788 12940
rect 8128 12434 8156 13398
rect 8312 13258 8340 13670
rect 8300 13252 8352 13258
rect 8220 13212 8300 13240
rect 8220 12646 8248 13212
rect 8300 13194 8352 13200
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 8312 12434 8340 12854
rect 8404 12442 8432 14758
rect 8496 14074 8524 14894
rect 8956 14414 8984 15438
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8772 14249 8800 14350
rect 8758 14240 8814 14249
rect 8758 14175 8814 14184
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8496 13161 8524 13398
rect 8956 13394 8984 14350
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 9048 13530 9076 13942
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 8482 13152 8538 13161
rect 8482 13087 8538 13096
rect 8482 12744 8538 12753
rect 8482 12679 8538 12688
rect 8036 12406 8156 12434
rect 8220 12406 8340 12434
rect 8392 12436 8444 12442
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7654 11520 7710 11529
rect 7654 11455 7710 11464
rect 7668 11286 7696 11455
rect 7656 11280 7708 11286
rect 7470 11248 7526 11257
rect 7760 11257 7788 11630
rect 7840 11280 7892 11286
rect 7656 11222 7708 11228
rect 7746 11248 7802 11257
rect 7470 11183 7526 11192
rect 7840 11222 7892 11228
rect 7746 11183 7802 11192
rect 7378 10840 7434 10849
rect 7010 10775 7066 10784
rect 7288 10804 7340 10810
rect 7484 10826 7512 11183
rect 7852 11082 7880 11222
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 8036 10826 8064 12406
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 7484 10798 7521 10826
rect 7378 10775 7434 10784
rect 7493 10792 7521 10798
rect 7564 10804 7616 10810
rect 7493 10764 7564 10792
rect 7288 10746 7340 10752
rect 7564 10746 7616 10752
rect 7944 10798 8064 10826
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 7392 10674 7788 10690
rect 6642 10639 6698 10648
rect 6828 10668 6880 10674
rect 6656 10033 6684 10639
rect 6828 10610 6880 10616
rect 7392 10668 7800 10674
rect 7392 10662 7748 10668
rect 6736 10600 6788 10606
rect 7392 10554 7420 10662
rect 7748 10610 7800 10616
rect 6788 10548 7420 10554
rect 6736 10542 7420 10548
rect 6748 10526 7420 10542
rect 6736 10464 6788 10470
rect 6734 10432 6736 10441
rect 6788 10432 6790 10441
rect 6734 10367 6790 10376
rect 7378 10432 7434 10441
rect 7944 10418 7972 10798
rect 6950 10364 7258 10373
rect 7378 10367 7434 10376
rect 7484 10390 7972 10418
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6734 10296 6790 10305
rect 6950 10299 7258 10308
rect 6920 10260 6972 10266
rect 6790 10240 6920 10248
rect 6734 10231 6920 10240
rect 6748 10220 6920 10231
rect 6920 10202 6972 10208
rect 6642 10024 6698 10033
rect 6552 9988 6604 9994
rect 6642 9959 6698 9968
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6552 9930 6604 9936
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5920 9042 5948 9454
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 6012 8634 6040 9522
rect 6472 9518 6500 9658
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6184 9376 6236 9382
rect 6090 9344 6146 9353
rect 6184 9318 6236 9324
rect 6366 9344 6422 9353
rect 6090 9279 6146 9288
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5920 8294 5948 8570
rect 6012 8498 6040 8570
rect 6104 8566 6132 9279
rect 6196 8945 6224 9318
rect 6366 9279 6422 9288
rect 6182 8936 6238 8945
rect 6182 8871 6238 8880
rect 6276 8900 6328 8906
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5920 8266 6132 8294
rect 5906 7984 5962 7993
rect 6104 7954 6132 8266
rect 5906 7919 5962 7928
rect 6092 7948 6144 7954
rect 5920 7478 5948 7919
rect 6092 7890 6144 7896
rect 6196 7886 6224 8871
rect 6276 8842 6328 8848
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5906 7304 5962 7313
rect 5906 7239 5962 7248
rect 5920 6390 5948 7239
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5920 6118 5948 6190
rect 6012 6118 6040 7754
rect 6184 7744 6236 7750
rect 6182 7712 6184 7721
rect 6236 7712 6238 7721
rect 6182 7647 6238 7656
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6104 6934 6132 7210
rect 6092 6928 6144 6934
rect 6196 6916 6224 7647
rect 6288 7041 6316 8842
rect 6380 7392 6408 9279
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6472 7546 6500 7754
rect 6564 7546 6592 9930
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6748 9722 6776 9862
rect 6736 9716 6788 9722
rect 6656 9676 6736 9704
rect 6656 8022 6684 9676
rect 6736 9658 6788 9664
rect 6840 9602 6868 9862
rect 6748 9574 6868 9602
rect 6748 9353 6776 9574
rect 6932 9364 6960 9959
rect 7392 9636 7420 10367
rect 7484 9704 7512 10390
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 8036 9722 8064 10066
rect 8024 9716 8076 9722
rect 7484 9676 7604 9704
rect 7392 9608 7491 9636
rect 7463 9602 7491 9608
rect 7463 9574 7512 9602
rect 7484 9500 7512 9574
rect 7392 9472 7512 9500
rect 6734 9344 6790 9353
rect 6734 9279 6790 9288
rect 6840 9336 6960 9364
rect 7288 9376 7340 9382
rect 6734 9208 6790 9217
rect 6734 9143 6790 9152
rect 6748 8498 6776 9143
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6840 8294 6868 9336
rect 7288 9318 7340 9324
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 7300 9110 7328 9318
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 6920 8968 6972 8974
rect 6918 8936 6920 8945
rect 6972 8936 6974 8945
rect 6918 8871 6974 8880
rect 6840 8248 6960 8294
rect 7196 8288 7248 8294
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6460 7404 6512 7410
rect 6380 7364 6460 7392
rect 6274 7032 6330 7041
rect 6274 6967 6330 6976
rect 6196 6888 6316 6916
rect 6092 6870 6144 6876
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6196 5914 6224 6734
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5920 5030 5948 5714
rect 5998 5536 6054 5545
rect 5998 5471 6054 5480
rect 6012 5030 6040 5471
rect 6196 5370 6224 5850
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6182 5264 6238 5273
rect 6182 5199 6238 5208
rect 6196 5098 6224 5199
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 4894 3088 4950 3097
rect 4894 3023 4950 3032
rect 5828 2514 5856 4558
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6012 3058 6040 4422
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6288 2650 6316 6888
rect 6380 6118 6408 7364
rect 6460 7346 6512 7352
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6472 6730 6500 6938
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6472 6322 6500 6666
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6380 5030 6408 6054
rect 6460 5296 6512 5302
rect 6458 5264 6460 5273
rect 6512 5264 6514 5273
rect 6458 5199 6514 5208
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6564 4554 6592 6054
rect 6656 5710 6684 7754
rect 6840 7546 6868 8248
rect 7248 8248 7328 8276
rect 7196 8230 7248 8236
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 7300 8072 7328 8248
rect 7208 8044 7328 8072
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6748 7313 6776 7482
rect 7116 7342 7144 7822
rect 7208 7410 7236 8044
rect 7392 7546 7420 9472
rect 7470 9208 7526 9217
rect 7470 9143 7526 9152
rect 7484 9042 7512 9143
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7576 8922 7604 9676
rect 8024 9658 8076 9664
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7484 8894 7604 8922
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7484 7426 7512 8894
rect 7668 8838 7696 9522
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 9042 7788 9318
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7852 8906 7880 9454
rect 8036 9382 8064 9522
rect 8128 9518 8156 12310
rect 8220 12170 8248 12406
rect 8392 12378 8444 12384
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8220 12073 8248 12106
rect 8206 12064 8262 12073
rect 8206 11999 8262 12008
rect 8312 11937 8340 12310
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 12073 8432 12174
rect 8390 12064 8446 12073
rect 8496 12050 8524 12679
rect 8588 12170 8616 13330
rect 9140 13274 9168 15438
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9232 13841 9260 14282
rect 9692 14006 9720 15846
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 14372 15632 14424 15638
rect 14186 15600 14242 15609
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 13728 15564 13780 15570
rect 14372 15574 14424 15580
rect 14186 15535 14188 15544
rect 13728 15506 13780 15512
rect 14240 15535 14242 15544
rect 14188 15506 14240 15512
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9588 14000 9640 14006
rect 9586 13968 9588 13977
rect 9680 14000 9732 14006
rect 9640 13968 9642 13977
rect 9680 13942 9732 13948
rect 9876 13938 9904 14214
rect 9586 13903 9642 13912
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9312 13864 9364 13870
rect 9218 13832 9274 13841
rect 9312 13806 9364 13812
rect 9218 13767 9274 13776
rect 8956 13246 9168 13274
rect 8758 13016 8814 13025
rect 8758 12951 8814 12960
rect 8772 12850 8800 12951
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8496 12022 8708 12050
rect 8390 11999 8446 12008
rect 8298 11928 8354 11937
rect 8298 11863 8354 11872
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8312 11558 8340 11698
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 11150 8340 11494
rect 8404 11393 8432 11834
rect 8588 11694 8616 11834
rect 8576 11688 8628 11694
rect 8574 11656 8576 11665
rect 8628 11656 8630 11665
rect 8574 11591 8630 11600
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8390 11384 8446 11393
rect 8390 11319 8446 11328
rect 8588 11218 8616 11494
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8496 10470 8524 11018
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8298 10160 8354 10169
rect 8298 10095 8354 10104
rect 8484 10124 8536 10130
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8220 9518 8248 9862
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8312 9466 8340 10095
rect 8484 10066 8536 10072
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8312 9438 8372 9466
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8344 9194 8372 9438
rect 8312 9166 8372 9194
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 8036 8650 8064 9046
rect 8208 9036 8260 9042
rect 7944 8622 8064 8650
rect 8128 8996 8208 9024
rect 7944 8514 7972 8622
rect 7852 8486 7972 8514
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 7886 7604 8298
rect 7852 7886 7880 8486
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7944 8265 7972 8366
rect 7930 8256 7986 8265
rect 7930 8191 7986 8200
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7300 7398 7512 7426
rect 7104 7336 7156 7342
rect 6734 7304 6790 7313
rect 7104 7278 7156 7284
rect 7300 7274 7328 7398
rect 7472 7336 7524 7342
rect 7472 7278 7524 7284
rect 6734 7239 6790 7248
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 6734 7168 6790 7177
rect 6734 7103 6790 7112
rect 6748 5846 6776 7103
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 7392 6848 7420 7210
rect 7116 6820 7420 6848
rect 6826 6624 6882 6633
rect 6826 6559 6882 6568
rect 6840 6458 6868 6559
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 7116 6322 7144 6820
rect 7484 6780 7512 7278
rect 8036 7018 8064 8502
rect 7208 6752 7512 6780
rect 7944 6990 8064 7018
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6840 5556 6868 6190
rect 7208 6118 7236 6752
rect 7944 6662 7972 6990
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7300 6322 7328 6598
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7470 6488 7526 6497
rect 7610 6491 7918 6500
rect 7470 6423 7526 6432
rect 7484 6390 7512 6423
rect 7472 6384 7524 6390
rect 7656 6384 7708 6390
rect 7472 6326 7524 6332
rect 7576 6344 7656 6372
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 6656 5528 6868 5556
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6564 3913 6592 3946
rect 6550 3904 6606 3913
rect 6550 3839 6606 3848
rect 6656 3466 6684 5528
rect 7196 5296 7248 5302
rect 7300 5284 7328 6258
rect 7392 6186 7420 6258
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7378 5944 7434 5953
rect 7378 5879 7434 5888
rect 7392 5574 7420 5879
rect 7576 5710 7604 6344
rect 7656 6326 7708 6332
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 6118 7880 6190
rect 8036 6118 8064 6870
rect 7840 6112 7892 6118
rect 7746 6080 7802 6089
rect 7840 6054 7892 6060
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7746 6015 7802 6024
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7760 5642 7788 6015
rect 7852 5710 7880 6054
rect 8036 5710 8064 6054
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7248 5256 7328 5284
rect 7196 5238 7248 5244
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6748 4690 6776 5102
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 6840 4690 6868 4966
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 7392 4826 7420 4966
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7484 4706 7512 5510
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 8024 5296 8076 5302
rect 7562 5264 7618 5273
rect 8024 5238 8076 5244
rect 7562 5199 7618 5208
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 7392 4678 7512 4706
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 4712 1896 4764 1902
rect 4712 1838 4764 1844
rect 6748 1698 6776 4626
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6840 2961 6868 4082
rect 7012 4072 7064 4078
rect 7010 4040 7012 4049
rect 7064 4040 7066 4049
rect 7010 3975 7066 3984
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 7392 3670 7420 4678
rect 7576 4468 7604 5199
rect 7930 4992 7986 5001
rect 7930 4927 7986 4936
rect 7944 4826 7972 4927
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7484 4440 7604 4468
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7484 3534 7512 4440
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 6826 2952 6882 2961
rect 6826 2887 6882 2896
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 7392 2378 7420 3402
rect 7576 3380 7604 3470
rect 7668 3398 7696 3674
rect 7484 3369 7604 3380
rect 7470 3360 7604 3369
rect 7526 3352 7604 3360
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7470 3295 7526 3304
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 8036 2774 8064 5238
rect 8128 3534 8156 8996
rect 8208 8978 8260 8984
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8673 8248 8774
rect 8206 8664 8262 8673
rect 8206 8599 8262 8608
rect 8220 6934 8248 8599
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8220 6730 8248 6870
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8312 6610 8340 9166
rect 8220 6582 8340 6610
rect 8220 6338 8248 6582
rect 8220 6310 8340 6338
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8220 4593 8248 6190
rect 8312 5914 8340 6310
rect 8404 6254 8432 9930
rect 8496 7206 8524 10066
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8588 9042 8616 9318
rect 8680 9042 8708 12022
rect 8864 11778 8892 12310
rect 8772 11750 8892 11778
rect 8772 11694 8800 11750
rect 8760 11688 8812 11694
rect 8852 11688 8904 11694
rect 8760 11630 8812 11636
rect 8850 11656 8852 11665
rect 8904 11656 8906 11665
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8772 8974 8800 11630
rect 8850 11591 8906 11600
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 10606 8892 11494
rect 8956 11354 8984 13246
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 11393 9076 13126
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9140 12646 9168 12786
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9232 12434 9260 12854
rect 9324 12782 9352 13806
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 13326 9444 13670
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9140 12406 9260 12434
rect 9034 11384 9090 11393
rect 8944 11348 8996 11354
rect 9034 11319 9090 11328
rect 8944 11290 8996 11296
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8956 9654 8984 11290
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8944 9376 8996 9382
rect 9048 9353 9076 10746
rect 9140 10033 9168 12406
rect 9324 12170 9352 12582
rect 9508 12434 9536 12650
rect 9600 12442 9628 12650
rect 9416 12406 9536 12434
rect 9588 12436 9640 12442
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9324 11694 9352 12106
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9324 11286 9352 11630
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9126 10024 9182 10033
rect 9126 9959 9182 9968
rect 9232 9926 9260 10610
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 8944 9318 8996 9324
rect 9034 9344 9090 9353
rect 8852 9104 8904 9110
rect 8956 9092 8984 9318
rect 9034 9279 9090 9288
rect 9140 9110 9168 9522
rect 9128 9104 9180 9110
rect 8956 9064 9100 9092
rect 8852 9046 8904 9052
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8482 7032 8538 7041
rect 8482 6967 8538 6976
rect 8496 6254 8524 6967
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8390 5808 8446 5817
rect 8390 5743 8446 5752
rect 8404 5710 8432 5743
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8206 4584 8262 4593
rect 8206 4519 8262 4528
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8312 2922 8340 5646
rect 8496 5574 8524 6190
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8390 5400 8446 5409
rect 8390 5335 8446 5344
rect 8404 5166 8432 5335
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8496 4570 8524 5510
rect 8588 5001 8616 8842
rect 8680 8498 8708 8842
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8666 8392 8722 8401
rect 8666 8327 8668 8336
rect 8720 8327 8722 8336
rect 8668 8298 8720 8304
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6089 8708 7142
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8772 6390 8800 6734
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8864 6225 8892 9046
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 6633 8984 8910
rect 9072 8888 9100 9064
rect 9128 9046 9180 9052
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9048 8860 9100 8888
rect 9048 8566 9076 8860
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 9140 8401 9168 8910
rect 9126 8392 9182 8401
rect 9126 8327 9182 8336
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 9048 8022 9076 8230
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 8942 6624 8998 6633
rect 8942 6559 8998 6568
rect 8850 6216 8906 6225
rect 8850 6151 8906 6160
rect 8666 6080 8722 6089
rect 8864 6066 8892 6151
rect 8666 6015 8722 6024
rect 8772 6038 8892 6066
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8574 4992 8630 5001
rect 8574 4927 8630 4936
rect 8680 4758 8708 5850
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8404 4078 8432 4558
rect 8496 4542 8616 4570
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8496 4214 8524 4422
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8588 3534 8616 4542
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8588 3194 8616 3470
rect 8680 3466 8708 4422
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8772 3398 8800 6038
rect 8942 5944 8998 5953
rect 8852 5908 8904 5914
rect 8942 5879 8998 5888
rect 8852 5850 8904 5856
rect 8864 5098 8892 5850
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8666 3224 8722 3233
rect 8576 3188 8628 3194
rect 8666 3159 8722 3168
rect 8576 3130 8628 3136
rect 8300 2916 8352 2922
rect 8680 2904 8708 3159
rect 8772 3126 8800 3334
rect 8864 3194 8892 4626
rect 8956 4554 8984 5879
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8956 3738 8984 4490
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8760 2916 8812 2922
rect 8680 2876 8760 2904
rect 8300 2858 8352 2864
rect 8760 2858 8812 2864
rect 8036 2746 8156 2774
rect 8128 2446 8156 2746
rect 9048 2650 9076 7958
rect 9140 7857 9168 7958
rect 9126 7848 9182 7857
rect 9126 7783 9182 7792
rect 9126 6896 9182 6905
rect 9126 6831 9128 6840
rect 9180 6831 9182 6840
rect 9128 6802 9180 6808
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9140 6497 9168 6666
rect 9126 6488 9182 6497
rect 9126 6423 9182 6432
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9140 4468 9168 5578
rect 9232 4622 9260 9862
rect 9324 9586 9352 11222
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9324 5710 9352 9386
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5234 9352 5510
rect 9416 5273 9444 12406
rect 9588 12378 9640 12384
rect 9600 11778 9628 12378
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9692 11830 9720 12242
rect 9508 11750 9628 11778
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9508 10198 9536 11750
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 9508 7002 9536 10134
rect 9600 8090 9628 11630
rect 9692 10606 9720 11766
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9217 9720 9862
rect 9784 9654 9812 13398
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9876 10742 9904 13126
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9761 9904 9862
rect 9862 9752 9918 9761
rect 9862 9687 9918 9696
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9678 9208 9734 9217
rect 9678 9143 9734 9152
rect 9862 9208 9918 9217
rect 9862 9143 9918 9152
rect 9678 9072 9734 9081
rect 9678 9007 9734 9016
rect 9692 8906 9720 9007
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9772 8832 9824 8838
rect 9876 8809 9904 9143
rect 9772 8774 9824 8780
rect 9862 8800 9918 8809
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9600 7177 9628 7822
rect 9586 7168 9642 7177
rect 9586 7103 9642 7112
rect 9600 7002 9628 7103
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9508 5522 9536 6938
rect 9586 6896 9642 6905
rect 9586 6831 9642 6840
rect 9600 6662 9628 6831
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9600 6390 9628 6598
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9692 6225 9720 8570
rect 9784 8265 9812 8774
rect 9862 8735 9918 8744
rect 9968 8514 9996 14214
rect 10046 12472 10102 12481
rect 10046 12407 10102 12416
rect 10060 12073 10088 12407
rect 10152 12374 10180 15370
rect 10336 14822 10364 15438
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10140 12368 10192 12374
rect 10336 12345 10364 14758
rect 10140 12310 10192 12316
rect 10322 12336 10378 12345
rect 10322 12271 10378 12280
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10140 12096 10192 12102
rect 10046 12064 10102 12073
rect 10140 12038 10192 12044
rect 10046 11999 10102 12008
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10060 10713 10088 11766
rect 10046 10704 10102 10713
rect 10046 10639 10102 10648
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9876 8486 9996 8514
rect 9770 8256 9826 8265
rect 9770 8191 9826 8200
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9678 6216 9734 6225
rect 9678 6151 9734 6160
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9508 5494 9628 5522
rect 9494 5400 9550 5409
rect 9494 5335 9550 5344
rect 9402 5264 9458 5273
rect 9312 5228 9364 5234
rect 9508 5234 9536 5335
rect 9402 5199 9458 5208
rect 9496 5228 9548 5234
rect 9312 5170 9364 5176
rect 9496 5170 9548 5176
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9140 4440 9260 4468
rect 9232 3602 9260 4440
rect 9324 4146 9352 5170
rect 9404 5024 9456 5030
rect 9600 4978 9628 5494
rect 9404 4966 9456 4972
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9416 4010 9444 4966
rect 9508 4950 9628 4978
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9402 3904 9458 3913
rect 9508 3890 9536 4950
rect 9586 4856 9642 4865
rect 9692 4826 9720 5578
rect 9784 5574 9812 8026
rect 9876 7410 9904 8486
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9876 5522 9904 7346
rect 9968 5778 9996 8298
rect 10060 8090 10088 9930
rect 10152 9353 10180 12038
rect 10230 11112 10286 11121
rect 10230 11047 10286 11056
rect 10244 10062 10272 11047
rect 10336 10810 10364 12174
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10336 9908 10364 10746
rect 10428 10062 10456 14758
rect 10520 12102 10548 14962
rect 10612 13025 10640 15506
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10598 13016 10654 13025
rect 10598 12951 10654 12960
rect 10704 12434 10732 15030
rect 10796 14618 10824 15098
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10888 14278 10916 15030
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 10980 14414 11008 14962
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 13297 10916 14214
rect 10874 13288 10930 13297
rect 10784 13252 10836 13258
rect 10874 13223 10930 13232
rect 10784 13194 10836 13200
rect 10796 12753 10824 13194
rect 10782 12744 10838 12753
rect 10782 12679 10838 12688
rect 10888 12442 10916 13223
rect 10876 12436 10928 12442
rect 10704 12406 10824 12434
rect 10598 12336 10654 12345
rect 10598 12271 10654 12280
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10612 10792 10640 12271
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10520 10764 10640 10792
rect 10520 10538 10548 10764
rect 10704 10742 10732 11494
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10336 9880 10456 9908
rect 10324 9648 10376 9654
rect 10322 9616 10324 9625
rect 10376 9616 10378 9625
rect 10322 9551 10378 9560
rect 10232 9376 10284 9382
rect 10138 9344 10194 9353
rect 10232 9318 10284 9324
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10138 9279 10194 9288
rect 10244 9178 10272 9318
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10152 8906 10180 9114
rect 10140 8900 10192 8906
rect 10336 8888 10364 9318
rect 10140 8842 10192 8848
rect 10244 8860 10364 8888
rect 10244 8616 10272 8860
rect 10428 8786 10456 9880
rect 10152 8588 10272 8616
rect 10336 8758 10456 8786
rect 10152 8537 10180 8588
rect 10138 8528 10194 8537
rect 10138 8463 10194 8472
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10244 8294 10272 8434
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 10060 7546 10088 7890
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10152 7478 10180 7822
rect 10140 7472 10192 7478
rect 10046 7440 10102 7449
rect 10140 7414 10192 7420
rect 10046 7375 10048 7384
rect 10100 7375 10102 7384
rect 10048 7346 10100 7352
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9876 5494 9996 5522
rect 9862 5400 9918 5409
rect 9862 5335 9864 5344
rect 9916 5335 9918 5344
rect 9864 5306 9916 5312
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9586 4791 9642 4800
rect 9680 4820 9732 4826
rect 9600 4622 9628 4791
rect 9680 4762 9732 4768
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9784 4690 9812 4762
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9600 4440 9720 4468
rect 9600 4146 9628 4440
rect 9692 4434 9720 4440
rect 9784 4434 9812 4490
rect 9692 4406 9812 4434
rect 9876 4321 9904 5102
rect 9862 4312 9918 4321
rect 9862 4247 9918 4256
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 4010 9628 4082
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9680 3936 9732 3942
rect 9508 3884 9680 3890
rect 9508 3878 9732 3884
rect 9508 3862 9720 3878
rect 9402 3839 9458 3848
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9140 3194 9168 3538
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9232 3126 9260 3334
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9416 2446 9444 3839
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9876 3194 9904 3674
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9876 3058 9904 3130
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9680 2576 9732 2582
rect 9678 2544 9680 2553
rect 9732 2544 9734 2553
rect 9968 2514 9996 5494
rect 10060 2990 10088 7346
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10152 3534 10180 7142
rect 10232 6384 10284 6390
rect 10336 6372 10364 8758
rect 10414 8664 10470 8673
rect 10520 8650 10548 10202
rect 10470 8622 10548 8650
rect 10414 8599 10470 8608
rect 10428 8430 10456 8599
rect 10612 8548 10640 10610
rect 10704 9994 10732 10678
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10704 8945 10732 9046
rect 10690 8936 10746 8945
rect 10796 8922 10824 12406
rect 10876 12378 10928 12384
rect 10980 12238 11008 14350
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10888 10713 10916 12106
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11150 11008 12038
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10874 10704 10930 10713
rect 10874 10639 10930 10648
rect 11072 10305 11100 14826
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 13462 11192 13670
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11164 12152 11192 12718
rect 11244 12640 11296 12646
rect 11242 12608 11244 12617
rect 11296 12608 11298 12617
rect 11242 12543 11298 12552
rect 11164 12124 11284 12152
rect 11150 12064 11206 12073
rect 11150 11999 11206 12008
rect 11164 11286 11192 11999
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11058 10296 11114 10305
rect 11058 10231 11114 10240
rect 11058 10160 11114 10169
rect 11058 10095 11060 10104
rect 11112 10095 11114 10104
rect 11060 10066 11112 10072
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9081 11100 9930
rect 11058 9072 11114 9081
rect 11058 9007 11114 9016
rect 10874 8936 10930 8945
rect 10796 8894 10874 8922
rect 10690 8871 10746 8880
rect 11072 8922 11100 9007
rect 10874 8871 10930 8880
rect 10980 8894 11100 8922
rect 10980 8634 11008 8894
rect 11164 8838 11192 11222
rect 11256 10033 11284 12124
rect 11242 10024 11298 10033
rect 11242 9959 11244 9968
rect 11296 9959 11298 9968
rect 11244 9930 11296 9936
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10520 8520 10640 8548
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10520 7750 10548 8520
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 8129 10732 8434
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10690 8120 10746 8129
rect 10690 8055 10746 8064
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 7478 10548 7686
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10416 6384 10468 6390
rect 10284 6344 10416 6372
rect 10232 6326 10284 6332
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5030 10272 6054
rect 10336 5914 10364 6344
rect 10416 6326 10468 6332
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10428 5778 10456 6122
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10428 5574 10456 5714
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 3058 10180 3334
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 10244 2854 10272 4422
rect 10336 3738 10364 5510
rect 10414 4992 10470 5001
rect 10414 4927 10470 4936
rect 10428 4321 10456 4927
rect 10414 4312 10470 4321
rect 10414 4247 10470 4256
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10520 3058 10548 7414
rect 10612 4706 10640 7482
rect 10796 4826 10824 8366
rect 10888 6662 10916 8570
rect 11164 8430 11192 8774
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10888 5914 10916 6258
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10874 5264 10930 5273
rect 10874 5199 10930 5208
rect 10888 5030 10916 5199
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10612 4678 10824 4706
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 4282 10732 4558
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10796 2990 10824 4678
rect 10888 4554 10916 4966
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10888 3534 10916 4014
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10980 3194 11008 7686
rect 11164 7410 11192 7686
rect 11256 7410 11284 9454
rect 11348 8566 11376 14010
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 13190 11468 13262
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11440 11937 11468 13126
rect 11532 12434 11560 14758
rect 11624 13705 11652 14758
rect 11610 13696 11666 13705
rect 11610 13631 11666 13640
rect 11716 12850 11744 14962
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 12360 14550 12388 14826
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12360 13938 12388 14350
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13326 11836 13670
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 12360 13410 12388 13874
rect 12268 13382 12388 13410
rect 12452 13410 12480 15302
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12544 14074 12572 14826
rect 13082 14512 13138 14521
rect 13082 14447 13138 14456
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12452 13382 12572 13410
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 12268 13258 12296 13382
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12254 13016 12310 13025
rect 12254 12951 12310 12960
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11716 12714 11744 12786
rect 12268 12714 12296 12951
rect 12360 12918 12388 13194
rect 12348 12912 12400 12918
rect 12452 12889 12480 13194
rect 12348 12854 12400 12860
rect 12438 12880 12494 12889
rect 12438 12815 12494 12824
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 11980 12436 12032 12442
rect 11532 12406 11928 12434
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11426 11928 11482 11937
rect 11532 11898 11560 12174
rect 11796 12096 11848 12102
rect 11794 12064 11796 12073
rect 11848 12064 11850 12073
rect 11794 11999 11850 12008
rect 11426 11863 11482 11872
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11440 7426 11468 11562
rect 11532 11218 11560 11698
rect 11610 11384 11666 11393
rect 11610 11319 11666 11328
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11532 10674 11560 11154
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 10062 11560 10406
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11532 9586 11560 9998
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11520 8968 11572 8974
rect 11518 8936 11520 8945
rect 11572 8936 11574 8945
rect 11518 8871 11574 8880
rect 11518 8664 11574 8673
rect 11624 8634 11652 11319
rect 11716 10198 11744 11698
rect 11900 11676 11928 12406
rect 11980 12378 12032 12384
rect 11992 12345 12020 12378
rect 11978 12336 12034 12345
rect 11978 12271 12034 12280
rect 12544 12238 12572 13382
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 12532 12232 12584 12238
rect 12070 12200 12126 12209
rect 12900 12232 12952 12238
rect 12532 12174 12584 12180
rect 12898 12200 12900 12209
rect 12952 12200 12954 12209
rect 12070 12135 12126 12144
rect 12898 12135 12954 12144
rect 12084 11898 12112 12135
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11808 11648 11928 11676
rect 11808 10248 11836 11648
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 12912 11286 12940 11494
rect 12900 11280 12952 11286
rect 12438 11248 12494 11257
rect 13004 11257 13032 12038
rect 13096 11286 13124 14447
rect 13188 12646 13216 15302
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 13938 13308 14418
rect 13450 14376 13506 14385
rect 13450 14311 13506 14320
rect 13464 13938 13492 14311
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 14006 13584 14214
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 12322 13216 12582
rect 13280 12442 13308 12922
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13266 12336 13322 12345
rect 13188 12294 13266 12322
rect 13266 12271 13322 12280
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13280 11558 13308 12174
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13084 11280 13136 11286
rect 12900 11222 12952 11228
rect 12990 11248 13046 11257
rect 12438 11183 12440 11192
rect 12492 11183 12494 11192
rect 12532 11212 12584 11218
rect 12440 11154 12492 11160
rect 12808 11212 12860 11218
rect 12584 11172 12808 11200
rect 12532 11154 12584 11160
rect 13084 11222 13136 11228
rect 12990 11183 13046 11192
rect 12808 11154 12860 11160
rect 12256 11076 12308 11082
rect 12452 11064 12480 11154
rect 12992 11144 13044 11150
rect 13268 11144 13320 11150
rect 13044 11104 13216 11132
rect 12992 11086 13044 11092
rect 12808 11076 12860 11082
rect 12452 11036 12808 11064
rect 12256 11018 12308 11024
rect 12808 11018 12860 11024
rect 12268 10452 12296 11018
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12346 10840 12402 10849
rect 12610 10843 12918 10852
rect 12346 10775 12402 10784
rect 12532 10804 12584 10810
rect 12360 10742 12388 10775
rect 12532 10746 12584 10752
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12544 10674 12572 10746
rect 12714 10704 12770 10713
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12532 10668 12584 10674
rect 12714 10639 12716 10648
rect 12532 10610 12584 10616
rect 12768 10639 12770 10648
rect 12716 10610 12768 10616
rect 12452 10470 12480 10610
rect 12624 10600 12676 10606
rect 12530 10568 12586 10577
rect 12624 10542 12676 10548
rect 12530 10503 12532 10512
rect 12584 10503 12586 10512
rect 12532 10474 12584 10480
rect 12440 10464 12492 10470
rect 12268 10424 12388 10452
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 11808 10220 11928 10248
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11518 8599 11574 8608
rect 11612 8628 11664 8634
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11348 7398 11468 7426
rect 11164 6610 11192 7346
rect 11072 6582 11192 6610
rect 11072 5817 11100 6582
rect 11242 6488 11298 6497
rect 11242 6423 11298 6432
rect 11152 5840 11204 5846
rect 11058 5808 11114 5817
rect 11152 5782 11204 5788
rect 11058 5743 11114 5752
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11072 4690 11100 5102
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11072 4457 11100 4490
rect 11058 4448 11114 4457
rect 11058 4383 11114 4392
rect 11058 4176 11114 4185
rect 11058 4111 11114 4120
rect 11072 3466 11100 4111
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11164 3126 11192 5782
rect 11256 4690 11284 6423
rect 11348 5166 11376 7398
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11440 7041 11468 7278
rect 11426 7032 11482 7041
rect 11426 6967 11428 6976
rect 11480 6967 11482 6976
rect 11428 6938 11480 6944
rect 11440 6798 11468 6938
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11440 5778 11468 6734
rect 11532 5846 11560 8599
rect 11612 8570 11664 8576
rect 11610 6896 11666 6905
rect 11610 6831 11666 6840
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11624 5658 11652 6831
rect 11716 6730 11744 9862
rect 11808 7478 11836 9862
rect 11900 9489 11928 10220
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11886 9480 11942 9489
rect 11886 9415 11942 9424
rect 12084 9382 12112 9590
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 11886 9072 11942 9081
rect 11886 9007 11942 9016
rect 11900 8974 11928 9007
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 11978 8800 12034 8809
rect 11978 8735 12034 8744
rect 11992 8430 12020 8735
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12268 8276 12296 8910
rect 12360 8634 12388 10424
rect 12440 10406 12492 10412
rect 12452 9674 12480 10406
rect 12636 10198 12664 10542
rect 13004 10266 13032 10950
rect 13188 10418 13216 11104
rect 13268 11086 13320 11092
rect 13280 10674 13308 11086
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13188 10390 13308 10418
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12990 10160 13046 10169
rect 12990 10095 12992 10104
rect 13044 10095 13046 10104
rect 12992 10066 13044 10072
rect 12624 10056 12676 10062
rect 12676 10004 13216 10010
rect 12624 9998 13216 10004
rect 12636 9982 13216 9998
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 12452 9646 12572 9674
rect 12544 9636 12572 9646
rect 12544 9608 12664 9636
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12452 9489 12480 9522
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12452 8566 12480 9046
rect 12636 8956 12664 9608
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12728 9382 12756 9522
rect 12820 9450 12848 9522
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12544 8928 12664 8956
rect 12544 8616 12572 8928
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 12544 8588 12664 8616
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12268 8248 12388 8276
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11900 7750 11928 8026
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 12360 7342 12388 8248
rect 12452 8022 12480 8366
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11808 6458 11836 7278
rect 12256 7200 12308 7206
rect 12308 7160 12388 7188
rect 12256 7142 12308 7148
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11900 6322 11928 6802
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12176 6322 12204 6734
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11794 6216 11850 6225
rect 11716 5914 11744 6190
rect 11794 6151 11850 6160
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11808 5710 11836 6151
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 11978 5808 12034 5817
rect 11888 5772 11940 5778
rect 11978 5743 12034 5752
rect 11888 5714 11940 5720
rect 11796 5704 11848 5710
rect 11532 5630 11652 5658
rect 11702 5672 11758 5681
rect 11336 5160 11388 5166
rect 11532 5114 11560 5630
rect 11796 5646 11848 5652
rect 11702 5607 11758 5616
rect 11716 5574 11744 5607
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11794 5536 11850 5545
rect 11336 5102 11388 5108
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11348 4298 11376 5102
rect 11256 4270 11376 4298
rect 11440 5086 11560 5114
rect 11256 3398 11284 4270
rect 11440 4146 11468 5086
rect 11520 4616 11572 4622
rect 11624 4604 11652 5510
rect 11794 5471 11850 5480
rect 11808 5302 11836 5471
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11900 5234 11928 5714
rect 11992 5302 12020 5743
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11900 5114 11928 5170
rect 11572 4576 11652 4604
rect 11716 5086 11928 5114
rect 11520 4558 11572 4564
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11440 3466 11468 3946
rect 11624 3641 11652 4218
rect 11610 3632 11666 3641
rect 11610 3567 11666 3576
rect 11518 3496 11574 3505
rect 11428 3460 11480 3466
rect 11518 3431 11574 3440
rect 11428 3402 11480 3408
rect 11532 3398 11560 3431
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11152 3120 11204 3126
rect 10966 3088 11022 3097
rect 11152 3062 11204 3068
rect 11716 3058 11744 5086
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4282 11836 4966
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11900 3924 11928 4558
rect 12176 4321 12204 4626
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12162 4312 12218 4321
rect 12162 4247 12218 4256
rect 12268 4214 12296 4558
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 11808 3896 11928 3924
rect 11808 3466 11836 3896
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 12360 3398 12388 7160
rect 12452 6866 12480 7686
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12452 6202 12480 6802
rect 12544 6390 12572 8298
rect 12636 7750 12664 8588
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 12714 7440 12770 7449
rect 12714 7375 12770 7384
rect 12898 7440 12954 7449
rect 12898 7375 12900 7384
rect 12728 7256 12756 7375
rect 12952 7375 12954 7384
rect 12900 7346 12952 7352
rect 12808 7268 12860 7274
rect 12728 7228 12808 7256
rect 12808 7210 12860 7216
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12452 6174 12572 6202
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12452 4282 12480 5306
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12544 3942 12572 6174
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 13004 5302 13032 8842
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 13096 5166 13124 9862
rect 13084 5160 13136 5166
rect 12898 5128 12954 5137
rect 13084 5102 13136 5108
rect 12898 5063 12954 5072
rect 12912 4622 12940 5063
rect 12900 4616 12952 4622
rect 13188 4570 13216 9982
rect 13280 9625 13308 10390
rect 13372 10266 13400 13806
rect 13556 13734 13584 13942
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13542 13424 13598 13433
rect 13542 13359 13598 13368
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13464 11898 13492 12106
rect 13556 12102 13584 13359
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13464 11626 13492 11834
rect 13740 11642 13768 15506
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 13912 15360 13964 15366
rect 13910 15328 13912 15337
rect 13964 15328 13966 15337
rect 13910 15263 13966 15272
rect 14292 15162 14320 15438
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 14006 13860 14214
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13648 11614 13768 11642
rect 13648 11082 13676 11614
rect 13832 11200 13860 11766
rect 13740 11172 13860 11200
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13464 10266 13492 10610
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13464 10169 13492 10202
rect 13450 10160 13506 10169
rect 13360 10124 13412 10130
rect 13450 10095 13506 10104
rect 13360 10066 13412 10072
rect 13266 9616 13322 9625
rect 13266 9551 13322 9560
rect 13372 9466 13400 10066
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 13280 9438 13400 9466
rect 13280 9382 13308 9438
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13360 9376 13412 9382
rect 13464 9330 13492 9930
rect 13412 9324 13492 9330
rect 13360 9318 13492 9324
rect 13280 5030 13308 9318
rect 13372 9302 13492 9318
rect 13372 6769 13400 9302
rect 13452 8968 13504 8974
rect 13556 8956 13584 11018
rect 13740 10810 13768 11172
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13504 8928 13584 8956
rect 13452 8910 13504 8916
rect 13464 8362 13492 8910
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13464 7546 13492 7754
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13358 6760 13414 6769
rect 13358 6695 13414 6704
rect 13464 6458 13492 7346
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13372 4826 13400 5850
rect 13450 5400 13506 5409
rect 13450 5335 13506 5344
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13464 4690 13492 5335
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 12900 4558 12952 4564
rect 13004 4542 13216 4570
rect 13268 4548 13320 4554
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 13004 3670 13032 4542
rect 13268 4490 13320 4496
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4078 13216 4422
rect 13176 4072 13228 4078
rect 13082 4040 13138 4049
rect 13176 4014 13228 4020
rect 13082 3975 13138 3984
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 10966 3023 11022 3032
rect 11704 3052 11756 3058
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10874 2544 10930 2553
rect 9678 2479 9734 2488
rect 9956 2508 10008 2514
rect 10874 2479 10930 2488
rect 9956 2450 10008 2456
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 7380 2372 7432 2378
rect 7380 2314 7432 2320
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 8036 2038 8064 2382
rect 9140 2038 9168 2382
rect 10888 2378 10916 2479
rect 10980 2378 11008 3023
rect 11704 2994 11756 3000
rect 11518 2680 11574 2689
rect 11518 2615 11574 2624
rect 11532 2582 11560 2615
rect 11808 2582 11836 3130
rect 12360 2990 12388 3334
rect 12452 3194 12480 3538
rect 13096 3534 13124 3975
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12716 3392 12768 3398
rect 12544 3352 12716 3380
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12348 2984 12400 2990
rect 12544 2961 12572 3352
rect 12716 3334 12768 3340
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 12348 2926 12400 2932
rect 12530 2952 12586 2961
rect 12530 2887 12586 2896
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 8024 2032 8076 2038
rect 8024 1974 8076 1980
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 9600 1902 9628 2246
rect 10152 2038 10180 2246
rect 10140 2032 10192 2038
rect 10140 1974 10192 1980
rect 9588 1896 9640 1902
rect 9588 1838 9640 1844
rect 11256 1698 11284 2246
rect 11716 1873 11744 2382
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12544 2106 12572 2246
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 12532 2100 12584 2106
rect 12532 2042 12584 2048
rect 11702 1864 11758 1873
rect 11702 1799 11758 1808
rect 13004 1737 13032 3470
rect 13188 2038 13216 3878
rect 13280 3126 13308 4490
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 13372 2972 13400 4082
rect 13450 4040 13506 4049
rect 13450 3975 13452 3984
rect 13504 3975 13506 3984
rect 13452 3946 13504 3952
rect 13464 3602 13492 3946
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13280 2944 13400 2972
rect 13280 2514 13308 2944
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13372 2582 13400 2790
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13280 2417 13308 2450
rect 13556 2446 13584 8774
rect 13648 7274 13676 10610
rect 13740 9586 13768 10746
rect 13832 9994 13860 11018
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13634 6896 13690 6905
rect 13634 6831 13690 6840
rect 13648 6322 13676 6831
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 2650 13676 6122
rect 13740 5114 13768 8570
rect 13832 5234 13860 9318
rect 13924 8634 13952 14282
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 14016 9897 14044 13942
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14108 13326 14136 13670
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14094 13152 14150 13161
rect 14094 13087 14150 13096
rect 14108 12986 14136 13087
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14002 9888 14058 9897
rect 14002 9823 14058 9832
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13924 8294 13952 8434
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7546 13952 8230
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13740 5086 13860 5114
rect 13832 4434 13860 5086
rect 13924 4729 13952 7346
rect 14016 4758 14044 9658
rect 14108 8634 14136 12786
rect 14200 9518 14228 13874
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14292 10674 14320 11698
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 9654 14320 10610
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14278 9480 14334 9489
rect 14278 9415 14334 9424
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14094 8392 14150 8401
rect 14094 8327 14150 8336
rect 14108 5846 14136 8327
rect 14292 8090 14320 9415
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14186 7576 14242 7585
rect 14186 7511 14188 7520
rect 14240 7511 14242 7520
rect 14188 7482 14240 7488
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14200 6633 14228 7142
rect 14186 6624 14242 6633
rect 14186 6559 14242 6568
rect 14292 6118 14320 7822
rect 14384 7562 14412 15574
rect 14476 15026 14504 16351
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14464 14272 14516 14278
rect 14462 14240 14464 14249
rect 14516 14240 14518 14249
rect 14462 14175 14518 14184
rect 14464 12096 14516 12102
rect 14462 12064 14464 12073
rect 14516 12064 14518 12073
rect 14462 11999 14518 12008
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14476 10985 14504 11018
rect 14462 10976 14518 10985
rect 14462 10911 14518 10920
rect 14464 9920 14516 9926
rect 14462 9888 14464 9897
rect 14516 9888 14518 9897
rect 14462 9823 14518 9832
rect 14464 8832 14516 8838
rect 14462 8800 14464 8809
rect 14516 8800 14518 8809
rect 14462 8735 14518 8744
rect 14464 7744 14516 7750
rect 14462 7712 14464 7721
rect 14516 7712 14518 7721
rect 14462 7647 14518 7656
rect 14384 7534 14504 7562
rect 14370 7032 14426 7041
rect 14476 7002 14504 7534
rect 14370 6967 14426 6976
rect 14464 6996 14516 7002
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 4826 14136 5510
rect 14200 5370 14228 5714
rect 14278 5400 14334 5409
rect 14188 5364 14240 5370
rect 14278 5335 14334 5344
rect 14188 5306 14240 5312
rect 14292 5302 14320 5335
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 14096 4820 14148 4826
rect 14148 4780 14228 4808
rect 14096 4762 14148 4768
rect 14004 4752 14056 4758
rect 13910 4720 13966 4729
rect 14004 4694 14056 4700
rect 13910 4655 13966 4664
rect 13912 4480 13964 4486
rect 13740 4406 13860 4434
rect 13910 4448 13912 4457
rect 13964 4448 13966 4457
rect 13740 3126 13768 4406
rect 13910 4383 13966 4392
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13544 2440 13596 2446
rect 13266 2408 13322 2417
rect 13544 2382 13596 2388
rect 13266 2343 13322 2352
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13176 2032 13228 2038
rect 13176 1974 13228 1980
rect 12990 1728 13046 1737
rect 6736 1692 6788 1698
rect 6736 1634 6788 1640
rect 11244 1692 11296 1698
rect 12990 1663 13046 1672
rect 11244 1634 11296 1640
rect 13648 1193 13676 2246
rect 13832 1601 13860 3946
rect 13924 3369 13952 4218
rect 14200 4214 14228 4780
rect 14384 4706 14412 6967
rect 14464 6938 14516 6944
rect 14462 5536 14518 5545
rect 14462 5471 14518 5480
rect 14476 4826 14504 5471
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14292 4678 14412 4706
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 4049 14136 4082
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 14096 3664 14148 3670
rect 14094 3632 14096 3641
rect 14148 3632 14150 3641
rect 14094 3567 14150 3576
rect 14200 3534 14228 4150
rect 14292 3738 14320 4678
rect 14370 4584 14426 4593
rect 14370 4519 14426 4528
rect 14384 4146 14412 4519
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 13910 3360 13966 3369
rect 13910 3295 13966 3304
rect 14568 2990 14596 15642
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14660 10606 14688 13262
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14752 8294 14780 15914
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14738 7304 14794 7313
rect 14648 7268 14700 7274
rect 14738 7239 14794 7248
rect 14648 7210 14700 7216
rect 14660 4214 14688 7210
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14752 3398 14780 7239
rect 14844 4622 14872 12582
rect 14936 11898 14964 15098
rect 15304 12434 15332 15370
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15120 12406 15332 12434
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 15028 11778 15056 12310
rect 14936 11750 15056 11778
rect 14936 5778 14964 11750
rect 15120 11665 15148 12406
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15106 11656 15162 11665
rect 15106 11591 15162 11600
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 15028 4185 15056 10406
rect 15120 6866 15148 11591
rect 15212 8634 15240 11834
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15304 6390 15332 9522
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15014 4176 15070 4185
rect 15014 4111 15070 4120
rect 15672 3602 15700 13806
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 13912 2304 13964 2310
rect 13910 2272 13912 2281
rect 13964 2272 13966 2281
rect 13910 2207 13966 2216
rect 13818 1592 13874 1601
rect 13818 1527 13874 1536
rect 13634 1184 13690 1193
rect 13634 1119 13690 1128
<< via2 >>
rect 14462 16360 14518 16416
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 2318 15544 2374 15600
rect 754 9968 810 10024
rect 1398 13368 1454 13424
rect 1030 12280 1086 12336
rect 938 4120 994 4176
rect 1122 3440 1178 3496
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 1582 14456 1638 14512
rect 1766 13912 1822 13968
rect 1766 13812 1768 13832
rect 1768 13812 1820 13832
rect 1820 13812 1822 13832
rect 1766 13776 1822 13812
rect 1398 11192 1454 11248
rect 1306 9560 1362 9616
rect 1766 11736 1822 11792
rect 1674 10648 1730 10704
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 1858 8336 1914 8392
rect 3606 15408 3662 15464
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 2410 10648 2466 10704
rect 2410 10376 2466 10432
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2410 8064 2466 8120
rect 1766 7420 1768 7440
rect 1768 7420 1820 7440
rect 1820 7420 1822 7440
rect 1766 7384 1822 7420
rect 1858 7248 1914 7304
rect 2318 7248 2374 7304
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 2778 11756 2834 11792
rect 2778 11736 2780 11756
rect 2780 11736 2832 11756
rect 2832 11736 2834 11756
rect 2594 11348 2650 11384
rect 2594 11328 2596 11348
rect 2596 11328 2648 11348
rect 2648 11328 2650 11348
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 2962 10104 3018 10160
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 2870 9152 2926 9208
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 3330 13368 3386 13424
rect 3606 13268 3608 13288
rect 3608 13268 3660 13288
rect 3660 13268 3662 13288
rect 3606 13232 3662 13268
rect 3514 11736 3570 11792
rect 3790 11600 3846 11656
rect 3422 11056 3478 11112
rect 3054 8744 3110 8800
rect 3054 8372 3056 8392
rect 3056 8372 3108 8392
rect 3108 8372 3110 8392
rect 3054 8336 3110 8372
rect 3054 6860 3110 6896
rect 3054 6840 3056 6860
rect 3056 6840 3108 6860
rect 3108 6840 3110 6860
rect 2778 6704 2834 6760
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2962 5752 3018 5808
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 2410 3848 2466 3904
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 3146 5888 3202 5944
rect 3330 8200 3386 8256
rect 3422 7928 3478 7984
rect 3330 6432 3386 6488
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 3238 5616 3294 5672
rect 3606 11056 3662 11112
rect 4250 14900 4252 14920
rect 4252 14900 4304 14920
rect 4304 14900 4306 14920
rect 4250 14864 4306 14900
rect 3974 13096 4030 13152
rect 4342 12960 4398 13016
rect 4342 12416 4398 12472
rect 3974 11328 4030 11384
rect 3790 8608 3846 8664
rect 3606 6568 3662 6624
rect 4250 10920 4306 10976
rect 4158 9424 4214 9480
rect 3974 8200 4030 8256
rect 3882 6160 3938 6216
rect 4158 8336 4214 8392
rect 4802 13948 4804 13968
rect 4804 13948 4856 13968
rect 4856 13948 4858 13968
rect 4802 13912 4858 13948
rect 4526 13776 4582 13832
rect 4526 12960 4582 13016
rect 4710 13132 4712 13152
rect 4712 13132 4764 13152
rect 4764 13132 4766 13152
rect 4710 13096 4766 13132
rect 5078 14184 5134 14240
rect 4986 12688 5042 12744
rect 4710 11772 4712 11792
rect 4712 11772 4764 11792
rect 4764 11772 4766 11792
rect 4710 11736 4766 11772
rect 4710 10376 4766 10432
rect 4526 9696 4582 9752
rect 4434 9288 4490 9344
rect 4434 9052 4436 9072
rect 4436 9052 4488 9072
rect 4488 9052 4490 9072
rect 4434 9016 4490 9052
rect 4434 7656 4490 7712
rect 4802 9288 4858 9344
rect 4158 5752 4214 5808
rect 3974 5480 4030 5536
rect 3790 5208 3846 5264
rect 3698 5072 3754 5128
rect 3606 3576 3662 3632
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 4434 6296 4490 6352
rect 4526 5208 4582 5264
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 2502 1944 2558 2000
rect 5630 13776 5686 13832
rect 5170 10920 5226 10976
rect 5538 12552 5594 12608
rect 5354 12280 5410 12336
rect 5354 11212 5410 11248
rect 5354 11192 5356 11212
rect 5356 11192 5408 11212
rect 5408 11192 5410 11212
rect 5538 10920 5594 10976
rect 5078 10376 5134 10432
rect 5722 11328 5778 11384
rect 5446 9832 5502 9888
rect 4986 8608 5042 8664
rect 5446 8608 5502 8664
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 6090 14220 6092 14240
rect 6092 14220 6144 14240
rect 6144 14220 6146 14240
rect 6090 14184 6146 14220
rect 6182 13912 6238 13968
rect 6182 12144 6238 12200
rect 5630 8608 5686 8664
rect 4986 7928 5042 7984
rect 4986 7520 5042 7576
rect 4986 6840 5042 6896
rect 5630 6704 5686 6760
rect 5446 5636 5502 5672
rect 5446 5616 5448 5636
rect 5448 5616 5500 5636
rect 5500 5616 5502 5636
rect 5354 4700 5356 4720
rect 5356 4700 5408 4720
rect 5408 4700 5410 4720
rect 5354 4664 5410 4700
rect 6366 11872 6422 11928
rect 6182 11192 6238 11248
rect 6090 10240 6146 10296
rect 6734 12552 6790 12608
rect 6734 12416 6790 12472
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 7194 13232 7250 13288
rect 7286 13096 7342 13152
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 6642 12144 6698 12200
rect 6918 11872 6974 11928
rect 7102 12008 7158 12064
rect 6366 10668 6422 10704
rect 6366 10648 6368 10668
rect 6368 10648 6420 10668
rect 6420 10648 6422 10668
rect 6274 10104 6330 10160
rect 6458 10104 6514 10160
rect 6642 10648 6698 10704
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 6918 11192 6974 11248
rect 7102 11192 7158 11248
rect 7194 10920 7250 10976
rect 7010 10784 7066 10840
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 8114 14048 8170 14104
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 7470 12960 7526 13016
rect 7562 12416 7618 12472
rect 8758 14184 8814 14240
rect 8482 13096 8538 13152
rect 8482 12688 8538 12744
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 7654 11464 7710 11520
rect 7470 11192 7526 11248
rect 7746 11192 7802 11248
rect 7378 10784 7434 10840
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 6734 10412 6736 10432
rect 6736 10412 6788 10432
rect 6788 10412 6790 10432
rect 6734 10376 6790 10412
rect 7378 10376 7434 10432
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 6734 10240 6790 10296
rect 6642 9968 6698 10024
rect 6918 9968 6974 10024
rect 6090 9288 6146 9344
rect 6366 9288 6422 9344
rect 6182 8880 6238 8936
rect 5906 7928 5962 7984
rect 5906 7248 5962 7304
rect 6182 7692 6184 7712
rect 6184 7692 6236 7712
rect 6236 7692 6238 7712
rect 6182 7656 6238 7692
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 6734 9288 6790 9344
rect 6734 9152 6790 9208
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 6918 8916 6920 8936
rect 6920 8916 6972 8936
rect 6972 8916 6974 8936
rect 6918 8880 6974 8916
rect 6274 6976 6330 7032
rect 5998 5480 6054 5536
rect 6182 5208 6238 5264
rect 4894 3032 4950 3088
rect 6458 5244 6460 5264
rect 6460 5244 6512 5264
rect 6512 5244 6514 5264
rect 6458 5208 6514 5244
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 7470 9152 7526 9208
rect 8206 12008 8262 12064
rect 8390 12008 8446 12064
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 14186 15564 14242 15600
rect 14186 15544 14188 15564
rect 14188 15544 14240 15564
rect 14240 15544 14242 15564
rect 9586 13948 9588 13968
rect 9588 13948 9640 13968
rect 9640 13948 9642 13968
rect 9586 13912 9642 13948
rect 9218 13776 9274 13832
rect 8758 12960 8814 13016
rect 8298 11872 8354 11928
rect 8574 11636 8576 11656
rect 8576 11636 8628 11656
rect 8628 11636 8630 11656
rect 8574 11600 8630 11636
rect 8390 11328 8446 11384
rect 8298 10104 8354 10160
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 7930 8200 7986 8256
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 6734 7248 6790 7304
rect 6734 7112 6790 7168
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 6826 6568 6882 6624
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 7470 6432 7526 6488
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 6550 3848 6606 3904
rect 7378 5888 7434 5944
rect 7746 6024 7802 6080
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 7562 5208 7618 5264
rect 7010 4020 7012 4040
rect 7012 4020 7064 4040
rect 7064 4020 7066 4040
rect 7010 3984 7066 4020
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 7930 4936 7986 4992
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 6826 2896 6882 2952
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 7470 3304 7526 3360
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 8206 8608 8262 8664
rect 8850 11636 8852 11656
rect 8852 11636 8904 11656
rect 8904 11636 8906 11656
rect 8850 11600 8906 11636
rect 9034 11328 9090 11384
rect 9126 9968 9182 10024
rect 9034 9288 9090 9344
rect 8482 6976 8538 7032
rect 8390 5752 8446 5808
rect 8206 4528 8262 4584
rect 8390 5344 8446 5400
rect 8666 8356 8722 8392
rect 8666 8336 8668 8356
rect 8668 8336 8720 8356
rect 8720 8336 8722 8356
rect 9126 8336 9182 8392
rect 8942 6568 8998 6624
rect 8850 6160 8906 6216
rect 8666 6024 8722 6080
rect 8574 4936 8630 4992
rect 8942 5888 8998 5944
rect 8666 3168 8722 3224
rect 9126 7792 9182 7848
rect 9126 6860 9182 6896
rect 9126 6840 9128 6860
rect 9128 6840 9180 6860
rect 9180 6840 9182 6860
rect 9126 6432 9182 6488
rect 9862 9696 9918 9752
rect 9678 9152 9734 9208
rect 9862 9152 9918 9208
rect 9678 9016 9734 9072
rect 9586 7112 9642 7168
rect 9586 6840 9642 6896
rect 9862 8744 9918 8800
rect 10046 12416 10102 12472
rect 10322 12280 10378 12336
rect 10046 12008 10102 12064
rect 10046 10648 10102 10704
rect 9770 8200 9826 8256
rect 9678 6160 9734 6216
rect 9494 5344 9550 5400
rect 9402 5208 9458 5264
rect 9402 3848 9458 3904
rect 9586 4800 9642 4856
rect 10230 11056 10286 11112
rect 10598 12960 10654 13016
rect 10874 13232 10930 13288
rect 10782 12688 10838 12744
rect 10598 12280 10654 12336
rect 10322 9596 10324 9616
rect 10324 9596 10376 9616
rect 10376 9596 10378 9616
rect 10322 9560 10378 9596
rect 10138 9288 10194 9344
rect 10138 8472 10194 8528
rect 10046 7404 10102 7440
rect 10046 7384 10048 7404
rect 10048 7384 10100 7404
rect 10100 7384 10102 7404
rect 9862 5364 9918 5400
rect 9862 5344 9864 5364
rect 9864 5344 9916 5364
rect 9916 5344 9918 5364
rect 9862 4256 9918 4312
rect 9678 2524 9680 2544
rect 9680 2524 9732 2544
rect 9732 2524 9734 2544
rect 9678 2488 9734 2524
rect 10414 8608 10470 8664
rect 10690 8880 10746 8936
rect 10874 10648 10930 10704
rect 11242 12588 11244 12608
rect 11244 12588 11296 12608
rect 11296 12588 11298 12608
rect 11242 12552 11298 12588
rect 11150 12008 11206 12064
rect 11058 10240 11114 10296
rect 11058 10124 11114 10160
rect 11058 10104 11060 10124
rect 11060 10104 11112 10124
rect 11112 10104 11114 10124
rect 11058 9016 11114 9072
rect 10874 8880 10930 8936
rect 11242 9988 11298 10024
rect 11242 9968 11244 9988
rect 11244 9968 11296 9988
rect 11296 9968 11298 9988
rect 10690 8064 10746 8120
rect 10414 4936 10470 4992
rect 10414 4256 10470 4312
rect 10874 5208 10930 5264
rect 11610 13640 11666 13696
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 13082 14456 13138 14512
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 12254 12960 12310 13016
rect 12438 12824 12494 12880
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 11426 11872 11482 11928
rect 11794 12044 11796 12064
rect 11796 12044 11848 12064
rect 11848 12044 11850 12064
rect 11794 12008 11850 12044
rect 11610 11328 11666 11384
rect 11518 8916 11520 8936
rect 11520 8916 11572 8936
rect 11572 8916 11574 8936
rect 11518 8880 11574 8916
rect 11518 8608 11574 8664
rect 11978 12280 12034 12336
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 12070 12144 12126 12200
rect 12898 12180 12900 12200
rect 12900 12180 12952 12200
rect 12952 12180 12954 12200
rect 12898 12144 12954 12180
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 12438 11212 12494 11248
rect 13450 14320 13506 14376
rect 13266 12280 13322 12336
rect 12438 11192 12440 11212
rect 12440 11192 12492 11212
rect 12492 11192 12494 11212
rect 12990 11192 13046 11248
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 12346 10784 12402 10840
rect 12714 10668 12770 10704
rect 12714 10648 12716 10668
rect 12716 10648 12768 10668
rect 12768 10648 12770 10668
rect 12530 10532 12586 10568
rect 12530 10512 12532 10532
rect 12532 10512 12584 10532
rect 12584 10512 12586 10532
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 11242 6432 11298 6488
rect 11058 5752 11114 5808
rect 11058 4392 11114 4448
rect 11058 4120 11114 4176
rect 11426 6996 11482 7032
rect 11426 6976 11428 6996
rect 11428 6976 11480 6996
rect 11480 6976 11482 6996
rect 11610 6840 11666 6896
rect 11886 9424 11942 9480
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 11886 9016 11942 9072
rect 11978 8744 12034 8800
rect 12990 10124 13046 10160
rect 12990 10104 12992 10124
rect 12992 10104 13044 10124
rect 13044 10104 13046 10124
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 12438 9424 12494 9480
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 11794 6160 11850 6216
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 11978 5752 12034 5808
rect 11702 5616 11758 5672
rect 11794 5480 11850 5536
rect 11610 3576 11666 3632
rect 11518 3440 11574 3496
rect 10966 3032 11022 3088
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 12162 4256 12218 4312
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 12714 7384 12770 7440
rect 12898 7404 12954 7440
rect 12898 7384 12900 7404
rect 12900 7384 12952 7404
rect 12952 7384 12954 7404
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 12898 5072 12954 5128
rect 13542 13368 13598 13424
rect 13910 15308 13912 15328
rect 13912 15308 13964 15328
rect 13964 15308 13966 15328
rect 13910 15272 13966 15308
rect 13450 10104 13506 10160
rect 13266 9560 13322 9616
rect 13358 6704 13414 6760
rect 13450 5344 13506 5400
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 13082 3984 13138 4040
rect 10874 2488 10930 2544
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 11518 2624 11574 2680
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 12530 2896 12586 2952
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 11702 1808 11758 1864
rect 13450 4004 13506 4040
rect 13450 3984 13452 4004
rect 13452 3984 13504 4004
rect 13504 3984 13506 4004
rect 13634 6840 13690 6896
rect 14094 13096 14150 13152
rect 14002 9832 14058 9888
rect 14278 9424 14334 9480
rect 14094 8336 14150 8392
rect 14186 7540 14242 7576
rect 14186 7520 14188 7540
rect 14188 7520 14240 7540
rect 14240 7520 14242 7540
rect 14186 6568 14242 6624
rect 14462 14220 14464 14240
rect 14464 14220 14516 14240
rect 14516 14220 14518 14240
rect 14462 14184 14518 14220
rect 14462 12044 14464 12064
rect 14464 12044 14516 12064
rect 14516 12044 14518 12064
rect 14462 12008 14518 12044
rect 14462 10920 14518 10976
rect 14462 9868 14464 9888
rect 14464 9868 14516 9888
rect 14516 9868 14518 9888
rect 14462 9832 14518 9868
rect 14462 8780 14464 8800
rect 14464 8780 14516 8800
rect 14516 8780 14518 8800
rect 14462 8744 14518 8780
rect 14462 7692 14464 7712
rect 14464 7692 14516 7712
rect 14516 7692 14518 7712
rect 14462 7656 14518 7692
rect 14370 6976 14426 7032
rect 14278 5344 14334 5400
rect 13910 4664 13966 4720
rect 13910 4428 13912 4448
rect 13912 4428 13964 4448
rect 13964 4428 13966 4448
rect 13910 4392 13966 4428
rect 13266 2352 13322 2408
rect 12990 1672 13046 1728
rect 14462 5480 14518 5536
rect 14094 3984 14150 4040
rect 14094 3612 14096 3632
rect 14096 3612 14148 3632
rect 14148 3612 14150 3632
rect 14094 3576 14150 3612
rect 14370 4528 14426 4584
rect 13910 3304 13966 3360
rect 14738 7248 14794 7304
rect 15106 11600 15162 11656
rect 15014 4120 15070 4176
rect 13910 2252 13912 2272
rect 13912 2252 13964 2272
rect 13964 2252 13966 2272
rect 13910 2216 13966 2252
rect 13818 1536 13874 1592
rect 13634 1128 13690 1184
<< metal3 >>
rect 14457 16418 14523 16421
rect 15200 16418 16000 16448
rect 14457 16416 16000 16418
rect 14457 16360 14462 16416
rect 14518 16360 16000 16416
rect 14457 16358 16000 16360
rect 14457 16355 14523 16358
rect 15200 16328 16000 16358
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 2313 15602 2379 15605
rect 14181 15602 14247 15605
rect 2313 15600 14247 15602
rect 2313 15544 2318 15600
rect 2374 15544 14186 15600
rect 14242 15544 14247 15600
rect 2313 15542 14247 15544
rect 2313 15539 2379 15542
rect 14181 15539 14247 15542
rect 3601 15466 3667 15469
rect 9254 15466 9260 15468
rect 3601 15464 9260 15466
rect 3601 15408 3606 15464
rect 3662 15408 9260 15464
rect 3601 15406 9260 15408
rect 3601 15403 3667 15406
rect 9254 15404 9260 15406
rect 9324 15404 9330 15468
rect 13905 15330 13971 15333
rect 15200 15330 16000 15360
rect 13905 15328 16000 15330
rect 13905 15272 13910 15328
rect 13966 15272 16000 15328
rect 13905 15270 16000 15272
rect 13905 15267 13971 15270
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 15200 15240 16000 15270
rect 12606 15199 12922 15200
rect 4245 14922 4311 14925
rect 10542 14922 10548 14924
rect 4245 14920 10548 14922
rect 4245 14864 4250 14920
rect 4306 14864 10548 14920
rect 4245 14862 10548 14864
rect 4245 14859 4311 14862
rect 10542 14860 10548 14862
rect 10612 14860 10618 14924
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 1577 14514 1643 14517
rect 13077 14514 13143 14517
rect 1577 14512 13143 14514
rect 1577 14456 1582 14512
rect 1638 14456 13082 14512
rect 13138 14456 13143 14512
rect 1577 14454 13143 14456
rect 1577 14451 1643 14454
rect 13077 14451 13143 14454
rect 790 14316 796 14380
rect 860 14378 866 14380
rect 13445 14378 13511 14381
rect 860 14376 13511 14378
rect 860 14320 13450 14376
rect 13506 14320 13511 14376
rect 860 14318 13511 14320
rect 860 14316 866 14318
rect 13445 14315 13511 14318
rect 5073 14242 5139 14245
rect 6085 14242 6151 14245
rect 5073 14240 6151 14242
rect 5073 14184 5078 14240
rect 5134 14184 6090 14240
rect 6146 14184 6151 14240
rect 5073 14182 6151 14184
rect 5073 14179 5139 14182
rect 6085 14179 6151 14182
rect 8753 14242 8819 14245
rect 11646 14242 11652 14244
rect 8753 14240 11652 14242
rect 8753 14184 8758 14240
rect 8814 14184 11652 14240
rect 8753 14182 11652 14184
rect 8753 14179 8819 14182
rect 11646 14180 11652 14182
rect 11716 14180 11722 14244
rect 14457 14242 14523 14245
rect 15200 14242 16000 14272
rect 14457 14240 16000 14242
rect 14457 14184 14462 14240
rect 14518 14184 16000 14240
rect 14457 14182 16000 14184
rect 14457 14179 14523 14182
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 15200 14152 16000 14182
rect 12606 14111 12922 14112
rect 8109 14106 8175 14109
rect 12382 14106 12388 14108
rect 8109 14104 12388 14106
rect 8109 14048 8114 14104
rect 8170 14048 12388 14104
rect 8109 14046 12388 14048
rect 8109 14043 8175 14046
rect 12382 14044 12388 14046
rect 12452 14044 12458 14108
rect 1158 13908 1164 13972
rect 1228 13970 1234 13972
rect 1761 13970 1827 13973
rect 1228 13968 1827 13970
rect 1228 13912 1766 13968
rect 1822 13912 1827 13968
rect 1228 13910 1827 13912
rect 1228 13908 1234 13910
rect 1761 13907 1827 13910
rect 4654 13908 4660 13972
rect 4724 13970 4730 13972
rect 4797 13970 4863 13973
rect 4724 13968 4863 13970
rect 4724 13912 4802 13968
rect 4858 13912 4863 13968
rect 4724 13910 4863 13912
rect 4724 13908 4730 13910
rect 4797 13907 4863 13910
rect 6177 13970 6243 13973
rect 9581 13970 9647 13973
rect 14038 13970 14044 13972
rect 6177 13968 9506 13970
rect 6177 13912 6182 13968
rect 6238 13912 9506 13968
rect 6177 13910 9506 13912
rect 6177 13907 6243 13910
rect 1761 13836 1827 13837
rect 1710 13834 1716 13836
rect 1670 13774 1716 13834
rect 1780 13832 1827 13836
rect 1822 13776 1827 13832
rect 1710 13772 1716 13774
rect 1780 13772 1827 13776
rect 1761 13771 1827 13772
rect 4521 13834 4587 13837
rect 5625 13836 5691 13837
rect 5390 13834 5396 13836
rect 4521 13832 5396 13834
rect 4521 13776 4526 13832
rect 4582 13776 5396 13832
rect 4521 13774 5396 13776
rect 4521 13771 4587 13774
rect 5390 13772 5396 13774
rect 5460 13772 5466 13836
rect 5574 13834 5580 13836
rect 5534 13774 5580 13834
rect 5644 13832 5691 13836
rect 5686 13776 5691 13832
rect 5574 13772 5580 13774
rect 5644 13772 5691 13776
rect 6678 13772 6684 13836
rect 6748 13834 6754 13836
rect 9213 13834 9279 13837
rect 6748 13832 9279 13834
rect 6748 13776 9218 13832
rect 9274 13776 9279 13832
rect 6748 13774 9279 13776
rect 9446 13834 9506 13910
rect 9581 13968 14044 13970
rect 9581 13912 9586 13968
rect 9642 13912 14044 13968
rect 9581 13910 14044 13912
rect 9581 13907 9647 13910
rect 14038 13908 14044 13910
rect 14108 13908 14114 13972
rect 13854 13834 13860 13836
rect 9446 13774 13860 13834
rect 6748 13772 6754 13774
rect 5625 13771 5691 13772
rect 9213 13771 9279 13774
rect 13854 13772 13860 13774
rect 13924 13772 13930 13836
rect 9806 13636 9812 13700
rect 9876 13698 9882 13700
rect 11605 13698 11671 13701
rect 9876 13696 11671 13698
rect 9876 13640 11610 13696
rect 11666 13640 11671 13696
rect 9876 13638 11671 13640
rect 9876 13636 9882 13638
rect 11605 13635 11671 13638
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 0 13426 800 13456
rect 1393 13426 1459 13429
rect 0 13424 1459 13426
rect 0 13368 1398 13424
rect 1454 13368 1459 13424
rect 0 13366 1459 13368
rect 0 13336 800 13366
rect 1393 13363 1459 13366
rect 3325 13426 3391 13429
rect 13537 13426 13603 13429
rect 3325 13424 13603 13426
rect 3325 13368 3330 13424
rect 3386 13368 13542 13424
rect 13598 13368 13603 13424
rect 3325 13366 13603 13368
rect 3325 13363 3391 13366
rect 13537 13363 13603 13366
rect 3601 13290 3667 13293
rect 7189 13290 7255 13293
rect 10869 13290 10935 13293
rect 3601 13288 10935 13290
rect 3601 13232 3606 13288
rect 3662 13232 7194 13288
rect 7250 13232 10874 13288
rect 10930 13232 10935 13288
rect 3601 13230 10935 13232
rect 3601 13227 3667 13230
rect 7189 13227 7255 13230
rect 10869 13227 10935 13230
rect 3969 13156 4035 13157
rect 3918 13154 3924 13156
rect 3878 13094 3924 13154
rect 3988 13152 4035 13156
rect 4030 13096 4035 13152
rect 3918 13092 3924 13094
rect 3988 13092 4035 13096
rect 3969 13091 4035 13092
rect 4705 13154 4771 13157
rect 5942 13154 5948 13156
rect 4705 13152 5948 13154
rect 4705 13096 4710 13152
rect 4766 13096 5948 13152
rect 4705 13094 5948 13096
rect 4705 13091 4771 13094
rect 5942 13092 5948 13094
rect 6012 13154 6018 13156
rect 7281 13154 7347 13157
rect 6012 13152 7347 13154
rect 6012 13096 7286 13152
rect 7342 13096 7347 13152
rect 6012 13094 7347 13096
rect 6012 13092 6018 13094
rect 7281 13091 7347 13094
rect 8334 13092 8340 13156
rect 8404 13154 8410 13156
rect 8477 13154 8543 13157
rect 8404 13152 8543 13154
rect 8404 13096 8482 13152
rect 8538 13096 8543 13152
rect 8404 13094 8543 13096
rect 8404 13092 8410 13094
rect 8477 13091 8543 13094
rect 14089 13154 14155 13157
rect 15200 13154 16000 13184
rect 14089 13152 16000 13154
rect 14089 13096 14094 13152
rect 14150 13096 16000 13152
rect 14089 13094 16000 13096
rect 14089 13091 14155 13094
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 15200 13064 16000 13094
rect 12606 13023 12922 13024
rect 3550 12956 3556 13020
rect 3620 13018 3626 13020
rect 4337 13018 4403 13021
rect 3620 13016 4403 13018
rect 3620 12960 4342 13016
rect 4398 12960 4403 13016
rect 3620 12958 4403 12960
rect 3620 12956 3626 12958
rect 4337 12955 4403 12958
rect 4521 13018 4587 13021
rect 7465 13018 7531 13021
rect 4521 13016 7531 13018
rect 4521 12960 4526 13016
rect 4582 12960 7470 13016
rect 7526 12960 7531 13016
rect 4521 12958 7531 12960
rect 4521 12955 4587 12958
rect 7465 12955 7531 12958
rect 8518 12956 8524 13020
rect 8588 13018 8594 13020
rect 8753 13018 8819 13021
rect 8588 13016 8819 13018
rect 8588 12960 8758 13016
rect 8814 12960 8819 13016
rect 8588 12958 8819 12960
rect 8588 12956 8594 12958
rect 8753 12955 8819 12958
rect 10593 13018 10659 13021
rect 12249 13018 12315 13021
rect 10593 13016 12315 13018
rect 10593 12960 10598 13016
rect 10654 12960 12254 13016
rect 12310 12960 12315 13016
rect 10593 12958 12315 12960
rect 10593 12955 10659 12958
rect 12249 12955 12315 12958
rect 974 12820 980 12884
rect 1044 12882 1050 12884
rect 12433 12882 12499 12885
rect 1044 12880 12499 12882
rect 1044 12824 12438 12880
rect 12494 12824 12499 12880
rect 1044 12822 12499 12824
rect 1044 12820 1050 12822
rect 12433 12819 12499 12822
rect 4981 12746 5047 12749
rect 8477 12746 8543 12749
rect 10777 12746 10843 12749
rect 4981 12744 7482 12746
rect 4981 12688 4986 12744
rect 5042 12688 7482 12744
rect 4981 12686 7482 12688
rect 4981 12683 5047 12686
rect 5533 12610 5599 12613
rect 6729 12610 6795 12613
rect 5533 12608 6795 12610
rect 5533 12552 5538 12608
rect 5594 12552 6734 12608
rect 6790 12552 6795 12608
rect 5533 12550 6795 12552
rect 7422 12610 7482 12686
rect 8477 12744 10843 12746
rect 8477 12688 8482 12744
rect 8538 12688 10782 12744
rect 10838 12688 10843 12744
rect 8477 12686 10843 12688
rect 8477 12683 8543 12686
rect 10777 12683 10843 12686
rect 11237 12610 11303 12613
rect 7422 12608 11303 12610
rect 7422 12552 11242 12608
rect 11298 12552 11303 12608
rect 7422 12550 11303 12552
rect 5533 12547 5599 12550
rect 6729 12547 6795 12550
rect 11237 12547 11303 12550
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 4337 12474 4403 12477
rect 6729 12474 6795 12477
rect 4337 12472 6795 12474
rect 4337 12416 4342 12472
rect 4398 12416 6734 12472
rect 6790 12416 6795 12472
rect 4337 12414 6795 12416
rect 4337 12411 4403 12414
rect 6729 12411 6795 12414
rect 7557 12474 7623 12477
rect 10041 12474 10107 12477
rect 7557 12472 10107 12474
rect 7557 12416 7562 12472
rect 7618 12416 10046 12472
rect 10102 12416 10107 12472
rect 7557 12414 10107 12416
rect 7557 12411 7623 12414
rect 10041 12411 10107 12414
rect 1025 12338 1091 12341
rect 5349 12338 5415 12341
rect 1025 12336 5415 12338
rect 1025 12280 1030 12336
rect 1086 12280 5354 12336
rect 5410 12280 5415 12336
rect 1025 12278 5415 12280
rect 1025 12275 1091 12278
rect 5349 12275 5415 12278
rect 6310 12276 6316 12340
rect 6380 12338 6386 12340
rect 10317 12338 10383 12341
rect 6380 12336 10383 12338
rect 6380 12280 10322 12336
rect 10378 12280 10383 12336
rect 6380 12278 10383 12280
rect 6380 12276 6386 12278
rect 10317 12275 10383 12278
rect 10593 12338 10659 12341
rect 11973 12338 12039 12341
rect 10593 12336 12039 12338
rect 10593 12280 10598 12336
rect 10654 12280 11978 12336
rect 12034 12280 12039 12336
rect 10593 12278 12039 12280
rect 10593 12275 10659 12278
rect 11973 12275 12039 12278
rect 12382 12276 12388 12340
rect 12452 12338 12458 12340
rect 13118 12338 13124 12340
rect 12452 12278 13124 12338
rect 12452 12276 12458 12278
rect 13118 12276 13124 12278
rect 13188 12276 13194 12340
rect 13261 12336 13327 12341
rect 13261 12280 13266 12336
rect 13322 12280 13327 12336
rect 13261 12275 13327 12280
rect 6177 12202 6243 12205
rect 6494 12202 6500 12204
rect 6177 12200 6500 12202
rect 6177 12144 6182 12200
rect 6238 12144 6500 12200
rect 6177 12142 6500 12144
rect 6177 12139 6243 12142
rect 6494 12140 6500 12142
rect 6564 12140 6570 12204
rect 6637 12202 6703 12205
rect 12065 12202 12131 12205
rect 6637 12200 12131 12202
rect 6637 12144 6642 12200
rect 6698 12144 12070 12200
rect 12126 12144 12131 12200
rect 6637 12142 12131 12144
rect 6637 12139 6703 12142
rect 12065 12139 12131 12142
rect 12893 12202 12959 12205
rect 13264 12202 13324 12275
rect 13486 12202 13492 12204
rect 12893 12200 13492 12202
rect 12893 12144 12898 12200
rect 12954 12144 13492 12200
rect 12893 12142 13492 12144
rect 12893 12139 12959 12142
rect 13486 12140 13492 12142
rect 13556 12140 13562 12204
rect 5022 12004 5028 12068
rect 5092 12066 5098 12068
rect 7097 12066 7163 12069
rect 8201 12068 8267 12069
rect 8150 12066 8156 12068
rect 5092 12064 7163 12066
rect 5092 12008 7102 12064
rect 7158 12008 7163 12064
rect 5092 12006 7163 12008
rect 8110 12006 8156 12066
rect 8220 12064 8267 12068
rect 8262 12008 8267 12064
rect 5092 12004 5098 12006
rect 7097 12003 7163 12006
rect 8150 12004 8156 12006
rect 8220 12004 8267 12008
rect 8201 12003 8267 12004
rect 8385 12066 8451 12069
rect 8518 12066 8524 12068
rect 8385 12064 8524 12066
rect 8385 12008 8390 12064
rect 8446 12008 8524 12064
rect 8385 12006 8524 12008
rect 8385 12003 8451 12006
rect 8518 12004 8524 12006
rect 8588 12004 8594 12068
rect 10041 12066 10107 12069
rect 11145 12066 11211 12069
rect 10041 12064 11211 12066
rect 10041 12008 10046 12064
rect 10102 12008 11150 12064
rect 11206 12008 11211 12064
rect 10041 12006 11211 12008
rect 10041 12003 10107 12006
rect 11145 12003 11211 12006
rect 11462 12004 11468 12068
rect 11532 12066 11538 12068
rect 11789 12066 11855 12069
rect 11532 12064 11855 12066
rect 11532 12008 11794 12064
rect 11850 12008 11855 12064
rect 11532 12006 11855 12008
rect 11532 12004 11538 12006
rect 11789 12003 11855 12006
rect 14457 12066 14523 12069
rect 15200 12066 16000 12096
rect 14457 12064 16000 12066
rect 14457 12008 14462 12064
rect 14518 12008 16000 12064
rect 14457 12006 16000 12008
rect 14457 12003 14523 12006
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 15200 11976 16000 12006
rect 12606 11935 12922 11936
rect 6361 11930 6427 11933
rect 6913 11930 6979 11933
rect 6361 11928 6979 11930
rect 6361 11872 6366 11928
rect 6422 11872 6918 11928
rect 6974 11872 6979 11928
rect 6361 11870 6979 11872
rect 6361 11867 6427 11870
rect 6913 11867 6979 11870
rect 8293 11932 8359 11933
rect 8293 11928 8340 11932
rect 8404 11930 8410 11932
rect 8293 11872 8298 11928
rect 8293 11868 8340 11872
rect 8404 11870 8450 11930
rect 8404 11868 8410 11870
rect 9990 11868 9996 11932
rect 10060 11930 10066 11932
rect 11421 11930 11487 11933
rect 10060 11928 11487 11930
rect 10060 11872 11426 11928
rect 11482 11872 11487 11928
rect 10060 11870 11487 11872
rect 10060 11868 10066 11870
rect 8293 11867 8359 11868
rect 11421 11867 11487 11870
rect 1761 11794 1827 11797
rect 2773 11794 2839 11797
rect 1761 11792 2839 11794
rect 1761 11736 1766 11792
rect 1822 11736 2778 11792
rect 2834 11736 2839 11792
rect 1761 11734 2839 11736
rect 1761 11731 1827 11734
rect 2773 11731 2839 11734
rect 3366 11732 3372 11796
rect 3436 11794 3442 11796
rect 3509 11794 3575 11797
rect 3436 11792 3575 11794
rect 3436 11736 3514 11792
rect 3570 11736 3575 11792
rect 3436 11734 3575 11736
rect 3436 11732 3442 11734
rect 3509 11731 3575 11734
rect 4705 11794 4771 11797
rect 13302 11794 13308 11796
rect 4705 11792 13308 11794
rect 4705 11736 4710 11792
rect 4766 11736 13308 11792
rect 4705 11734 13308 11736
rect 4705 11731 4771 11734
rect 13302 11732 13308 11734
rect 13372 11732 13378 11796
rect 1526 11596 1532 11660
rect 1596 11658 1602 11660
rect 3785 11658 3851 11661
rect 8569 11658 8635 11661
rect 1596 11656 3851 11658
rect 1596 11600 3790 11656
rect 3846 11600 3851 11656
rect 1596 11598 3851 11600
rect 1596 11596 1602 11598
rect 3785 11595 3851 11598
rect 6686 11656 8635 11658
rect 6686 11600 8574 11656
rect 8630 11600 8635 11656
rect 6686 11598 8635 11600
rect 6686 11522 6746 11598
rect 8569 11595 8635 11598
rect 8845 11658 8911 11661
rect 15101 11658 15167 11661
rect 8845 11656 15167 11658
rect 8845 11600 8850 11656
rect 8906 11600 15106 11656
rect 15162 11600 15167 11656
rect 8845 11598 15167 11600
rect 8845 11595 8911 11598
rect 15101 11595 15167 11598
rect 2730 11462 6746 11522
rect 7649 11522 7715 11525
rect 11278 11522 11284 11524
rect 7649 11520 11284 11522
rect 7649 11464 7654 11520
rect 7710 11464 11284 11520
rect 7649 11462 11284 11464
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 2589 11386 2655 11389
rect 2730 11386 2790 11462
rect 7649 11459 7715 11462
rect 11278 11460 11284 11462
rect 11348 11460 11354 11524
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 2589 11384 2790 11386
rect 2589 11328 2594 11384
rect 2650 11328 2790 11384
rect 2589 11326 2790 11328
rect 3969 11386 4035 11389
rect 4102 11386 4108 11388
rect 3969 11384 4108 11386
rect 3969 11328 3974 11384
rect 4030 11328 4108 11384
rect 3969 11326 4108 11328
rect 2589 11323 2655 11326
rect 3969 11323 4035 11326
rect 4102 11324 4108 11326
rect 4172 11324 4178 11388
rect 5574 11324 5580 11388
rect 5644 11386 5650 11388
rect 5717 11386 5783 11389
rect 5644 11384 5783 11386
rect 5644 11328 5722 11384
rect 5778 11328 5783 11384
rect 5644 11326 5783 11328
rect 5644 11324 5650 11326
rect 5717 11323 5783 11326
rect 8385 11386 8451 11389
rect 9029 11386 9095 11389
rect 8385 11384 9690 11386
rect 8385 11328 8390 11384
rect 8446 11328 9034 11384
rect 9090 11328 9690 11384
rect 8385 11326 9690 11328
rect 8385 11323 8451 11326
rect 9029 11323 9095 11326
rect 1393 11250 1459 11253
rect 5349 11250 5415 11253
rect 1393 11248 5415 11250
rect 1393 11192 1398 11248
rect 1454 11192 5354 11248
rect 5410 11192 5415 11248
rect 1393 11190 5415 11192
rect 1393 11187 1459 11190
rect 5349 11187 5415 11190
rect 6177 11250 6243 11253
rect 6913 11250 6979 11253
rect 6177 11248 6979 11250
rect 6177 11192 6182 11248
rect 6238 11192 6918 11248
rect 6974 11192 6979 11248
rect 6177 11190 6979 11192
rect 6177 11187 6243 11190
rect 6913 11187 6979 11190
rect 7097 11250 7163 11253
rect 7465 11250 7531 11253
rect 7097 11248 7531 11250
rect 7097 11192 7102 11248
rect 7158 11192 7470 11248
rect 7526 11192 7531 11248
rect 7097 11190 7531 11192
rect 7097 11187 7163 11190
rect 7465 11187 7531 11190
rect 7741 11250 7807 11253
rect 9438 11250 9444 11252
rect 7741 11248 9444 11250
rect 7741 11192 7746 11248
rect 7802 11192 9444 11248
rect 7741 11190 9444 11192
rect 7741 11187 7807 11190
rect 9438 11188 9444 11190
rect 9508 11188 9514 11252
rect 9630 11250 9690 11326
rect 10542 11324 10548 11388
rect 10612 11386 10618 11388
rect 11605 11386 11671 11389
rect 10612 11384 11671 11386
rect 10612 11328 11610 11384
rect 11666 11328 11671 11384
rect 10612 11326 11671 11328
rect 10612 11324 10618 11326
rect 11605 11323 11671 11326
rect 12433 11250 12499 11253
rect 12985 11250 13051 11253
rect 9630 11248 12499 11250
rect 9630 11192 12438 11248
rect 12494 11192 12499 11248
rect 9630 11190 12499 11192
rect 12433 11187 12499 11190
rect 12758 11248 13051 11250
rect 12758 11192 12990 11248
rect 13046 11192 13051 11248
rect 12758 11190 13051 11192
rect 606 11052 612 11116
rect 676 11114 682 11116
rect 3417 11114 3483 11117
rect 676 11112 3483 11114
rect 676 11056 3422 11112
rect 3478 11056 3483 11112
rect 676 11054 3483 11056
rect 676 11052 682 11054
rect 3417 11051 3483 11054
rect 3601 11114 3667 11117
rect 10225 11114 10291 11117
rect 12758 11114 12818 11190
rect 12985 11187 13051 11190
rect 3601 11112 10291 11114
rect 3601 11056 3606 11112
rect 3662 11056 10230 11112
rect 10286 11056 10291 11112
rect 3601 11054 10291 11056
rect 3601 11051 3667 11054
rect 10225 11051 10291 11054
rect 12390 11054 12818 11114
rect 2998 10916 3004 10980
rect 3068 10978 3074 10980
rect 4245 10978 4311 10981
rect 3068 10976 4311 10978
rect 3068 10920 4250 10976
rect 4306 10920 4311 10976
rect 3068 10918 4311 10920
rect 3068 10916 3074 10918
rect 4245 10915 4311 10918
rect 5165 10980 5231 10981
rect 5165 10976 5212 10980
rect 5276 10978 5282 10980
rect 5533 10978 5599 10981
rect 7189 10978 7255 10981
rect 5165 10920 5170 10976
rect 5165 10916 5212 10920
rect 5276 10918 5322 10978
rect 5533 10976 7255 10978
rect 5533 10920 5538 10976
rect 5594 10920 7194 10976
rect 7250 10920 7255 10976
rect 5533 10918 7255 10920
rect 5276 10916 5282 10918
rect 5165 10915 5231 10916
rect 5533 10915 5599 10918
rect 7189 10915 7255 10918
rect 9622 10916 9628 10980
rect 9692 10978 9698 10980
rect 12390 10978 12450 11054
rect 9692 10918 12450 10978
rect 14457 10978 14523 10981
rect 15200 10978 16000 11008
rect 14457 10976 16000 10978
rect 14457 10920 14462 10976
rect 14518 10920 16000 10976
rect 14457 10918 16000 10920
rect 9692 10916 9698 10918
rect 14457 10915 14523 10918
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 15200 10888 16000 10918
rect 12606 10847 12922 10848
rect 3734 10780 3740 10844
rect 3804 10842 3810 10844
rect 7005 10842 7071 10845
rect 7373 10844 7439 10845
rect 7373 10842 7420 10844
rect 3804 10840 7071 10842
rect 3804 10784 7010 10840
rect 7066 10784 7071 10840
rect 3804 10782 7071 10784
rect 7328 10840 7420 10842
rect 7328 10784 7378 10840
rect 7328 10782 7420 10784
rect 3804 10780 3810 10782
rect 7005 10779 7071 10782
rect 7373 10780 7420 10782
rect 7484 10780 7490 10844
rect 11646 10780 11652 10844
rect 11716 10842 11722 10844
rect 12341 10842 12407 10845
rect 11716 10840 12407 10842
rect 11716 10784 12346 10840
rect 12402 10784 12407 10840
rect 11716 10782 12407 10784
rect 11716 10780 11722 10782
rect 7373 10779 7439 10780
rect 12341 10779 12407 10782
rect 1669 10706 1735 10709
rect 2405 10706 2471 10709
rect 1669 10704 2471 10706
rect 1669 10648 1674 10704
rect 1730 10648 2410 10704
rect 2466 10648 2471 10704
rect 1669 10646 2471 10648
rect 1669 10643 1735 10646
rect 2405 10643 2471 10646
rect 6126 10644 6132 10708
rect 6196 10706 6202 10708
rect 6361 10706 6427 10709
rect 6196 10704 6427 10706
rect 6196 10648 6366 10704
rect 6422 10648 6427 10704
rect 6196 10646 6427 10648
rect 6196 10644 6202 10646
rect 6361 10643 6427 10646
rect 6637 10706 6703 10709
rect 10041 10706 10107 10709
rect 6637 10704 10107 10706
rect 6637 10648 6642 10704
rect 6698 10648 10046 10704
rect 10102 10648 10107 10704
rect 6637 10646 10107 10648
rect 6637 10643 6703 10646
rect 10041 10643 10107 10646
rect 10869 10706 10935 10709
rect 12709 10706 12775 10709
rect 10869 10704 12775 10706
rect 10869 10648 10874 10704
rect 10930 10648 12714 10704
rect 12770 10648 12775 10704
rect 10869 10646 12775 10648
rect 10869 10643 10935 10646
rect 12709 10643 12775 10646
rect 12525 10570 12591 10573
rect 2730 10568 12591 10570
rect 2730 10512 12530 10568
rect 12586 10512 12591 10568
rect 2730 10510 12591 10512
rect 2405 10434 2471 10437
rect 2730 10434 2790 10510
rect 12525 10507 12591 10510
rect 2405 10432 2790 10434
rect 2405 10376 2410 10432
rect 2466 10376 2790 10432
rect 2405 10374 2790 10376
rect 4705 10434 4771 10437
rect 4838 10434 4844 10436
rect 4705 10432 4844 10434
rect 4705 10376 4710 10432
rect 4766 10376 4844 10432
rect 4705 10374 4844 10376
rect 2405 10371 2471 10374
rect 4705 10371 4771 10374
rect 4838 10372 4844 10374
rect 4908 10372 4914 10436
rect 5073 10434 5139 10437
rect 6729 10434 6795 10437
rect 5073 10432 6795 10434
rect 5073 10376 5078 10432
rect 5134 10376 6734 10432
rect 6790 10376 6795 10432
rect 5073 10374 6795 10376
rect 5073 10371 5139 10374
rect 6729 10371 6795 10374
rect 7373 10436 7439 10437
rect 7373 10432 7420 10436
rect 7484 10434 7490 10436
rect 7373 10376 7378 10432
rect 7373 10372 7420 10376
rect 7484 10374 7530 10434
rect 7484 10372 7490 10374
rect 7373 10371 7439 10372
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 6085 10298 6151 10301
rect 6729 10298 6795 10301
rect 6085 10296 6795 10298
rect 6085 10240 6090 10296
rect 6146 10240 6734 10296
rect 6790 10240 6795 10296
rect 6085 10238 6795 10240
rect 6085 10235 6151 10238
rect 6729 10235 6795 10238
rect 7414 10236 7420 10300
rect 7484 10298 7490 10300
rect 11053 10298 11119 10301
rect 7484 10296 11119 10298
rect 7484 10240 11058 10296
rect 11114 10240 11119 10296
rect 7484 10238 11119 10240
rect 7484 10236 7490 10238
rect 11053 10235 11119 10238
rect 2957 10162 3023 10165
rect 6269 10162 6335 10165
rect 2957 10160 6335 10162
rect 2957 10104 2962 10160
rect 3018 10104 6274 10160
rect 6330 10104 6335 10160
rect 2957 10102 6335 10104
rect 2957 10099 3023 10102
rect 6269 10099 6335 10102
rect 6453 10162 6519 10165
rect 8293 10162 8359 10165
rect 6453 10160 8359 10162
rect 6453 10104 6458 10160
rect 6514 10104 8298 10160
rect 8354 10104 8359 10160
rect 6453 10102 8359 10104
rect 6453 10099 6519 10102
rect 8293 10099 8359 10102
rect 11053 10162 11119 10165
rect 12985 10162 13051 10165
rect 11053 10160 13051 10162
rect 11053 10104 11058 10160
rect 11114 10104 12990 10160
rect 13046 10104 13051 10160
rect 11053 10102 13051 10104
rect 11053 10099 11119 10102
rect 12985 10099 13051 10102
rect 13445 10160 13511 10165
rect 13445 10104 13450 10160
rect 13506 10104 13511 10160
rect 13445 10099 13511 10104
rect 749 10026 815 10029
rect 6637 10026 6703 10029
rect 749 10024 6703 10026
rect 749 9968 754 10024
rect 810 9968 6642 10024
rect 6698 9968 6703 10024
rect 749 9966 6703 9968
rect 749 9963 815 9966
rect 6637 9963 6703 9966
rect 6913 10026 6979 10029
rect 9121 10026 9187 10029
rect 6913 10024 9187 10026
rect 6913 9968 6918 10024
rect 6974 9968 9126 10024
rect 9182 9968 9187 10024
rect 6913 9966 9187 9968
rect 6913 9963 6979 9966
rect 9121 9963 9187 9966
rect 11237 10026 11303 10029
rect 13448 10026 13508 10099
rect 11237 10024 13508 10026
rect 11237 9968 11242 10024
rect 11298 9968 13508 10024
rect 11237 9966 13508 9968
rect 11237 9963 11303 9966
rect 5441 9890 5507 9893
rect 7414 9890 7420 9892
rect 5441 9888 7420 9890
rect 5441 9832 5446 9888
rect 5502 9832 7420 9888
rect 5441 9830 7420 9832
rect 5441 9827 5507 9830
rect 7414 9828 7420 9830
rect 7484 9828 7490 9892
rect 13997 9890 14063 9893
rect 14457 9890 14523 9893
rect 15200 9890 16000 9920
rect 13997 9888 14106 9890
rect 13997 9832 14002 9888
rect 14058 9832 14106 9888
rect 13997 9827 14106 9832
rect 14457 9888 16000 9890
rect 14457 9832 14462 9888
rect 14518 9832 16000 9888
rect 14457 9830 16000 9832
rect 14457 9827 14523 9830
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 4521 9754 4587 9757
rect 4654 9754 4660 9756
rect 4521 9752 4660 9754
rect 4521 9696 4526 9752
rect 4582 9696 4660 9752
rect 4521 9694 4660 9696
rect 4521 9691 4587 9694
rect 4654 9692 4660 9694
rect 4724 9692 4730 9756
rect 9857 9754 9923 9757
rect 11462 9754 11468 9756
rect 9857 9752 11468 9754
rect 9857 9696 9862 9752
rect 9918 9696 11468 9752
rect 9857 9694 11468 9696
rect 9857 9691 9923 9694
rect 11462 9692 11468 9694
rect 11532 9692 11538 9756
rect 1301 9618 1367 9621
rect 6502 9618 7252 9652
rect 10317 9618 10383 9621
rect 1301 9616 10383 9618
rect 1301 9560 1306 9616
rect 1362 9592 10322 9616
rect 1362 9560 6562 9592
rect 1301 9558 6562 9560
rect 7192 9560 10322 9592
rect 10378 9560 10383 9616
rect 7192 9558 10383 9560
rect 1301 9555 1367 9558
rect 10317 9555 10383 9558
rect 13261 9616 13327 9621
rect 13261 9560 13266 9616
rect 13322 9560 13327 9616
rect 13261 9555 13327 9560
rect 4153 9482 4219 9485
rect 6640 9482 7068 9516
rect 9622 9482 9628 9484
rect 4153 9480 9628 9482
rect 4153 9424 4158 9480
rect 4214 9456 9628 9480
rect 4214 9424 6700 9456
rect 4153 9422 6700 9424
rect 7008 9422 9628 9456
rect 4153 9419 4219 9422
rect 9622 9420 9628 9422
rect 9692 9420 9698 9484
rect 11881 9482 11947 9485
rect 12433 9484 12499 9485
rect 11700 9480 11947 9482
rect 11700 9424 11886 9480
rect 11942 9424 11947 9480
rect 11700 9422 11947 9424
rect 4429 9346 4495 9349
rect 4797 9346 4863 9349
rect 4429 9344 4863 9346
rect 4429 9288 4434 9344
rect 4490 9288 4802 9344
rect 4858 9288 4863 9344
rect 4429 9286 4863 9288
rect 4429 9283 4495 9286
rect 4797 9283 4863 9286
rect 5942 9284 5948 9348
rect 6012 9346 6018 9348
rect 6085 9346 6151 9349
rect 6012 9344 6151 9346
rect 6012 9288 6090 9344
rect 6146 9288 6151 9344
rect 6012 9286 6151 9288
rect 6012 9284 6018 9286
rect 6085 9283 6151 9286
rect 6361 9346 6427 9349
rect 6494 9346 6500 9348
rect 6361 9344 6500 9346
rect 6361 9288 6366 9344
rect 6422 9288 6500 9344
rect 6361 9286 6500 9288
rect 6361 9283 6427 9286
rect 6494 9284 6500 9286
rect 6564 9346 6570 9348
rect 6729 9346 6795 9349
rect 6564 9344 6795 9346
rect 6564 9288 6734 9344
rect 6790 9288 6795 9344
rect 6564 9286 6795 9288
rect 6564 9284 6570 9286
rect 6729 9283 6795 9286
rect 9029 9348 9095 9349
rect 9029 9344 9076 9348
rect 9140 9346 9146 9348
rect 9029 9288 9034 9344
rect 9029 9284 9076 9288
rect 9140 9286 9186 9346
rect 9140 9284 9146 9286
rect 9622 9284 9628 9348
rect 9692 9346 9698 9348
rect 10133 9346 10199 9349
rect 9692 9344 10199 9346
rect 9692 9288 10138 9344
rect 10194 9288 10199 9344
rect 9692 9286 10199 9288
rect 9692 9284 9698 9286
rect 9029 9283 9095 9284
rect 10133 9283 10199 9286
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 2865 9210 2931 9213
rect 6729 9210 6795 9213
rect 2865 9208 6795 9210
rect 2865 9152 2870 9208
rect 2926 9152 6734 9208
rect 6790 9152 6795 9208
rect 2865 9150 6795 9152
rect 2865 9147 2931 9150
rect 6729 9147 6795 9150
rect 7465 9210 7531 9213
rect 9673 9210 9739 9213
rect 9857 9210 9923 9213
rect 7465 9208 9923 9210
rect 7465 9152 7470 9208
rect 7526 9152 9678 9208
rect 9734 9152 9862 9208
rect 9918 9152 9923 9208
rect 7465 9150 9923 9152
rect 7465 9147 7531 9150
rect 9673 9147 9739 9150
rect 9857 9147 9923 9150
rect 4429 9074 4495 9077
rect 9673 9074 9739 9077
rect 4429 9072 9739 9074
rect 4429 9016 4434 9072
rect 4490 9016 9678 9072
rect 9734 9016 9739 9072
rect 4429 9014 9739 9016
rect 4429 9011 4495 9014
rect 9673 9011 9739 9014
rect 11053 9076 11119 9077
rect 11053 9072 11100 9076
rect 11164 9074 11170 9076
rect 11700 9074 11760 9422
rect 11881 9419 11947 9422
rect 12382 9420 12388 9484
rect 12452 9482 12499 9484
rect 13264 9482 13324 9555
rect 12452 9480 13324 9482
rect 12494 9424 13324 9480
rect 12452 9422 13324 9424
rect 14046 9482 14106 9827
rect 15200 9800 16000 9830
rect 14273 9482 14339 9485
rect 14046 9480 14339 9482
rect 14046 9424 14278 9480
rect 14334 9424 14339 9480
rect 14046 9422 14339 9424
rect 12452 9420 12499 9422
rect 12433 9419 12499 9420
rect 14273 9419 14339 9422
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 11881 9074 11947 9077
rect 11053 9016 11058 9072
rect 11053 9012 11100 9016
rect 11164 9014 11210 9074
rect 11700 9072 11947 9074
rect 11700 9016 11886 9072
rect 11942 9016 11947 9072
rect 11700 9014 11947 9016
rect 11164 9012 11170 9014
rect 11053 9011 11119 9012
rect 11881 9011 11947 9014
rect 6177 8938 6243 8941
rect 6913 8938 6979 8941
rect 6177 8936 6979 8938
rect 6177 8880 6182 8936
rect 6238 8880 6918 8936
rect 6974 8880 6979 8936
rect 6177 8878 6979 8880
rect 6177 8875 6243 8878
rect 6913 8875 6979 8878
rect 7422 8878 8218 8938
rect 3049 8802 3115 8805
rect 7422 8802 7482 8878
rect 3049 8800 7482 8802
rect 3049 8744 3054 8800
rect 3110 8744 7482 8800
rect 3049 8742 7482 8744
rect 8158 8802 8218 8878
rect 8334 8876 8340 8940
rect 8404 8938 8410 8940
rect 10685 8938 10751 8941
rect 8404 8936 10751 8938
rect 8404 8880 10690 8936
rect 10746 8880 10751 8936
rect 8404 8878 10751 8880
rect 8404 8876 8410 8878
rect 10685 8875 10751 8878
rect 10869 8940 10935 8941
rect 10869 8936 10916 8940
rect 10980 8938 10986 8940
rect 11513 8938 11579 8941
rect 10980 8936 11579 8938
rect 10869 8880 10874 8936
rect 10980 8880 11518 8936
rect 11574 8880 11579 8936
rect 10869 8876 10916 8880
rect 10980 8878 11579 8880
rect 10980 8876 10986 8878
rect 10869 8875 10935 8876
rect 11513 8875 11579 8878
rect 9622 8802 9628 8804
rect 8158 8742 9628 8802
rect 3049 8739 3115 8742
rect 9622 8740 9628 8742
rect 9692 8740 9698 8804
rect 9857 8802 9923 8805
rect 11973 8802 12039 8805
rect 9857 8800 12039 8802
rect 9857 8744 9862 8800
rect 9918 8744 11978 8800
rect 12034 8744 12039 8800
rect 9857 8742 12039 8744
rect 9857 8739 9923 8742
rect 11973 8739 12039 8742
rect 14457 8802 14523 8805
rect 15200 8802 16000 8832
rect 14457 8800 16000 8802
rect 14457 8744 14462 8800
rect 14518 8744 16000 8800
rect 14457 8742 16000 8744
rect 14457 8739 14523 8742
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 15200 8712 16000 8742
rect 12606 8671 12922 8672
rect 3785 8666 3851 8669
rect 4981 8668 5047 8669
rect 4470 8666 4476 8668
rect 3785 8664 4476 8666
rect 3785 8608 3790 8664
rect 3846 8608 4476 8664
rect 3785 8606 4476 8608
rect 3785 8603 3851 8606
rect 4470 8604 4476 8606
rect 4540 8604 4546 8668
rect 4981 8666 5028 8668
rect 4936 8664 5028 8666
rect 4936 8608 4986 8664
rect 4936 8606 5028 8608
rect 4981 8604 5028 8606
rect 5092 8604 5098 8668
rect 5206 8604 5212 8668
rect 5276 8666 5282 8668
rect 5441 8666 5507 8669
rect 5276 8664 5507 8666
rect 5276 8608 5446 8664
rect 5502 8608 5507 8664
rect 5276 8606 5507 8608
rect 5276 8604 5282 8606
rect 4981 8603 5047 8604
rect 5441 8603 5507 8606
rect 5625 8666 5691 8669
rect 8201 8668 8267 8669
rect 10409 8668 10475 8669
rect 5758 8666 5764 8668
rect 5625 8664 5764 8666
rect 5625 8608 5630 8664
rect 5686 8608 5764 8664
rect 5625 8606 5764 8608
rect 5625 8603 5691 8606
rect 5758 8604 5764 8606
rect 5828 8604 5834 8668
rect 8150 8666 8156 8668
rect 8110 8606 8156 8666
rect 8220 8664 8267 8668
rect 8262 8608 8267 8664
rect 8150 8604 8156 8606
rect 8220 8604 8267 8608
rect 10358 8604 10364 8668
rect 10428 8666 10475 8668
rect 10428 8664 10520 8666
rect 10470 8608 10520 8664
rect 10428 8606 10520 8608
rect 10428 8604 10475 8606
rect 11278 8604 11284 8668
rect 11348 8666 11354 8668
rect 11513 8666 11579 8669
rect 11348 8664 11579 8666
rect 11348 8608 11518 8664
rect 11574 8608 11579 8664
rect 11348 8606 11579 8608
rect 11348 8604 11354 8606
rect 8201 8603 8267 8604
rect 10409 8603 10475 8604
rect 11513 8603 11579 8606
rect 10133 8530 10199 8533
rect 2730 8528 10199 8530
rect 2730 8472 10138 8528
rect 10194 8472 10199 8528
rect 2730 8470 10199 8472
rect 1853 8394 1919 8397
rect 2730 8394 2790 8470
rect 10133 8467 10199 8470
rect 1853 8392 2790 8394
rect 1853 8336 1858 8392
rect 1914 8336 2790 8392
rect 1853 8334 2790 8336
rect 3049 8394 3115 8397
rect 4153 8394 4219 8397
rect 3049 8392 4219 8394
rect 3049 8336 3054 8392
rect 3110 8336 4158 8392
rect 4214 8336 4219 8392
rect 3049 8334 4219 8336
rect 1853 8331 1919 8334
rect 3049 8331 3115 8334
rect 4153 8331 4219 8334
rect 4286 8332 4292 8396
rect 4356 8394 4362 8396
rect 8661 8394 8727 8397
rect 4356 8392 8727 8394
rect 4356 8336 8666 8392
rect 8722 8336 8727 8392
rect 4356 8334 8727 8336
rect 4356 8332 4362 8334
rect 8661 8331 8727 8334
rect 9121 8394 9187 8397
rect 14089 8394 14155 8397
rect 9121 8392 14155 8394
rect 9121 8336 9126 8392
rect 9182 8336 14094 8392
rect 14150 8336 14155 8392
rect 9121 8334 14155 8336
rect 9121 8331 9187 8334
rect 14089 8331 14155 8334
rect 3325 8258 3391 8261
rect 2730 8256 3391 8258
rect 2730 8200 3330 8256
rect 3386 8200 3391 8256
rect 2730 8198 3391 8200
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 2405 8122 2471 8125
rect 2730 8122 2790 8198
rect 3325 8195 3391 8198
rect 3969 8258 4035 8261
rect 5574 8258 5580 8260
rect 3969 8256 5580 8258
rect 3969 8200 3974 8256
rect 4030 8200 5580 8256
rect 3969 8198 5580 8200
rect 3969 8195 4035 8198
rect 5574 8196 5580 8198
rect 5644 8196 5650 8260
rect 7925 8258 7991 8261
rect 8518 8258 8524 8260
rect 7925 8256 8524 8258
rect 7925 8200 7930 8256
rect 7986 8200 8524 8256
rect 7925 8198 8524 8200
rect 7925 8195 7991 8198
rect 8518 8196 8524 8198
rect 8588 8196 8594 8260
rect 9765 8258 9831 8261
rect 10174 8258 10180 8260
rect 9765 8256 10180 8258
rect 9765 8200 9770 8256
rect 9826 8200 10180 8256
rect 9765 8198 10180 8200
rect 9765 8195 9831 8198
rect 10174 8196 10180 8198
rect 10244 8196 10250 8260
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 2405 8120 2790 8122
rect 2405 8064 2410 8120
rect 2466 8064 2790 8120
rect 2405 8062 2790 8064
rect 2405 8059 2471 8062
rect 7414 8060 7420 8124
rect 7484 8122 7490 8124
rect 10685 8122 10751 8125
rect 7484 8120 10751 8122
rect 7484 8064 10690 8120
rect 10746 8064 10751 8120
rect 7484 8062 10751 8064
rect 7484 8060 7490 8062
rect 10685 8059 10751 8062
rect 3417 7986 3483 7989
rect 4981 7986 5047 7989
rect 3417 7984 5047 7986
rect 3417 7928 3422 7984
rect 3478 7928 4986 7984
rect 5042 7928 5047 7984
rect 3417 7926 5047 7928
rect 3417 7923 3483 7926
rect 4981 7923 5047 7926
rect 5901 7986 5967 7989
rect 9806 7986 9812 7988
rect 5901 7984 9812 7986
rect 5901 7928 5906 7984
rect 5962 7928 9812 7984
rect 5901 7926 9812 7928
rect 5901 7923 5967 7926
rect 9806 7924 9812 7926
rect 9876 7924 9882 7988
rect 5390 7788 5396 7852
rect 5460 7850 5466 7852
rect 9121 7850 9187 7853
rect 5460 7848 9187 7850
rect 5460 7792 9126 7848
rect 9182 7792 9187 7848
rect 5460 7790 9187 7792
rect 5460 7788 5466 7790
rect 9121 7787 9187 7790
rect 4429 7714 4495 7717
rect 6177 7714 6243 7717
rect 7414 7714 7420 7716
rect 4429 7712 6056 7714
rect 4429 7656 4434 7712
rect 4490 7656 6056 7712
rect 4429 7654 6056 7656
rect 4429 7651 4495 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 4838 7516 4844 7580
rect 4908 7578 4914 7580
rect 4981 7578 5047 7581
rect 4908 7576 5047 7578
rect 4908 7520 4986 7576
rect 5042 7520 5047 7576
rect 4908 7518 5047 7520
rect 5996 7578 6056 7654
rect 6177 7712 7420 7714
rect 6177 7656 6182 7712
rect 6238 7656 7420 7712
rect 6177 7654 7420 7656
rect 6177 7651 6243 7654
rect 7414 7652 7420 7654
rect 7484 7652 7490 7716
rect 14457 7714 14523 7717
rect 15200 7714 16000 7744
rect 14457 7712 16000 7714
rect 14457 7656 14462 7712
rect 14518 7656 16000 7712
rect 14457 7654 16000 7656
rect 14457 7651 14523 7654
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 15200 7624 16000 7654
rect 12606 7583 12922 7584
rect 7414 7578 7420 7580
rect 5996 7518 7420 7578
rect 4908 7516 4914 7518
rect 4981 7515 5047 7518
rect 7414 7516 7420 7518
rect 7484 7516 7490 7580
rect 14038 7516 14044 7580
rect 14108 7578 14114 7580
rect 14181 7578 14247 7581
rect 14108 7576 14247 7578
rect 14108 7520 14186 7576
rect 14242 7520 14247 7576
rect 14108 7518 14247 7520
rect 14108 7516 14114 7518
rect 14181 7515 14247 7518
rect 1761 7442 1827 7445
rect 8150 7442 8156 7444
rect 1761 7440 8156 7442
rect 1761 7384 1766 7440
rect 1822 7384 8156 7440
rect 1761 7382 8156 7384
rect 1761 7379 1827 7382
rect 8150 7380 8156 7382
rect 8220 7380 8226 7444
rect 10041 7442 10107 7445
rect 12709 7442 12775 7445
rect 10041 7440 12775 7442
rect 10041 7384 10046 7440
rect 10102 7384 12714 7440
rect 12770 7384 12775 7440
rect 10041 7382 12775 7384
rect 10041 7379 10107 7382
rect 12709 7379 12775 7382
rect 12893 7442 12959 7445
rect 13118 7442 13124 7444
rect 12893 7440 13124 7442
rect 12893 7384 12898 7440
rect 12954 7384 13124 7440
rect 12893 7382 13124 7384
rect 12893 7379 12959 7382
rect 13118 7380 13124 7382
rect 13188 7380 13194 7444
rect 1853 7306 1919 7309
rect 2313 7306 2379 7309
rect 5758 7306 5764 7308
rect 1853 7304 5764 7306
rect 1853 7248 1858 7304
rect 1914 7248 2318 7304
rect 2374 7248 5764 7304
rect 1853 7246 5764 7248
rect 1853 7243 1919 7246
rect 2313 7243 2379 7246
rect 5758 7244 5764 7246
rect 5828 7244 5834 7308
rect 5901 7306 5967 7309
rect 6126 7306 6132 7308
rect 5901 7304 6132 7306
rect 5901 7248 5906 7304
rect 5962 7248 6132 7304
rect 5901 7246 6132 7248
rect 5901 7243 5967 7246
rect 6126 7244 6132 7246
rect 6196 7244 6202 7308
rect 6729 7306 6795 7309
rect 14733 7306 14799 7309
rect 6729 7304 14799 7306
rect 6729 7248 6734 7304
rect 6790 7248 14738 7304
rect 14794 7248 14799 7304
rect 6729 7246 14799 7248
rect 6729 7243 6795 7246
rect 14733 7243 14799 7246
rect 4102 7108 4108 7172
rect 4172 7170 4178 7172
rect 6729 7170 6795 7173
rect 4172 7168 6795 7170
rect 4172 7112 6734 7168
rect 6790 7112 6795 7168
rect 4172 7110 6795 7112
rect 4172 7108 4178 7110
rect 6729 7107 6795 7110
rect 8886 7108 8892 7172
rect 8956 7170 8962 7172
rect 9581 7170 9647 7173
rect 8956 7168 9647 7170
rect 8956 7112 9586 7168
rect 9642 7112 9647 7168
rect 8956 7110 9647 7112
rect 8956 7108 8962 7110
rect 9581 7107 9647 7110
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 2446 6972 2452 7036
rect 2516 7034 2522 7036
rect 6269 7034 6335 7037
rect 2516 7032 6335 7034
rect 2516 6976 6274 7032
rect 6330 6976 6335 7032
rect 2516 6974 6335 6976
rect 2516 6972 2522 6974
rect 6269 6971 6335 6974
rect 7414 6972 7420 7036
rect 7484 7034 7490 7036
rect 8477 7034 8543 7037
rect 9990 7034 9996 7036
rect 7484 7032 9996 7034
rect 7484 6976 8482 7032
rect 8538 6976 9996 7032
rect 7484 6974 9996 6976
rect 7484 6972 7490 6974
rect 8477 6971 8543 6974
rect 9990 6972 9996 6974
rect 10060 6972 10066 7036
rect 10174 6972 10180 7036
rect 10244 7034 10250 7036
rect 11421 7034 11487 7037
rect 10244 7032 11487 7034
rect 10244 6976 11426 7032
rect 11482 6976 11487 7032
rect 10244 6974 11487 6976
rect 10244 6972 10250 6974
rect 11421 6971 11487 6974
rect 13854 6972 13860 7036
rect 13924 7034 13930 7036
rect 14365 7034 14431 7037
rect 13924 7032 14431 7034
rect 13924 6976 14370 7032
rect 14426 6976 14431 7032
rect 13924 6974 14431 6976
rect 13924 6972 13930 6974
rect 14365 6971 14431 6974
rect 974 6836 980 6900
rect 1044 6898 1050 6900
rect 3049 6898 3115 6901
rect 1044 6896 3115 6898
rect 1044 6840 3054 6896
rect 3110 6840 3115 6896
rect 1044 6838 3115 6840
rect 1044 6836 1050 6838
rect 3049 6835 3115 6838
rect 4981 6898 5047 6901
rect 8334 6898 8340 6900
rect 4981 6896 8340 6898
rect 4981 6840 4986 6896
rect 5042 6840 8340 6896
rect 4981 6838 8340 6840
rect 4981 6835 5047 6838
rect 8334 6836 8340 6838
rect 8404 6836 8410 6900
rect 9121 6898 9187 6901
rect 9254 6898 9260 6900
rect 9121 6896 9260 6898
rect 9121 6840 9126 6896
rect 9182 6840 9260 6896
rect 9121 6838 9260 6840
rect 9121 6835 9187 6838
rect 9254 6836 9260 6838
rect 9324 6836 9330 6900
rect 9581 6898 9647 6901
rect 11094 6898 11100 6900
rect 9581 6896 11100 6898
rect 9581 6840 9586 6896
rect 9642 6840 11100 6896
rect 9581 6838 11100 6840
rect 9581 6835 9647 6838
rect 11094 6836 11100 6838
rect 11164 6898 11170 6900
rect 11605 6898 11671 6901
rect 11164 6896 11671 6898
rect 11164 6840 11610 6896
rect 11666 6840 11671 6896
rect 11164 6838 11671 6840
rect 11164 6836 11170 6838
rect 11605 6835 11671 6838
rect 13302 6836 13308 6900
rect 13372 6898 13378 6900
rect 13629 6898 13695 6901
rect 13372 6896 13695 6898
rect 13372 6840 13634 6896
rect 13690 6840 13695 6896
rect 13372 6838 13695 6840
rect 13372 6836 13378 6838
rect 13629 6835 13695 6838
rect 2773 6762 2839 6765
rect 5625 6762 5691 6765
rect 13353 6762 13419 6765
rect 2773 6760 5691 6762
rect 2773 6704 2778 6760
rect 2834 6704 5630 6760
rect 5686 6704 5691 6760
rect 2773 6702 5691 6704
rect 2773 6699 2839 6702
rect 5625 6699 5691 6702
rect 5766 6760 13419 6762
rect 5766 6704 13358 6760
rect 13414 6704 13419 6760
rect 5766 6702 13419 6704
rect 3601 6626 3667 6629
rect 5766 6626 5826 6702
rect 13353 6699 13419 6702
rect 3601 6624 5826 6626
rect 3601 6568 3606 6624
rect 3662 6568 5826 6624
rect 3601 6566 5826 6568
rect 3601 6563 3667 6566
rect 5942 6564 5948 6628
rect 6012 6626 6018 6628
rect 6821 6626 6887 6629
rect 6012 6624 6887 6626
rect 6012 6568 6826 6624
rect 6882 6568 6887 6624
rect 6012 6566 6887 6568
rect 6012 6564 6018 6566
rect 6821 6563 6887 6566
rect 8937 6626 9003 6629
rect 11278 6626 11284 6628
rect 8937 6624 11284 6626
rect 8937 6568 8942 6624
rect 8998 6568 11284 6624
rect 8937 6566 11284 6568
rect 8937 6563 9003 6566
rect 11278 6564 11284 6566
rect 11348 6564 11354 6628
rect 14181 6626 14247 6629
rect 15200 6626 16000 6656
rect 14181 6624 16000 6626
rect 14181 6568 14186 6624
rect 14242 6568 16000 6624
rect 14181 6566 16000 6568
rect 14181 6563 14247 6566
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 15200 6536 16000 6566
rect 12606 6495 12922 6496
rect 3325 6490 3391 6493
rect 4470 6490 4476 6492
rect 3325 6488 4476 6490
rect 3325 6432 3330 6488
rect 3386 6432 4476 6488
rect 3325 6430 4476 6432
rect 3325 6427 3391 6430
rect 4470 6428 4476 6430
rect 4540 6490 4546 6492
rect 4540 6430 4722 6490
rect 4540 6428 4546 6430
rect 790 6292 796 6356
rect 860 6354 866 6356
rect 4429 6354 4495 6357
rect 860 6352 4495 6354
rect 860 6296 4434 6352
rect 4490 6296 4495 6352
rect 860 6294 4495 6296
rect 4662 6354 4722 6430
rect 6678 6428 6684 6492
rect 6748 6490 6754 6492
rect 7465 6490 7531 6493
rect 6748 6488 7531 6490
rect 6748 6432 7470 6488
rect 7526 6432 7531 6488
rect 6748 6430 7531 6432
rect 6748 6428 6754 6430
rect 7465 6427 7531 6430
rect 9121 6490 9187 6493
rect 11237 6490 11303 6493
rect 9121 6488 11303 6490
rect 9121 6432 9126 6488
rect 9182 6432 11242 6488
rect 11298 6432 11303 6488
rect 9121 6430 11303 6432
rect 9121 6427 9187 6430
rect 11237 6427 11303 6430
rect 10358 6354 10364 6356
rect 4662 6294 10364 6354
rect 860 6292 866 6294
rect 4429 6291 4495 6294
rect 10358 6292 10364 6294
rect 10428 6292 10434 6356
rect 3877 6218 3943 6221
rect 8845 6218 8911 6221
rect 3877 6216 8911 6218
rect 3877 6160 3882 6216
rect 3938 6160 8850 6216
rect 8906 6160 8911 6216
rect 3877 6158 8911 6160
rect 3877 6155 3943 6158
rect 8845 6155 8911 6158
rect 9673 6218 9739 6221
rect 11789 6218 11855 6221
rect 9673 6216 11855 6218
rect 9673 6160 9678 6216
rect 9734 6160 11794 6216
rect 11850 6160 11855 6216
rect 9673 6158 11855 6160
rect 9673 6155 9739 6158
rect 11789 6155 11855 6158
rect 7741 6082 7807 6085
rect 8661 6082 8727 6085
rect 7741 6080 8727 6082
rect 7741 6024 7746 6080
rect 7802 6024 8666 6080
rect 8722 6024 8727 6080
rect 7741 6022 8727 6024
rect 7741 6019 7807 6022
rect 8661 6019 8727 6022
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 3141 5946 3207 5949
rect 4286 5946 4292 5948
rect 3141 5944 4292 5946
rect 3141 5888 3146 5944
rect 3202 5888 4292 5944
rect 3141 5886 4292 5888
rect 3141 5883 3207 5886
rect 4286 5884 4292 5886
rect 4356 5884 4362 5948
rect 7373 5946 7439 5949
rect 8937 5946 9003 5949
rect 9070 5946 9076 5948
rect 7373 5944 9076 5946
rect 7373 5888 7378 5944
rect 7434 5888 8942 5944
rect 8998 5888 9076 5944
rect 7373 5886 9076 5888
rect 7373 5883 7439 5886
rect 8937 5883 9003 5886
rect 9070 5884 9076 5886
rect 9140 5884 9146 5948
rect 10358 5884 10364 5948
rect 10428 5946 10434 5948
rect 10428 5886 11714 5946
rect 10428 5884 10434 5886
rect 2957 5812 3023 5813
rect 2957 5810 3004 5812
rect 2912 5808 3004 5810
rect 2912 5752 2962 5808
rect 2912 5750 3004 5752
rect 2957 5748 3004 5750
rect 3068 5748 3074 5812
rect 4153 5810 4219 5813
rect 8385 5810 8451 5813
rect 11053 5810 11119 5813
rect 4153 5808 11119 5810
rect 4153 5752 4158 5808
rect 4214 5752 8390 5808
rect 8446 5752 11058 5808
rect 11114 5752 11119 5808
rect 4153 5750 11119 5752
rect 11654 5810 11714 5886
rect 11973 5810 12039 5813
rect 11654 5808 12039 5810
rect 11654 5752 11978 5808
rect 12034 5752 12039 5808
rect 11654 5750 12039 5752
rect 2957 5747 3023 5748
rect 4153 5747 4219 5750
rect 8385 5747 8451 5750
rect 11053 5747 11119 5750
rect 11973 5747 12039 5750
rect 3233 5674 3299 5677
rect 3550 5674 3556 5676
rect 3233 5672 3556 5674
rect 3233 5616 3238 5672
rect 3294 5616 3556 5672
rect 3233 5614 3556 5616
rect 3233 5611 3299 5614
rect 3550 5612 3556 5614
rect 3620 5612 3626 5676
rect 5441 5674 5507 5677
rect 11697 5674 11763 5677
rect 5441 5672 11763 5674
rect 5441 5616 5446 5672
rect 5502 5616 11702 5672
rect 11758 5616 11763 5672
rect 5441 5614 11763 5616
rect 5441 5611 5507 5614
rect 11697 5611 11763 5614
rect 3969 5538 4035 5541
rect 5993 5538 6059 5541
rect 3969 5536 6059 5538
rect 3969 5480 3974 5536
rect 4030 5480 5998 5536
rect 6054 5480 6059 5536
rect 3969 5478 6059 5480
rect 3969 5475 4035 5478
rect 5993 5475 6059 5478
rect 11789 5538 11855 5541
rect 12382 5538 12388 5540
rect 11789 5536 12388 5538
rect 11789 5480 11794 5536
rect 11850 5480 12388 5536
rect 11789 5478 12388 5480
rect 11789 5475 11855 5478
rect 12382 5476 12388 5478
rect 12452 5476 12458 5540
rect 14457 5538 14523 5541
rect 15200 5538 16000 5568
rect 14457 5536 16000 5538
rect 14457 5480 14462 5536
rect 14518 5480 16000 5536
rect 14457 5478 16000 5480
rect 14457 5475 14523 5478
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 15200 5448 16000 5478
rect 12606 5407 12922 5408
rect 8385 5402 8451 5405
rect 8886 5402 8892 5404
rect 8385 5400 8892 5402
rect 8385 5344 8390 5400
rect 8446 5344 8892 5400
rect 8385 5342 8892 5344
rect 8385 5339 8451 5342
rect 8886 5340 8892 5342
rect 8956 5340 8962 5404
rect 9489 5402 9555 5405
rect 9622 5402 9628 5404
rect 9489 5400 9628 5402
rect 9489 5344 9494 5400
rect 9550 5344 9628 5400
rect 9489 5342 9628 5344
rect 9489 5339 9555 5342
rect 9622 5340 9628 5342
rect 9692 5340 9698 5404
rect 9857 5402 9923 5405
rect 13445 5404 13511 5405
rect 10174 5402 10180 5404
rect 9857 5400 10180 5402
rect 9857 5344 9862 5400
rect 9918 5344 10180 5400
rect 9857 5342 10180 5344
rect 9857 5339 9923 5342
rect 10174 5340 10180 5342
rect 10244 5340 10250 5404
rect 13445 5402 13492 5404
rect 13364 5400 13492 5402
rect 13556 5402 13562 5404
rect 14273 5402 14339 5405
rect 13556 5400 14339 5402
rect 13364 5344 13450 5400
rect 13556 5344 14278 5400
rect 14334 5344 14339 5400
rect 13364 5342 13492 5344
rect 13445 5340 13492 5342
rect 13556 5342 14339 5344
rect 13556 5340 13562 5342
rect 13445 5339 13511 5340
rect 14273 5339 14339 5342
rect 3366 5204 3372 5268
rect 3436 5266 3442 5268
rect 3785 5266 3851 5269
rect 4521 5266 4587 5269
rect 3436 5264 4587 5266
rect 3436 5208 3790 5264
rect 3846 5208 4526 5264
rect 4582 5208 4587 5264
rect 3436 5206 4587 5208
rect 3436 5204 3442 5206
rect 3785 5203 3851 5206
rect 4521 5203 4587 5206
rect 6177 5266 6243 5269
rect 6310 5266 6316 5268
rect 6177 5264 6316 5266
rect 6177 5208 6182 5264
rect 6238 5208 6316 5264
rect 6177 5206 6316 5208
rect 6177 5203 6243 5206
rect 6310 5204 6316 5206
rect 6380 5204 6386 5268
rect 6453 5266 6519 5269
rect 7557 5266 7623 5269
rect 9397 5266 9463 5269
rect 6453 5264 9463 5266
rect 6453 5208 6458 5264
rect 6514 5208 7562 5264
rect 7618 5208 9402 5264
rect 9458 5208 9463 5264
rect 6453 5206 9463 5208
rect 6453 5203 6519 5206
rect 7557 5203 7623 5206
rect 9397 5203 9463 5206
rect 10869 5266 10935 5269
rect 11646 5266 11652 5268
rect 10869 5264 11652 5266
rect 10869 5208 10874 5264
rect 10930 5208 11652 5264
rect 10869 5206 11652 5208
rect 10869 5203 10935 5206
rect 11646 5204 11652 5206
rect 11716 5204 11722 5268
rect 3693 5130 3759 5133
rect 12893 5130 12959 5133
rect 3693 5128 12959 5130
rect 3693 5072 3698 5128
rect 3754 5072 12898 5128
rect 12954 5072 12959 5128
rect 3693 5070 12959 5072
rect 3693 5067 3759 5070
rect 12893 5067 12959 5070
rect 7925 4994 7991 4997
rect 8150 4994 8156 4996
rect 7925 4992 8156 4994
rect 7925 4936 7930 4992
rect 7986 4936 8156 4992
rect 7925 4934 8156 4936
rect 7925 4931 7991 4934
rect 8150 4932 8156 4934
rect 8220 4932 8226 4996
rect 8569 4994 8635 4997
rect 10409 4994 10475 4997
rect 8569 4992 10475 4994
rect 8569 4936 8574 4992
rect 8630 4936 10414 4992
rect 10470 4936 10475 4992
rect 8569 4934 10475 4936
rect 8569 4931 8635 4934
rect 10409 4931 10475 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 9438 4796 9444 4860
rect 9508 4858 9514 4860
rect 9581 4858 9647 4861
rect 9508 4856 9647 4858
rect 9508 4800 9586 4856
rect 9642 4800 9647 4856
rect 9508 4798 9647 4800
rect 9508 4796 9514 4798
rect 9581 4795 9647 4798
rect 5349 4722 5415 4725
rect 13905 4722 13971 4725
rect 5349 4720 13971 4722
rect 5349 4664 5354 4720
rect 5410 4664 13910 4720
rect 13966 4664 13971 4720
rect 5349 4662 13971 4664
rect 5349 4659 5415 4662
rect 13905 4659 13971 4662
rect 8201 4586 8267 4589
rect 14365 4586 14431 4589
rect 8201 4584 14431 4586
rect 8201 4528 8206 4584
rect 8262 4528 14370 4584
rect 14426 4528 14431 4584
rect 8201 4526 14431 4528
rect 8201 4523 8267 4526
rect 14365 4523 14431 4526
rect 0 4450 800 4480
rect 2446 4450 2452 4452
rect 0 4390 2452 4450
rect 0 4360 800 4390
rect 2446 4388 2452 4390
rect 2516 4388 2522 4452
rect 9070 4388 9076 4452
rect 9140 4450 9146 4452
rect 11053 4450 11119 4453
rect 9140 4448 11119 4450
rect 9140 4392 11058 4448
rect 11114 4392 11119 4448
rect 9140 4390 11119 4392
rect 9140 4388 9146 4390
rect 11053 4387 11119 4390
rect 13905 4450 13971 4453
rect 15200 4450 16000 4480
rect 13905 4448 16000 4450
rect 13905 4392 13910 4448
rect 13966 4392 16000 4448
rect 13905 4390 16000 4392
rect 13905 4387 13971 4390
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 15200 4360 16000 4390
rect 12606 4319 12922 4320
rect 9857 4314 9923 4317
rect 8158 4312 9923 4314
rect 8158 4256 9862 4312
rect 9918 4256 9923 4312
rect 8158 4254 9923 4256
rect 933 4178 999 4181
rect 8158 4178 8218 4254
rect 9857 4251 9923 4254
rect 10409 4314 10475 4317
rect 12157 4314 12223 4317
rect 10409 4312 12223 4314
rect 10409 4256 10414 4312
rect 10470 4256 12162 4312
rect 12218 4256 12223 4312
rect 10409 4254 12223 4256
rect 10409 4251 10475 4254
rect 12157 4251 12223 4254
rect 933 4176 8218 4178
rect 933 4120 938 4176
rect 994 4120 8218 4176
rect 933 4118 8218 4120
rect 11053 4178 11119 4181
rect 15009 4178 15075 4181
rect 11053 4176 15075 4178
rect 11053 4120 11058 4176
rect 11114 4120 15014 4176
rect 15070 4120 15075 4176
rect 11053 4118 15075 4120
rect 933 4115 999 4118
rect 11053 4115 11119 4118
rect 15009 4115 15075 4118
rect 7005 4042 7071 4045
rect 13077 4042 13143 4045
rect 2730 4040 13143 4042
rect 2730 3984 7010 4040
rect 7066 3984 13082 4040
rect 13138 3984 13143 4040
rect 2730 3982 13143 3984
rect 2405 3906 2471 3909
rect 2730 3906 2790 3982
rect 7005 3979 7071 3982
rect 13077 3979 13143 3982
rect 13445 4042 13511 4045
rect 14089 4042 14155 4045
rect 13445 4040 14155 4042
rect 13445 3984 13450 4040
rect 13506 3984 14094 4040
rect 14150 3984 14155 4040
rect 13445 3982 14155 3984
rect 13445 3979 13511 3982
rect 14089 3979 14155 3982
rect 2405 3904 2790 3906
rect 2405 3848 2410 3904
rect 2466 3848 2790 3904
rect 2405 3846 2790 3848
rect 2405 3843 2471 3846
rect 3918 3844 3924 3908
rect 3988 3906 3994 3908
rect 6545 3906 6611 3909
rect 3988 3904 6611 3906
rect 3988 3848 6550 3904
rect 6606 3848 6611 3904
rect 3988 3846 6611 3848
rect 3988 3844 3994 3846
rect 6545 3843 6611 3846
rect 8886 3844 8892 3908
rect 8956 3906 8962 3908
rect 9397 3906 9463 3909
rect 8956 3904 9463 3906
rect 8956 3848 9402 3904
rect 9458 3848 9463 3904
rect 8956 3846 9463 3848
rect 8956 3844 8962 3846
rect 9397 3843 9463 3846
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 3601 3634 3667 3637
rect 11605 3634 11671 3637
rect 14089 3634 14155 3637
rect 3601 3632 11671 3634
rect 3601 3576 3606 3632
rect 3662 3576 11610 3632
rect 11666 3576 11671 3632
rect 3601 3574 11671 3576
rect 3601 3571 3667 3574
rect 11605 3571 11671 3574
rect 12390 3632 14155 3634
rect 12390 3576 14094 3632
rect 14150 3576 14155 3632
rect 12390 3574 14155 3576
rect 1117 3498 1183 3501
rect 11513 3498 11579 3501
rect 1117 3496 11579 3498
rect 1117 3440 1122 3496
rect 1178 3440 11518 3496
rect 11574 3440 11579 3496
rect 1117 3438 11579 3440
rect 1117 3435 1183 3438
rect 11513 3435 11579 3438
rect 2998 3300 3004 3364
rect 3068 3362 3074 3364
rect 7465 3362 7531 3365
rect 3068 3360 7531 3362
rect 3068 3304 7470 3360
rect 7526 3304 7531 3360
rect 3068 3302 7531 3304
rect 3068 3300 3074 3302
rect 7465 3299 7531 3302
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 8518 3164 8524 3228
rect 8588 3226 8594 3228
rect 8661 3226 8727 3229
rect 12390 3226 12450 3574
rect 14089 3571 14155 3574
rect 13905 3362 13971 3365
rect 15200 3362 16000 3392
rect 13905 3360 16000 3362
rect 13905 3304 13910 3360
rect 13966 3304 16000 3360
rect 13905 3302 16000 3304
rect 13905 3299 13971 3302
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 15200 3272 16000 3302
rect 12606 3231 12922 3232
rect 8588 3224 8727 3226
rect 8588 3168 8666 3224
rect 8722 3168 8727 3224
rect 8588 3166 8727 3168
rect 8588 3164 8594 3166
rect 8661 3163 8727 3166
rect 10734 3166 12450 3226
rect 4889 3090 4955 3093
rect 10734 3090 10794 3166
rect 10961 3092 11027 3093
rect 4889 3088 10794 3090
rect 4889 3032 4894 3088
rect 4950 3032 10794 3088
rect 4889 3030 10794 3032
rect 4889 3027 4955 3030
rect 10910 3028 10916 3092
rect 10980 3090 11027 3092
rect 10980 3088 11072 3090
rect 11022 3032 11072 3088
rect 10980 3030 11072 3032
rect 10980 3028 11027 3030
rect 10961 3027 11027 3028
rect 6821 2954 6887 2957
rect 12525 2954 12591 2957
rect 6821 2952 12591 2954
rect 6821 2896 6826 2952
rect 6882 2896 12530 2952
rect 12586 2896 12591 2952
rect 6821 2894 12591 2896
rect 6821 2891 6887 2894
rect 12525 2891 12591 2894
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 11278 2620 11284 2684
rect 11348 2682 11354 2684
rect 11513 2682 11579 2685
rect 11348 2680 11579 2682
rect 11348 2624 11518 2680
rect 11574 2624 11579 2680
rect 11348 2622 11579 2624
rect 11348 2620 11354 2622
rect 11513 2619 11579 2622
rect 1526 2484 1532 2548
rect 1596 2546 1602 2548
rect 9070 2546 9076 2548
rect 1596 2486 9076 2546
rect 1596 2484 1602 2486
rect 9070 2484 9076 2486
rect 9140 2484 9146 2548
rect 9673 2546 9739 2549
rect 10869 2546 10935 2549
rect 9673 2544 10935 2546
rect 9673 2488 9678 2544
rect 9734 2488 10874 2544
rect 10930 2488 10935 2544
rect 9673 2486 10935 2488
rect 9673 2483 9739 2486
rect 10869 2483 10935 2486
rect 1710 2348 1716 2412
rect 1780 2410 1786 2412
rect 13261 2410 13327 2413
rect 1780 2408 13327 2410
rect 1780 2352 13266 2408
rect 13322 2352 13327 2408
rect 1780 2350 13327 2352
rect 1780 2348 1786 2350
rect 13261 2347 13327 2350
rect 13905 2274 13971 2277
rect 15200 2274 16000 2304
rect 13905 2272 16000 2274
rect 13905 2216 13910 2272
rect 13966 2216 16000 2272
rect 13905 2214 16000 2216
rect 13905 2211 13971 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 15200 2184 16000 2214
rect 12606 2143 12922 2144
rect 2497 2002 2563 2005
rect 11462 2002 11468 2004
rect 2497 2000 11468 2002
rect 2497 1944 2502 2000
rect 2558 1944 11468 2000
rect 2497 1942 11468 1944
rect 2497 1939 2563 1942
rect 11462 1940 11468 1942
rect 11532 1940 11538 2004
rect 1158 1804 1164 1868
rect 1228 1866 1234 1868
rect 11697 1866 11763 1869
rect 1228 1864 11763 1866
rect 1228 1808 11702 1864
rect 11758 1808 11763 1864
rect 1228 1806 11763 1808
rect 1228 1804 1234 1806
rect 11697 1803 11763 1806
rect 606 1668 612 1732
rect 676 1730 682 1732
rect 12985 1730 13051 1733
rect 676 1728 13051 1730
rect 676 1672 12990 1728
rect 13046 1672 13051 1728
rect 676 1670 13051 1672
rect 676 1668 682 1670
rect 12985 1667 13051 1670
rect 3734 1532 3740 1596
rect 3804 1594 3810 1596
rect 13813 1594 13879 1597
rect 3804 1592 13879 1594
rect 3804 1536 13818 1592
rect 13874 1536 13879 1592
rect 3804 1534 13879 1536
rect 3804 1532 3810 1534
rect 13813 1531 13879 1534
rect 13629 1186 13695 1189
rect 15200 1186 16000 1216
rect 13629 1184 16000 1186
rect 13629 1128 13634 1184
rect 13690 1128 16000 1184
rect 13629 1126 16000 1128
rect 13629 1123 13695 1126
rect 15200 1096 16000 1126
<< via3 >>
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 9260 15404 9324 15468
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 10548 14860 10612 14924
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 796 14316 860 14380
rect 11652 14180 11716 14244
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 12388 14044 12452 14108
rect 1164 13908 1228 13972
rect 4660 13908 4724 13972
rect 1716 13832 1780 13836
rect 1716 13776 1766 13832
rect 1766 13776 1780 13832
rect 1716 13772 1780 13776
rect 5396 13772 5460 13836
rect 5580 13832 5644 13836
rect 5580 13776 5630 13832
rect 5630 13776 5644 13832
rect 5580 13772 5644 13776
rect 6684 13772 6748 13836
rect 14044 13908 14108 13972
rect 13860 13772 13924 13836
rect 9812 13636 9876 13700
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 3924 13152 3988 13156
rect 3924 13096 3974 13152
rect 3974 13096 3988 13152
rect 3924 13092 3988 13096
rect 5948 13092 6012 13156
rect 8340 13092 8404 13156
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 3556 12956 3620 13020
rect 8524 12956 8588 13020
rect 980 12820 1044 12884
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 6316 12276 6380 12340
rect 12388 12276 12452 12340
rect 13124 12276 13188 12340
rect 6500 12140 6564 12204
rect 13492 12140 13556 12204
rect 5028 12004 5092 12068
rect 8156 12064 8220 12068
rect 8156 12008 8206 12064
rect 8206 12008 8220 12064
rect 8156 12004 8220 12008
rect 8524 12004 8588 12068
rect 11468 12004 11532 12068
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 8340 11928 8404 11932
rect 8340 11872 8354 11928
rect 8354 11872 8404 11928
rect 8340 11868 8404 11872
rect 9996 11868 10060 11932
rect 3372 11732 3436 11796
rect 13308 11732 13372 11796
rect 1532 11596 1596 11660
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 11284 11460 11348 11524
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 4108 11324 4172 11388
rect 5580 11324 5644 11388
rect 9444 11188 9508 11252
rect 10548 11324 10612 11388
rect 612 11052 676 11116
rect 3004 10916 3068 10980
rect 5212 10976 5276 10980
rect 5212 10920 5226 10976
rect 5226 10920 5276 10976
rect 5212 10916 5276 10920
rect 9628 10916 9692 10980
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 3740 10780 3804 10844
rect 7420 10840 7484 10844
rect 7420 10784 7434 10840
rect 7434 10784 7484 10840
rect 7420 10780 7484 10784
rect 11652 10780 11716 10844
rect 6132 10644 6196 10708
rect 4844 10372 4908 10436
rect 7420 10432 7484 10436
rect 7420 10376 7434 10432
rect 7434 10376 7484 10432
rect 7420 10372 7484 10376
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 7420 10236 7484 10300
rect 7420 9828 7484 9892
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 4660 9692 4724 9756
rect 11468 9692 11532 9756
rect 9628 9420 9692 9484
rect 5948 9284 6012 9348
rect 6500 9284 6564 9348
rect 9076 9344 9140 9348
rect 9076 9288 9090 9344
rect 9090 9288 9140 9344
rect 9076 9284 9140 9288
rect 9628 9284 9692 9348
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11100 9072 11164 9076
rect 12388 9480 12452 9484
rect 12388 9424 12438 9480
rect 12438 9424 12452 9480
rect 12388 9420 12452 9424
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 11100 9016 11114 9072
rect 11114 9016 11164 9072
rect 11100 9012 11164 9016
rect 8340 8876 8404 8940
rect 10916 8936 10980 8940
rect 10916 8880 10930 8936
rect 10930 8880 10980 8936
rect 10916 8876 10980 8880
rect 9628 8740 9692 8804
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 4476 8604 4540 8668
rect 5028 8664 5092 8668
rect 5028 8608 5042 8664
rect 5042 8608 5092 8664
rect 5028 8604 5092 8608
rect 5212 8604 5276 8668
rect 5764 8604 5828 8668
rect 8156 8664 8220 8668
rect 8156 8608 8206 8664
rect 8206 8608 8220 8664
rect 8156 8604 8220 8608
rect 10364 8664 10428 8668
rect 10364 8608 10414 8664
rect 10414 8608 10428 8664
rect 10364 8604 10428 8608
rect 11284 8604 11348 8668
rect 4292 8332 4356 8396
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 5580 8196 5644 8260
rect 8524 8196 8588 8260
rect 10180 8196 10244 8260
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 7420 8060 7484 8124
rect 9812 7924 9876 7988
rect 5396 7788 5460 7852
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 4844 7516 4908 7580
rect 7420 7652 7484 7716
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 7420 7516 7484 7580
rect 14044 7516 14108 7580
rect 8156 7380 8220 7444
rect 13124 7380 13188 7444
rect 5764 7244 5828 7308
rect 6132 7244 6196 7308
rect 4108 7108 4172 7172
rect 8892 7108 8956 7172
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 2452 6972 2516 7036
rect 7420 6972 7484 7036
rect 9996 6972 10060 7036
rect 10180 6972 10244 7036
rect 13860 6972 13924 7036
rect 980 6836 1044 6900
rect 8340 6836 8404 6900
rect 9260 6836 9324 6900
rect 11100 6836 11164 6900
rect 13308 6836 13372 6900
rect 5948 6564 6012 6628
rect 11284 6564 11348 6628
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 4476 6428 4540 6492
rect 796 6292 860 6356
rect 6684 6428 6748 6492
rect 10364 6292 10428 6356
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 4292 5884 4356 5948
rect 9076 5884 9140 5948
rect 10364 5884 10428 5948
rect 3004 5808 3068 5812
rect 3004 5752 3018 5808
rect 3018 5752 3068 5808
rect 3004 5748 3068 5752
rect 3556 5612 3620 5676
rect 12388 5476 12452 5540
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 8892 5340 8956 5404
rect 9628 5340 9692 5404
rect 10180 5340 10244 5404
rect 13492 5400 13556 5404
rect 13492 5344 13506 5400
rect 13506 5344 13556 5400
rect 13492 5340 13556 5344
rect 3372 5204 3436 5268
rect 6316 5204 6380 5268
rect 11652 5204 11716 5268
rect 8156 4932 8220 4996
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 9444 4796 9508 4860
rect 2452 4388 2516 4452
rect 9076 4388 9140 4452
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 3924 3844 3988 3908
rect 8892 3844 8956 3908
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 3004 3300 3068 3364
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 8524 3164 8588 3228
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 10916 3088 10980 3092
rect 10916 3032 10966 3088
rect 10966 3032 10980 3088
rect 10916 3028 10980 3032
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 11284 2620 11348 2684
rect 1532 2484 1596 2548
rect 9076 2484 9140 2548
rect 1716 2348 1780 2412
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 11468 1940 11532 2004
rect 1164 1804 1228 1868
rect 612 1668 676 1732
rect 3740 1532 3804 1596
<< metal4 >>
rect 1944 15808 2264 15824
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 795 14380 861 14381
rect 795 14316 796 14380
rect 860 14316 861 14380
rect 795 14315 861 14316
rect 611 11116 677 11117
rect 611 11052 612 11116
rect 676 11052 677 11116
rect 611 11051 677 11052
rect 614 1733 674 11051
rect 798 6357 858 14315
rect 1163 13972 1229 13973
rect 1163 13908 1164 13972
rect 1228 13908 1229 13972
rect 1163 13907 1229 13908
rect 979 12884 1045 12885
rect 979 12820 980 12884
rect 1044 12820 1045 12884
rect 979 12819 1045 12820
rect 982 6901 1042 12819
rect 979 6900 1045 6901
rect 979 6836 980 6900
rect 1044 6836 1045 6900
rect 979 6835 1045 6836
rect 795 6356 861 6357
rect 795 6292 796 6356
rect 860 6292 861 6356
rect 795 6291 861 6292
rect 1166 1869 1226 13907
rect 1715 13836 1781 13837
rect 1715 13772 1716 13836
rect 1780 13772 1781 13836
rect 1715 13771 1781 13772
rect 1531 11660 1597 11661
rect 1531 11596 1532 11660
rect 1596 11596 1597 11660
rect 1531 11595 1597 11596
rect 1534 2549 1594 11595
rect 1531 2548 1597 2549
rect 1531 2484 1532 2548
rect 1596 2484 1597 2548
rect 1531 2483 1597 2484
rect 1718 2413 1778 13771
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 2604 15264 2924 15824
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 6944 15808 7264 15824
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 4659 13972 4725 13973
rect 4659 13908 4660 13972
rect 4724 13908 4725 13972
rect 4659 13907 4725 13908
rect 2604 13088 2924 13718
rect 3923 13156 3989 13157
rect 3923 13092 3924 13156
rect 3988 13092 3989 13156
rect 3923 13091 3989 13092
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 3555 13020 3621 13021
rect 3555 12956 3556 13020
rect 3620 12956 3621 13020
rect 3555 12955 3621 12956
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 3371 11796 3437 11797
rect 3371 11732 3372 11796
rect 3436 11732 3437 11796
rect 3371 11731 3437 11732
rect 3003 10980 3069 10981
rect 3003 10916 3004 10980
rect 3068 10916 3069 10980
rect 3003 10915 3069 10916
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2451 7036 2517 7037
rect 2451 6972 2452 7036
rect 2516 6972 2517 7036
rect 2451 6971 2517 6972
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 2454 4453 2514 6971
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 3006 5813 3066 10915
rect 3003 5812 3069 5813
rect 3003 5748 3004 5812
rect 3068 5748 3069 5812
rect 3003 5747 3069 5748
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2451 4452 2517 4453
rect 2451 4388 2452 4452
rect 2516 4388 2517 4452
rect 2451 4387 2517 4388
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1715 2412 1781 2413
rect 1715 2348 1716 2412
rect 1780 2348 1781 2412
rect 1715 2347 1781 2348
rect 1944 2128 2264 2688
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 3006 3365 3066 5747
rect 3374 5269 3434 11731
rect 3558 5677 3618 12955
rect 3739 10844 3805 10845
rect 3739 10780 3740 10844
rect 3804 10780 3805 10844
rect 3739 10779 3805 10780
rect 3555 5676 3621 5677
rect 3555 5612 3556 5676
rect 3620 5612 3621 5676
rect 3555 5611 3621 5612
rect 3371 5268 3437 5269
rect 3371 5204 3372 5268
rect 3436 5204 3437 5268
rect 3371 5203 3437 5204
rect 3003 3364 3069 3365
rect 3003 3300 3004 3364
rect 3068 3300 3069 3364
rect 3003 3299 3069 3300
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 1163 1868 1229 1869
rect 1163 1804 1164 1868
rect 1228 1804 1229 1868
rect 1163 1803 1229 1804
rect 611 1732 677 1733
rect 611 1668 612 1732
rect 676 1668 677 1732
rect 611 1667 677 1668
rect 3742 1597 3802 10779
rect 3926 3909 3986 13091
rect 4107 11388 4173 11389
rect 4107 11324 4108 11388
rect 4172 11324 4173 11388
rect 4107 11323 4173 11324
rect 4110 7173 4170 11323
rect 4662 9757 4722 13907
rect 5395 13836 5461 13837
rect 5395 13772 5396 13836
rect 5460 13772 5461 13836
rect 5395 13771 5461 13772
rect 5579 13836 5645 13837
rect 5579 13772 5580 13836
rect 5644 13772 5645 13836
rect 5579 13771 5645 13772
rect 6683 13836 6749 13837
rect 6683 13772 6684 13836
rect 6748 13772 6749 13836
rect 6683 13771 6749 13772
rect 5027 12068 5093 12069
rect 5027 12004 5028 12068
rect 5092 12004 5093 12068
rect 5027 12003 5093 12004
rect 4843 10436 4909 10437
rect 4843 10372 4844 10436
rect 4908 10372 4909 10436
rect 4843 10371 4909 10372
rect 4659 9756 4725 9757
rect 4659 9692 4660 9756
rect 4724 9692 4725 9756
rect 4659 9691 4725 9692
rect 4475 8668 4541 8669
rect 4475 8604 4476 8668
rect 4540 8604 4541 8668
rect 4475 8603 4541 8604
rect 4291 8396 4357 8397
rect 4291 8332 4292 8396
rect 4356 8332 4357 8396
rect 4291 8331 4357 8332
rect 4107 7172 4173 7173
rect 4107 7108 4108 7172
rect 4172 7108 4173 7172
rect 4107 7107 4173 7108
rect 4294 5949 4354 8331
rect 4478 6493 4538 8603
rect 4846 7581 4906 10371
rect 5030 8669 5090 12003
rect 5211 10980 5277 10981
rect 5211 10916 5212 10980
rect 5276 10916 5277 10980
rect 5211 10915 5277 10916
rect 5214 8669 5274 10915
rect 5027 8668 5093 8669
rect 5027 8604 5028 8668
rect 5092 8604 5093 8668
rect 5027 8603 5093 8604
rect 5211 8668 5277 8669
rect 5211 8604 5212 8668
rect 5276 8604 5277 8668
rect 5211 8603 5277 8604
rect 5398 7853 5458 13771
rect 5582 12450 5642 13771
rect 5947 13156 6013 13157
rect 5947 13092 5948 13156
rect 6012 13092 6013 13156
rect 5947 13091 6013 13092
rect 5582 12390 5826 12450
rect 5579 11388 5645 11389
rect 5579 11324 5580 11388
rect 5644 11324 5645 11388
rect 5579 11323 5645 11324
rect 5582 8261 5642 11323
rect 5766 8669 5826 12390
rect 5950 9349 6010 13091
rect 6315 12340 6381 12341
rect 6315 12276 6316 12340
rect 6380 12276 6381 12340
rect 6315 12275 6381 12276
rect 6131 10708 6197 10709
rect 6131 10644 6132 10708
rect 6196 10644 6197 10708
rect 6131 10643 6197 10644
rect 5947 9348 6013 9349
rect 5947 9284 5948 9348
rect 6012 9284 6013 9348
rect 5947 9283 6013 9284
rect 5763 8668 5829 8669
rect 5763 8604 5764 8668
rect 5828 8604 5829 8668
rect 5763 8603 5829 8604
rect 5579 8260 5645 8261
rect 5579 8196 5580 8260
rect 5644 8196 5645 8260
rect 5579 8195 5645 8196
rect 5395 7852 5461 7853
rect 5395 7788 5396 7852
rect 5460 7788 5461 7852
rect 5395 7787 5461 7788
rect 4843 7580 4909 7581
rect 4843 7516 4844 7580
rect 4908 7516 4909 7580
rect 4843 7515 4909 7516
rect 6134 7309 6194 10643
rect 5763 7308 5829 7309
rect 5763 7244 5764 7308
rect 5828 7306 5829 7308
rect 6131 7308 6197 7309
rect 5828 7246 6010 7306
rect 5828 7244 5829 7246
rect 5763 7243 5829 7244
rect 5950 6629 6010 7246
rect 6131 7244 6132 7308
rect 6196 7244 6197 7308
rect 6131 7243 6197 7244
rect 5947 6628 6013 6629
rect 5947 6564 5948 6628
rect 6012 6564 6013 6628
rect 5947 6563 6013 6564
rect 4475 6492 4541 6493
rect 4475 6428 4476 6492
rect 4540 6428 4541 6492
rect 4475 6427 4541 6428
rect 4291 5948 4357 5949
rect 4291 5884 4292 5948
rect 4356 5884 4357 5948
rect 4291 5883 4357 5884
rect 6318 5269 6378 12275
rect 6499 12204 6565 12205
rect 6499 12140 6500 12204
rect 6564 12140 6565 12204
rect 6499 12139 6565 12140
rect 6502 9349 6562 12139
rect 6499 9348 6565 9349
rect 6499 9284 6500 9348
rect 6564 9284 6565 9348
rect 6499 9283 6565 9284
rect 6686 6493 6746 13771
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6944 10368 7264 11392
rect 7604 15264 7924 15824
rect 11944 15808 12264 15824
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 9259 15468 9325 15469
rect 9259 15404 9260 15468
rect 9324 15404 9325 15468
rect 9259 15403 9325 15404
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 8339 13156 8405 13157
rect 8339 13092 8340 13156
rect 8404 13092 8405 13156
rect 8339 13091 8405 13092
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 8155 12068 8221 12069
rect 8155 12004 8156 12068
rect 8220 12004 8221 12068
rect 8155 12003 8221 12004
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7419 10844 7485 10845
rect 7419 10780 7420 10844
rect 7484 10780 7485 10844
rect 7419 10779 7485 10780
rect 7422 10437 7482 10779
rect 7419 10436 7485 10437
rect 7419 10372 7420 10436
rect 7484 10372 7485 10436
rect 7419 10371 7485 10372
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6944 9280 7264 10304
rect 7419 10300 7485 10301
rect 7419 10236 7420 10300
rect 7484 10236 7485 10300
rect 7419 10235 7485 10236
rect 7422 9893 7482 10235
rect 7419 9892 7485 9893
rect 7419 9828 7420 9892
rect 7484 9828 7485 9892
rect 7419 9827 7485 9828
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7419 8124 7485 8125
rect 7419 8060 7420 8124
rect 7484 8060 7485 8124
rect 7419 8059 7485 8060
rect 6944 7104 7264 8058
rect 7422 7717 7482 8059
rect 7419 7716 7485 7717
rect 7419 7652 7420 7716
rect 7484 7652 7485 7716
rect 7419 7651 7485 7652
rect 7604 7648 7924 8672
rect 8158 8669 8218 12003
rect 8342 11933 8402 13091
rect 8523 13020 8589 13021
rect 8523 12956 8524 13020
rect 8588 12956 8589 13020
rect 8523 12955 8589 12956
rect 8526 12069 8586 12955
rect 8523 12068 8589 12069
rect 8523 12004 8524 12068
rect 8588 12004 8589 12068
rect 8523 12003 8589 12004
rect 8339 11932 8405 11933
rect 8339 11868 8340 11932
rect 8404 11868 8405 11932
rect 8339 11867 8405 11868
rect 9075 9348 9141 9349
rect 9075 9284 9076 9348
rect 9140 9284 9141 9348
rect 9075 9283 9141 9284
rect 8339 8940 8405 8941
rect 8339 8876 8340 8940
rect 8404 8876 8405 8940
rect 8339 8875 8405 8876
rect 8155 8668 8221 8669
rect 8155 8604 8156 8668
rect 8220 8604 8221 8668
rect 8155 8603 8221 8604
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7419 7580 7485 7581
rect 7419 7516 7420 7580
rect 7484 7516 7485 7580
rect 7419 7515 7485 7516
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6683 6492 6749 6493
rect 6683 6428 6684 6492
rect 6748 6428 6749 6492
rect 6683 6427 6749 6428
rect 6944 6016 7264 7040
rect 7422 7037 7482 7515
rect 7419 7036 7485 7037
rect 7419 6972 7420 7036
rect 7484 6972 7485 7036
rect 7419 6971 7485 6972
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6315 5268 6381 5269
rect 6315 5204 6316 5268
rect 6380 5204 6381 5268
rect 6315 5203 6381 5204
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 3923 3908 3989 3909
rect 3923 3844 3924 3908
rect 3988 3844 3989 3908
rect 3923 3843 3989 3844
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 6560 7924 7584
rect 8155 7444 8221 7445
rect 8155 7380 8156 7444
rect 8220 7380 8221 7444
rect 8155 7379 8221 7380
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 8158 4997 8218 7379
rect 8342 6901 8402 8875
rect 8523 8260 8589 8261
rect 8523 8196 8524 8260
rect 8588 8196 8589 8260
rect 8523 8195 8589 8196
rect 8339 6900 8405 6901
rect 8339 6836 8340 6900
rect 8404 6836 8405 6900
rect 8339 6835 8405 6836
rect 8155 4996 8221 4997
rect 8155 4932 8156 4996
rect 8220 4932 8221 4996
rect 8155 4931 8221 4932
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 8526 3229 8586 8195
rect 8891 7172 8957 7173
rect 8891 7108 8892 7172
rect 8956 7108 8957 7172
rect 8891 7107 8957 7108
rect 8894 5405 8954 7107
rect 9078 5949 9138 9283
rect 9262 6901 9322 15403
rect 10547 14924 10613 14925
rect 10547 14860 10548 14924
rect 10612 14860 10613 14924
rect 10547 14859 10613 14860
rect 9811 13700 9877 13701
rect 9811 13636 9812 13700
rect 9876 13636 9877 13700
rect 9811 13635 9877 13636
rect 9443 11252 9509 11253
rect 9443 11188 9444 11252
rect 9508 11188 9509 11252
rect 9443 11187 9509 11188
rect 9259 6900 9325 6901
rect 9259 6836 9260 6900
rect 9324 6836 9325 6900
rect 9259 6835 9325 6836
rect 9075 5948 9141 5949
rect 9075 5884 9076 5948
rect 9140 5884 9141 5948
rect 9075 5883 9141 5884
rect 8891 5404 8957 5405
rect 8891 5340 8892 5404
rect 8956 5340 8957 5404
rect 8891 5339 8957 5340
rect 8894 3909 8954 5339
rect 9446 4861 9506 11187
rect 9627 10980 9693 10981
rect 9627 10916 9628 10980
rect 9692 10916 9693 10980
rect 9627 10915 9693 10916
rect 9630 9485 9690 10915
rect 9627 9484 9693 9485
rect 9627 9420 9628 9484
rect 9692 9420 9693 9484
rect 9627 9419 9693 9420
rect 9627 9348 9693 9349
rect 9627 9284 9628 9348
rect 9692 9284 9693 9348
rect 9627 9283 9693 9284
rect 9630 8805 9690 9283
rect 9627 8804 9693 8805
rect 9627 8740 9628 8804
rect 9692 8740 9693 8804
rect 9627 8739 9693 8740
rect 9630 5405 9690 8739
rect 9814 7989 9874 13635
rect 9995 11932 10061 11933
rect 9995 11868 9996 11932
rect 10060 11868 10061 11932
rect 9995 11867 10061 11868
rect 9811 7988 9877 7989
rect 9811 7924 9812 7988
rect 9876 7924 9877 7988
rect 9811 7923 9877 7924
rect 9998 7037 10058 11867
rect 10550 11389 10610 14859
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11651 14244 11717 14245
rect 11651 14180 11652 14244
rect 11716 14180 11717 14244
rect 11651 14179 11717 14180
rect 11467 12068 11533 12069
rect 11467 12004 11468 12068
rect 11532 12004 11533 12068
rect 11467 12003 11533 12004
rect 11283 11524 11349 11525
rect 11283 11460 11284 11524
rect 11348 11460 11349 11524
rect 11283 11459 11349 11460
rect 10547 11388 10613 11389
rect 10547 11324 10548 11388
rect 10612 11324 10613 11388
rect 10547 11323 10613 11324
rect 11099 9076 11165 9077
rect 11099 9012 11100 9076
rect 11164 9012 11165 9076
rect 11099 9011 11165 9012
rect 10915 8940 10981 8941
rect 10915 8876 10916 8940
rect 10980 8876 10981 8940
rect 10915 8875 10981 8876
rect 10363 8668 10429 8669
rect 10363 8604 10364 8668
rect 10428 8604 10429 8668
rect 10363 8603 10429 8604
rect 10179 8260 10245 8261
rect 10179 8196 10180 8260
rect 10244 8196 10245 8260
rect 10179 8195 10245 8196
rect 10182 7037 10242 8195
rect 9995 7036 10061 7037
rect 9995 6972 9996 7036
rect 10060 6972 10061 7036
rect 9995 6971 10061 6972
rect 10179 7036 10245 7037
rect 10179 6972 10180 7036
rect 10244 6972 10245 7036
rect 10179 6971 10245 6972
rect 10182 5405 10242 6971
rect 10366 6357 10426 8603
rect 10363 6356 10429 6357
rect 10363 6292 10364 6356
rect 10428 6292 10429 6356
rect 10363 6291 10429 6292
rect 10366 5949 10426 6291
rect 10363 5948 10429 5949
rect 10363 5884 10364 5948
rect 10428 5884 10429 5948
rect 10363 5883 10429 5884
rect 9627 5404 9693 5405
rect 9627 5340 9628 5404
rect 9692 5340 9693 5404
rect 9627 5339 9693 5340
rect 10179 5404 10245 5405
rect 10179 5340 10180 5404
rect 10244 5340 10245 5404
rect 10179 5339 10245 5340
rect 9443 4860 9509 4861
rect 9443 4796 9444 4860
rect 9508 4796 9509 4860
rect 9443 4795 9509 4796
rect 9075 4452 9141 4453
rect 9075 4388 9076 4452
rect 9140 4388 9141 4452
rect 9075 4387 9141 4388
rect 8891 3908 8957 3909
rect 8891 3844 8892 3908
rect 8956 3844 8957 3908
rect 8891 3843 8957 3844
rect 8523 3228 8589 3229
rect 8523 3164 8524 3228
rect 8588 3164 8589 3228
rect 8523 3163 8589 3164
rect 9078 2549 9138 4387
rect 10918 3093 10978 8875
rect 11102 6901 11162 9011
rect 11286 8669 11346 11459
rect 11470 10570 11530 12003
rect 11654 10845 11714 14179
rect 11944 13632 12264 14656
rect 12604 15264 12924 15824
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12387 14108 12453 14109
rect 12387 14044 12388 14108
rect 12452 14044 12453 14108
rect 12387 14043 12453 14044
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11944 11456 12264 12480
rect 12390 12341 12450 14043
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 14043 13972 14109 13973
rect 14043 13908 14044 13972
rect 14108 13908 14109 13972
rect 14043 13907 14109 13908
rect 13859 13836 13925 13837
rect 13859 13772 13860 13836
rect 13924 13772 13925 13836
rect 13859 13771 13925 13772
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12387 12340 12453 12341
rect 12387 12276 12388 12340
rect 12452 12276 12453 12340
rect 12387 12275 12453 12276
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11651 10844 11717 10845
rect 11651 10780 11652 10844
rect 11716 10780 11717 10844
rect 11651 10779 11717 10780
rect 11470 10510 11714 10570
rect 11467 9756 11533 9757
rect 11467 9692 11468 9756
rect 11532 9692 11533 9756
rect 11467 9691 11533 9692
rect 11283 8668 11349 8669
rect 11283 8604 11284 8668
rect 11348 8604 11349 8668
rect 11283 8603 11349 8604
rect 11099 6900 11165 6901
rect 11099 6836 11100 6900
rect 11164 6836 11165 6900
rect 11099 6835 11165 6836
rect 11283 6628 11349 6629
rect 11283 6564 11284 6628
rect 11348 6564 11349 6628
rect 11283 6563 11349 6564
rect 10915 3092 10981 3093
rect 10915 3028 10916 3092
rect 10980 3028 10981 3092
rect 10915 3027 10981 3028
rect 11286 2685 11346 6563
rect 11283 2684 11349 2685
rect 11283 2620 11284 2684
rect 11348 2620 11349 2684
rect 11283 2619 11349 2620
rect 9075 2548 9141 2549
rect 9075 2484 9076 2548
rect 9140 2484 9141 2548
rect 9075 2483 9141 2484
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11470 2005 11530 9691
rect 11654 5269 11714 10510
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 12604 12000 12924 13024
rect 13123 12340 13189 12341
rect 13123 12276 13124 12340
rect 13188 12276 13189 12340
rect 13123 12275 13189 12276
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12387 9484 12453 9485
rect 12387 9420 12388 9484
rect 12452 9420 12453 9484
rect 12387 9419 12453 9420
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11651 5268 11717 5269
rect 11651 5204 11652 5268
rect 11716 5204 11717 5268
rect 11651 5203 11717 5204
rect 11944 4928 12264 5952
rect 12390 5541 12450 9419
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 13126 7445 13186 12275
rect 13491 12204 13557 12205
rect 13491 12140 13492 12204
rect 13556 12140 13557 12204
rect 13491 12139 13557 12140
rect 13307 11796 13373 11797
rect 13307 11732 13308 11796
rect 13372 11732 13373 11796
rect 13307 11731 13373 11732
rect 13123 7444 13189 7445
rect 13123 7380 13124 7444
rect 13188 7380 13189 7444
rect 13123 7379 13189 7380
rect 13310 6901 13370 11731
rect 13307 6900 13373 6901
rect 13307 6836 13308 6900
rect 13372 6836 13373 6900
rect 13307 6835 13373 6836
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12387 5540 12453 5541
rect 12387 5476 12388 5540
rect 12452 5476 12453 5540
rect 12387 5475 12453 5476
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11944 3294 12264 3776
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 11944 2128 12264 2688
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 13494 5405 13554 12139
rect 13862 7037 13922 13771
rect 14046 7581 14106 13907
rect 14043 7580 14109 7581
rect 14043 7516 14044 7580
rect 14108 7516 14109 7580
rect 14043 7515 14109 7516
rect 13859 7036 13925 7037
rect 13859 6972 13860 7036
rect 13924 6972 13925 7036
rect 13859 6971 13925 6972
rect 13491 5404 13557 5405
rect 13491 5340 13492 5404
rect 13556 5340 13557 5404
rect 13491 5339 13557 5340
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 11467 2004 11533 2005
rect 11467 1940 11468 2004
rect 11532 1940 11533 2004
rect 11467 1939 11533 1940
rect 3739 1596 3805 1597
rect 3739 1532 3740 1596
rect 3804 1532 3805 1596
rect 3739 1531 3805 1532
<< via4 >>
rect 1986 13058 2222 13294
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 2646 13718 2882 13954
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 1986 3058 2222 3294
rect 2646 3718 2882 3954
rect 6986 13058 7222 13294
rect 7646 13718 7882 13954
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 6986 3058 7222 3294
rect 7646 3718 7882 3954
rect 11986 13058 12222 13294
rect 12646 13718 12882 13954
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 11986 3058 12222 3294
rect 12646 3718 12882 3954
<< metal5 >>
rect 1056 13954 14860 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 14860 13954
rect 1056 13676 14860 13718
rect 1056 13294 14860 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 14860 13294
rect 1056 13016 14860 13058
rect 1056 8954 14860 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 14860 8954
rect 1056 8676 14860 8718
rect 1056 8294 14860 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 14860 8294
rect 1056 8016 14860 8058
rect 1056 3954 14860 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 14860 3954
rect 1056 3676 14860 3718
rect 1056 3294 14860 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 14860 3294
rect 1056 3016 14860 3058
use sky130_fd_sc_hd__and3_1  _162_
timestamp 0
transform -1 0 8280 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _163_
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _164_
timestamp 0
transform -1 0 7176 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _165_
timestamp 0
transform 1 0 12512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _166_
timestamp 0
transform -1 0 2484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _167_
timestamp 0
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _168_
timestamp 0
transform -1 0 3496 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _169_
timestamp 0
transform -1 0 13248 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 0
transform -1 0 2760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _171_
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 0
transform -1 0 10488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _173_
timestamp 0
transform 1 0 1472 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _174_
timestamp 0
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 0
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _176_
timestamp 0
transform 1 0 3312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _177_
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _178_
timestamp 0
transform -1 0 9476 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _179_
timestamp 0
transform -1 0 4324 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _180_
timestamp 0
transform 1 0 12512 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _181_
timestamp 0
transform 1 0 12880 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _182_
timestamp 0
transform -1 0 9292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _183_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _184_
timestamp 0
transform 1 0 12972 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _185_
timestamp 0
transform 1 0 10672 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _186_
timestamp 0
transform -1 0 2944 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_2  _187_
timestamp 0
transform -1 0 10304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 0
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _189_
timestamp 0
transform -1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _190_
timestamp 0
transform -1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _191_
timestamp 0
transform 1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _192_
timestamp 0
transform -1 0 5980 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _193_
timestamp 0
transform 1 0 3772 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 0
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _195_
timestamp 0
transform -1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _196_
timestamp 0
transform 1 0 13984 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _197_
timestamp 0
transform 1 0 9292 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _199_
timestamp 0
transform -1 0 10672 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _200_
timestamp 0
transform -1 0 11500 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _201_
timestamp 0
transform 1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _202_
timestamp 0
transform -1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _203_
timestamp 0
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _204_
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _205_
timestamp 0
transform -1 0 14536 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 0
transform -1 0 5520 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _207_
timestamp 0
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _208_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _209_
timestamp 0
transform -1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _210_
timestamp 0
transform 1 0 13984 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _211_
timestamp 0
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _212_
timestamp 0
transform -1 0 11960 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 0
transform -1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 0
transform 1 0 9476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _215_
timestamp 0
transform 1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _216_
timestamp 0
transform 1 0 4140 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _217_
timestamp 0
transform -1 0 12052 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _218_
timestamp 0
transform 1 0 8096 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _219_
timestamp 0
transform -1 0 12052 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _220_
timestamp 0
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _221_
timestamp 0
transform -1 0 8648 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _222_
timestamp 0
transform -1 0 4140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _223_
timestamp 0
transform 1 0 12604 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _224_
timestamp 0
transform 1 0 12512 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _225_
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _227_
timestamp 0
transform 1 0 3496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _228_
timestamp 0
transform -1 0 12052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _229_
timestamp 0
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _230_
timestamp 0
transform 1 0 10764 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _231_
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _232_
timestamp 0
transform -1 0 14536 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _233_
timestamp 0
transform -1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _234_
timestamp 0
transform 1 0 12512 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _235_
timestamp 0
transform -1 0 2116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _236_
timestamp 0
transform -1 0 7728 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 0
transform 1 0 4140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 0
transform -1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _239_
timestamp 0
transform 1 0 3864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _240_
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _241_
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 0
transform -1 0 10580 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 0
transform -1 0 5612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _244_
timestamp 0
transform -1 0 3404 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _245_
timestamp 0
transform -1 0 3404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _246_
timestamp 0
transform -1 0 7360 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _247_
timestamp 0
transform 1 0 4600 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _248_
timestamp 0
transform 1 0 5520 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _249_
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 0
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _251_
timestamp 0
transform 1 0 5520 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _252_
timestamp 0
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _253_
timestamp 0
transform -1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _254_
timestamp 0
transform -1 0 7912 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _255_
timestamp 0
transform 1 0 11316 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _256_
timestamp 0
transform -1 0 5704 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _257_
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _258_
timestamp 0
transform 1 0 11592 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 0
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _260_
timestamp 0
transform 1 0 9108 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _261_
timestamp 0
transform -1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp 0
transform -1 0 7084 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 0
transform -1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _264_
timestamp 0
transform -1 0 14536 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _265_
timestamp 0
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 0
transform -1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _267_
timestamp 0
transform -1 0 9844 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _268_
timestamp 0
transform -1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp 0
transform 1 0 10488 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _270_
timestamp 0
transform 1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _271_
timestamp 0
transform 1 0 5244 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _272_
timestamp 0
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 0
transform -1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _274_
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_2  _275_
timestamp 0
transform -1 0 7820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _276_
timestamp 0
transform -1 0 7636 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _277_
timestamp 0
transform 1 0 4324 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _278_
timestamp 0
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _279_
timestamp 0
transform 1 0 6532 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _280_
timestamp 0
transform 1 0 3128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _281_
timestamp 0
transform -1 0 13524 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 0
transform -1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _283_
timestamp 0
transform -1 0 6992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _284_
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _285_
timestamp 0
transform -1 0 13524 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _286_
timestamp 0
transform -1 0 10856 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _287_
timestamp 0
transform 1 0 2392 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _288_
timestamp 0
transform -1 0 13432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _289_
timestamp 0
transform -1 0 2300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _290_
timestamp 0
transform 1 0 3864 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp 0
transform -1 0 14444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _292_
timestamp 0
transform -1 0 9568 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 0
transform -1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _294_
timestamp 0
transform 1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _295_
timestamp 0
transform 1 0 11960 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _296_
timestamp 0
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _297_
timestamp 0
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 0
transform 1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 0
transform -1 0 12788 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 0
transform 1 0 6440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 0
transform 1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _302_
timestamp 0
transform -1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _303_
timestamp 0
transform 1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 0
transform -1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 0
transform -1 0 11776 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _306_
timestamp 0
transform 1 0 13432 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _310_
timestamp 0
transform -1 0 7268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _311_
timestamp 0
transform 1 0 10488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _312_
timestamp 0
transform -1 0 8188 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _313_
timestamp 0
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 0
transform -1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 0
transform -1 0 12788 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 0
transform -1 0 12512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _317_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 0
transform 1 0 5888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 0
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 0
transform -1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 0
transform -1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp 0
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 0
transform 1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 0
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 0
transform -1 0 13616 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 0
transform 1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 0
transform 1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 0
transform -1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 0
transform -1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _330_
timestamp 0
transform 1 0 9292 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _331_
timestamp 0
transform 1 0 12236 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _332_
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 0
transform 1 0 9568 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _334_
timestamp 0
transform 1 0 5796 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _335_
timestamp 0
transform 1 0 11960 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _336_
timestamp 0
transform 1 0 9568 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _337_
timestamp 0
transform -1 0 10764 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _338_
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 0
transform 1 0 4232 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _340_
timestamp 0
transform -1 0 11132 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _341_
timestamp 0
transform 1 0 8648 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _342_
timestamp 0
transform 1 0 12420 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _343_
timestamp 0
transform -1 0 4232 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _344_
timestamp 0
transform 1 0 12144 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _345_
timestamp 0
transform 1 0 4416 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _346_
timestamp 0
transform -1 0 8832 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _347_
timestamp 0
transform -1 0 7268 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _348_
timestamp 0
transform -1 0 5796 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _349_
timestamp 0
transform -1 0 4600 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _350_
timestamp 0
transform -1 0 8648 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _351_
timestamp 0
transform 1 0 3496 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _352_
timestamp 0
transform -1 0 3404 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _353_
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _354_
timestamp 0
transform 1 0 12052 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _355_
timestamp 0
transform 1 0 9384 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _356_
timestamp 0
transform 1 0 6532 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _357_
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _358_
timestamp 0
transform 1 0 11868 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _359_
timestamp 0
transform -1 0 6440 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _360_
timestamp 0
transform 1 0 4508 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _361_
timestamp 0
transform -1 0 4416 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_1  _370_
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform 1 0 12420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 0
transform -1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 0
transform 1 0 10304 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 0
transform 1 0 7544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__B
timestamp 0
transform -1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__C
timestamp 0
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 0
transform -1 0 6256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A
timestamp 0
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__B
timestamp 0
transform 1 0 12052 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 0
transform 1 0 1564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A1_N
timestamp 0
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A2_N
timestamp 0
transform 1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A1
timestamp 0
transform -1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A2
timestamp 0
transform 1 0 11684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__B1
timestamp 0
transform 1 0 11316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A1
timestamp 0
transform 1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__B1
timestamp 0
transform 1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A1
timestamp 0
transform 1 0 7176 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A2
timestamp 0
transform 1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 0
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__C
timestamp 0
transform 1 0 12420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__D
timestamp 0
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 0
transform 1 0 4508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__C
timestamp 0
transform -1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__D
timestamp 0
transform -1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__B
timestamp 0
transform -1 0 13156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__D
timestamp 0
transform -1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__B
timestamp 0
transform 1 0 8372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A1
timestamp 0
transform 1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A2
timestamp 0
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A2
timestamp 0
transform -1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__C1
timestamp 0
transform 1 0 3128 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 0
transform -1 0 10028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 0
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 0
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__B
timestamp 0
transform -1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 0
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__B
timestamp 0
transform 1 0 5060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 0
transform 1 0 4416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 0
transform 1 0 12512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__B
timestamp 0
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__C
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A1
timestamp 0
transform -1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A2
timestamp 0
transform 1 0 13800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__B
timestamp 0
transform 1 0 9936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A2
timestamp 0
transform -1 0 11408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A3
timestamp 0
transform -1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A_N
timestamp 0
transform -1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__B
timestamp 0
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 0
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__B
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__B
timestamp 0
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 0
transform 1 0 12696 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A2
timestamp 0
transform -1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__C
timestamp 0
transform 1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__C
timestamp 0
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__B
timestamp 0
transform -1 0 13984 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B
timestamp 0
transform 1 0 11684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 0
transform 1 0 11316 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 0
transform -1 0 2760 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__C1
timestamp 0
transform -1 0 11960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 0
transform -1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__B
timestamp 0
transform -1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 0
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__B
timestamp 0
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__B
timestamp 0
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 0
transform 1 0 8372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A2
timestamp 0
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__B
timestamp 0
transform -1 0 7912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__C
timestamp 0
transform 1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 0
transform 1 0 12420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 0
transform 1 0 12328 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 0
transform -1 0 2208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 0
transform -1 0 12144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A1
timestamp 0
transform 1 0 4048 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__B
timestamp 0
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__C
timestamp 0
transform -1 0 3864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__B
timestamp 0
transform 1 0 10580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 0
transform 1 0 13524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A1
timestamp 0
transform 1 0 13064 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__A2
timestamp 0
transform 1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__B1
timestamp 0
transform 1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A
timestamp 0
transform -1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__C
timestamp 0
transform -1 0 2852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 0
transform 1 0 7084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A
timestamp 0
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__B
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__C
timestamp 0
transform 1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__B1
timestamp 0
transform 1 0 6624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__B
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__B
timestamp 0
transform 1 0 5336 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A
timestamp 0
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A3
timestamp 0
transform 1 0 8096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__C1
timestamp 0
transform 1 0 11132 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A4
timestamp 0
transform 1 0 4784 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A
timestamp 0
transform 1 0 11408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__A
timestamp 0
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A
timestamp 0
transform 1 0 13248 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__C
timestamp 0
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A
timestamp 0
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__B2
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A1
timestamp 0
transform 1 0 7084 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__B1
timestamp 0
transform -1 0 8004 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A
timestamp 0
transform -1 0 5152 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__B
timestamp 0
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 0
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 0
transform 1 0 12880 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A2
timestamp 0
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__B1
timestamp 0
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A
timestamp 0
transform -1 0 13892 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A_N
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__B
timestamp 0
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__C
timestamp 0
transform 1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A2
timestamp 0
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__B1
timestamp 0
transform 1 0 2208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__D1
timestamp 0
transform 1 0 3404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__A
timestamp 0
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__B
timestamp 0
transform -1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A1
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__A2
timestamp 0
transform -1 0 3036 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__C
timestamp 0
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 0
transform 1 0 9476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__B
timestamp 0
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A1
timestamp 0
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A2
timestamp 0
transform -1 0 11040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A
timestamp 0
transform -1 0 11960 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A
timestamp 0
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__297__A
timestamp 0
transform 1 0 4416 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 0
transform 1 0 7544 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 0
transform 1 0 12052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__A
timestamp 0
transform 1 0 12972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__302__A
timestamp 0
transform 1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A
timestamp 0
transform -1 0 13248 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A
timestamp 0
transform 1 0 11960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__305__A
timestamp 0
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A
timestamp 0
transform -1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 0
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A
timestamp 0
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__309__A
timestamp 0
transform 1 0 11960 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__A
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A
timestamp 0
transform 1 0 10948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__A
timestamp 0
transform 1 0 8372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A
timestamp 0
transform 1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__A
timestamp 0
transform -1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__316__A
timestamp 0
transform 1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__A
timestamp 0
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A
timestamp 0
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__319__A
timestamp 0
transform 1 0 13892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__320__A
timestamp 0
transform 1 0 9568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__321__A
timestamp 0
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A
timestamp 0
transform -1 0 2944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__323__A
timestamp 0
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__A
timestamp 0
transform -1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A
timestamp 0
transform 1 0 13800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A
timestamp 0
transform -1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__A
timestamp 0
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__A
timestamp 0
transform 1 0 8740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__A
timestamp 0
transform 1 0 9476 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 0
transform 1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output2_A
timestamp 0
transform 1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output4_A
timestamp 0
transform -1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 6992 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 7820 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform 1 0 10120 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform -1 0 8280 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 9016 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_1  clkload0
timestamp 0
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp 0
transform 1 0 5060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 0
transform 1 0 9016 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 0
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_95
timestamp 0
transform 1 0 9844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_99
timestamp 0
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_103
timestamp 0
transform 1 0 10580 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 0
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_116
timestamp 0
transform 1 0 11776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_120
timestamp 0
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 0
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_130
timestamp 0
transform 1 0 13064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_21
timestamp 0
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_26
timestamp 0
transform 1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_30
timestamp 0
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_42
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 0
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_74
timestamp 0
transform 1 0 7912 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_89
timestamp 0
transform 1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_104
timestamp 0
transform 1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_108
timestamp 0
transform 1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_144
timestamp 0
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_8
timestamp 0
transform 1 0 1840 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_12
timestamp 0
transform 1 0 2208 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_16
timestamp 0
transform 1 0 2576 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_59
timestamp 0
transform 1 0 6532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_68
timestamp 0
transform 1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_72
timestamp 0
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 0
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_94
timestamp 0
transform 1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_98
timestamp 0
transform 1 0 10120 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_110
timestamp 0
transform 1 0 11224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_118
timestamp 0
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_122
timestamp 0
transform 1 0 12328 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_125
timestamp 0
transform 1 0 12604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_132
timestamp 0
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_138
timestamp 0
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_18
timestamp 0
transform 1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_22
timestamp 0
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_26
timestamp 0
transform 1 0 3496 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_38
timestamp 0
transform 1 0 4600 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_46
timestamp 0
transform 1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_66
timestamp 0
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_70
timestamp 0
transform 1 0 7544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_73
timestamp 0
transform 1 0 7820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_77
timestamp 0
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_80
timestamp 0
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_85
timestamp 0
transform 1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_89
timestamp 0
transform 1 0 9292 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_101
timestamp 0
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_124
timestamp 0
transform 1 0 12512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_128
timestamp 0
transform 1 0 12880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_132
timestamp 0
transform 1 0 13248 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_136
timestamp 0
transform 1 0 13616 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_24
timestamp 0
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_33
timestamp 0
transform 1 0 4140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_72
timestamp 0
transform 1 0 7728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 0
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_93
timestamp 0
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_110
timestamp 0
transform 1 0 11224 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_119
timestamp 0
transform 1 0 12052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_123
timestamp 0
transform 1 0 12420 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_127
timestamp 0
transform 1 0 12788 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_131
timestamp 0
transform 1 0 13156 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_21
timestamp 0
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_24
timestamp 0
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_29
timestamp 0
transform 1 0 3772 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_33
timestamp 0
transform 1 0 4140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_36
timestamp 0
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_41
timestamp 0
transform 1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_50
timestamp 0
transform 1 0 5704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_62
timestamp 0
transform 1 0 6808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_84
timestamp 0
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_119
timestamp 0
transform 1 0 12052 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_9
timestamp 0
transform 1 0 1932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_13
timestamp 0
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_17
timestamp 0
transform 1 0 2668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp 0
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_34
timestamp 0
transform 1 0 4232 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_44
timestamp 0
transform 1 0 5152 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_69
timestamp 0
transform 1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_80
timestamp 0
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_89
timestamp 0
transform 1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_93
timestamp 0
transform 1 0 9660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_105
timestamp 0
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_108
timestamp 0
transform 1 0 11040 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_23
timestamp 0
transform 1 0 3220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_37
timestamp 0
transform 1 0 4508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_41
timestamp 0
transform 1 0 4876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_73
timestamp 0
transform 1 0 7820 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_77
timestamp 0
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_85
timestamp 0
transform 1 0 8924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_97
timestamp 0
transform 1 0 10028 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_106
timestamp 0
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_119
timestamp 0
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_144
timestamp 0
transform 1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_23
timestamp 0
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 0
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_73
timestamp 0
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 0
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_89
timestamp 0
transform 1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_93
timestamp 0
transform 1 0 9660 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_118
timestamp 0
transform 1 0 11960 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_144
timestamp 0
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_6
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_12
timestamp 0
transform 1 0 2208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 0
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_76
timestamp 0
transform 1 0 8096 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_88
timestamp 0
transform 1 0 9200 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_96
timestamp 0
transform 1 0 9936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_103
timestamp 0
transform 1 0 10580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_107
timestamp 0
transform 1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_136
timestamp 0
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_11
timestamp 0
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_21
timestamp 0
transform 1 0 3036 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_24
timestamp 0
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_49
timestamp 0
transform 1 0 5612 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_57
timestamp 0
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_64
timestamp 0
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_68
timestamp 0
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 0
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_103
timestamp 0
transform 1 0 10580 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_113
timestamp 0
transform 1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_117
timestamp 0
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_137
timestamp 0
transform 1 0 13708 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_23
timestamp 0
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_46
timestamp 0
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_61
timestamp 0
transform 1 0 6716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_73
timestamp 0
transform 1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_107
timestamp 0
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_122
timestamp 0
transform 1 0 12328 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_130
timestamp 0
transform 1 0 13064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_134
timestamp 0
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_11
timestamp 0
transform 1 0 2116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_23
timestamp 0
transform 1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_54
timestamp 0
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_58
timestamp 0
transform 1 0 6440 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_111
timestamp 0
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_117
timestamp 0
transform 1 0 11868 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_134
timestamp 0
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 0
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_11
timestamp 0
transform 1 0 2116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_23
timestamp 0
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_30
timestamp 0
transform 1 0 3864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_64
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_74
timestamp 0
transform 1 0 7912 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_78
timestamp 0
transform 1 0 8280 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_91
timestamp 0
transform 1 0 9476 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_116
timestamp 0
transform 1 0 11776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_120
timestamp 0
transform 1 0 12144 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_127
timestamp 0
transform 1 0 12788 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_131
timestamp 0
transform 1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_136
timestamp 0
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_140
timestamp 0
transform 1 0 13984 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_25
timestamp 0
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_79
timestamp 0
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_91
timestamp 0
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_105
timestamp 0
transform 1 0 10764 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_117
timestamp 0
transform 1 0 11868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_127
timestamp 0
transform 1 0 12788 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_134
timestamp 0
transform 1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 0
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_9
timestamp 0
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_19
timestamp 0
transform 1 0 2852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_25
timestamp 0
transform 1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_29
timestamp 0
transform 1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_37
timestamp 0
transform 1 0 4508 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_50
timestamp 0
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_72
timestamp 0
transform 1 0 7728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_84
timestamp 0
transform 1 0 8832 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_100
timestamp 0
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_117
timestamp 0
transform 1 0 11868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_127
timestamp 0
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_131
timestamp 0
transform 1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_25
timestamp 0
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_33
timestamp 0
transform 1 0 4140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_64
timestamp 0
transform 1 0 6992 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_68
timestamp 0
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_72
timestamp 0
transform 1 0 7728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 0
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_105
timestamp 0
transform 1 0 10764 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_113
timestamp 0
transform 1 0 11500 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_135
timestamp 0
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_30
timestamp 0
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_34
timestamp 0
transform 1 0 4232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_41
timestamp 0
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_52
timestamp 0
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_67
timestamp 0
transform 1 0 7268 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_71
timestamp 0
transform 1 0 7636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_121
timestamp 0
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_130
timestamp 0
transform 1 0 13064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_135
timestamp 0
transform 1 0 13524 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_143
timestamp 0
transform 1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_23
timestamp 0
transform 1 0 3220 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_78
timestamp 0
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_92
timestamp 0
transform 1 0 9568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_96
timestamp 0
transform 1 0 9936 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_106
timestamp 0
transform 1 0 10856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_110
timestamp 0
transform 1 0 11224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_114
timestamp 0
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_118
timestamp 0
transform 1 0 11960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_122
timestamp 0
transform 1 0 12328 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 0
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_34
timestamp 0
transform 1 0 4232 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_41
timestamp 0
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_45
timestamp 0
transform 1 0 5244 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_64
timestamp 0
transform 1 0 6992 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_68
timestamp 0
transform 1 0 7360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_80
timestamp 0
transform 1 0 8464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_106
timestamp 0
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_116
timestamp 0
transform 1 0 11776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_120
timestamp 0
transform 1 0 12144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_124
timestamp 0
transform 1 0 12512 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_132
timestamp 0
transform 1 0 13248 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_138
timestamp 0
transform 1 0 13800 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_145
timestamp 0
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_10
timestamp 0
transform 1 0 2024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_14
timestamp 0
transform 1 0 2392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_21
timestamp 0
transform 1 0 3036 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_25
timestamp 0
transform 1 0 3404 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_40
timestamp 0
transform 1 0 4784 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_71
timestamp 0
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_75
timestamp 0
transform 1 0 8004 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_114
timestamp 0
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_144
timestamp 0
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_7
timestamp 0
transform 1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_36
timestamp 0
transform 1 0 4416 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_40
timestamp 0
transform 1 0 4784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_44
timestamp 0
transform 1 0 5152 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_61
timestamp 0
transform 1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_67
timestamp 0
transform 1 0 7268 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_75
timestamp 0
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_92
timestamp 0
transform 1 0 9568 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_104
timestamp 0
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_117
timestamp 0
transform 1 0 11868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_121
timestamp 0
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_127
timestamp 0
transform 1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_136
timestamp 0
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_145
timestamp 0
transform 1 0 14444 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_8
timestamp 0
transform 1 0 1840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_12
timestamp 0
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_17
timestamp 0
transform 1 0 2668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_21
timestamp 0
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_51
timestamp 0
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_63
timestamp 0
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_75
timestamp 0
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_105
timestamp 0
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_113
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_117
timestamp 0
transform 1 0 11868 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_125
timestamp 0
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_129
timestamp 0
transform 1 0 12972 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_137
timestamp 0
transform 1 0 13708 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_11
timestamp 0
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_17
timestamp 0
transform 1 0 2668 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_38
timestamp 0
transform 1 0 4600 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_68
timestamp 0
transform 1 0 7360 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_72
timestamp 0
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_84
timestamp 0
transform 1 0 8832 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_96
timestamp 0
transform 1 0 9936 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_102
timestamp 0
transform 1 0 10488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_109
timestamp 0
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_119
timestamp 0
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_123
timestamp 0
transform 1 0 12420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_135
timestamp 0
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_141
timestamp 0
transform 1 0 14076 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_11
timestamp 0
transform 1 0 2116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_19
timestamp 0
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_35
timestamp 0
transform 1 0 4324 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_39
timestamp 0
transform 1 0 4692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_51
timestamp 0
transform 1 0 5796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_55
timestamp 0
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_57
timestamp 0
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_61
timestamp 0
transform 1 0 6716 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 0
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_94
timestamp 0
transform 1 0 9752 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_103
timestamp 0
transform 1 0 10580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_111
timestamp 0
transform 1 0 11316 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_113
timestamp 0
transform 1 0 11500 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_131
timestamp 0
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_135
timestamp 0
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_144
timestamp 0
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output2
timestamp 0
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output3
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output4
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 0
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output6
timestamp 0
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 0
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 0
transform 1 0 14260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_25
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_26
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_27
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_28
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_29
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_30
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_31
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_32
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_33
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_34
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_35
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_36
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_37
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_38
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_39
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_40
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_41
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_42
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_43
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_44
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_45
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_46
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_47
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_48
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_49
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  project3_9
timestamp 0
transform 1 0 14260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  project3_10
timestamp 0
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  project3_11
timestamp 0
transform -1 0 14536 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  project3_12
timestamp 0
transform -1 0 14536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  project3_13
timestamp 0
transform -1 0 14536 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  project3_14
timestamp 0
transform -1 0 14168 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  project3_15
timestamp 0
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  project3_16
timestamp 0
transform -1 0 13984 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_50
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_51
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_52
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_53
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_54
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_55
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_56
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_57
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_58
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_59
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_60
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_61
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_62
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_63
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_65
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_66
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_67
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_68
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_70
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_71
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_72
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_73
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_74
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_75
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_76
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_77
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_78
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_79
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_80
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_81
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_82
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_83
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_84
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_85
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_86
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_87
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_88
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_89
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_90
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_91
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_92
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_93
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_94
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_95
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_96
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_97
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_98
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_99
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_100
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_101
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_102
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_103
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_104
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_105
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_106
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_107
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_108
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_109
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_110
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_111
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_112
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_113
timestamp 0
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_114
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_115
timestamp 0
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_116
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
<< labels >>
rlabel metal1 s 7958 15232 7958 15232 4 VGND
rlabel metal1 s 7958 15776 7958 15776 4 VPWR
rlabel metal1 s 8280 8058 8280 8058 4 _000_
rlabel metal3 s 9660 12716 9660 12716 4 _001_
rlabel metal2 s 3174 4539 3174 4539 4 _002_
rlabel metal2 s 13018 7072 13018 7072 4 _003_
rlabel metal1 s 4002 7446 4002 7446 4 _004_
rlabel metal2 s 14444 7548 14444 7548 4 _005_
rlabel metal1 s 5842 3706 5842 3706 4 _006_
rlabel metal1 s 8924 5134 8924 5134 4 _007_
rlabel metal1 s 7360 7514 7360 7514 4 _008_
rlabel metal4 s 1564 7072 1564 7072 4 _009_
rlabel metal3 s 4278 14909 4278 14909 4 _010_
rlabel metal1 s 13984 2618 13984 2618 4 _011_
rlabel metal2 s 12282 12835 12282 12835 4 _012_
rlabel metal1 s 4094 5814 4094 5814 4 _013_
rlabel metal1 s 2392 2482 2392 2482 4 _014_
rlabel metal3 s 7981 13804 7981 13804 4 _015_
rlabel metal1 s 10810 12886 10810 12886 4 _016_
rlabel metal3 s 4462 9061 4462 9061 4 _017_
rlabel metal2 s 14030 7208 14030 7208 4 _018_
rlabel metal1 s 12052 9894 12052 9894 4 _019_
rlabel metal1 s 1334 14518 1334 14518 4 _020_
rlabel metal1 s 5796 4522 5796 4522 4 _021_
rlabel metal1 s 11730 3094 11730 3094 4 _022_
rlabel metal1 s 9384 13430 9384 13430 4 _023_
rlabel metal1 s 14030 3094 14030 3094 4 _024_
rlabel metal1 s 11454 14858 11454 14858 4 _025_
rlabel metal1 s 4462 7446 4462 7446 4 _026_
rlabel metal2 s 4462 4386 4462 4386 4 _027_
rlabel metal2 s 6670 10336 6670 10336 4 _028_
rlabel metal4 s 13340 9316 13340 9316 4 _029_
rlabel metal4 s 13156 9860 13156 9860 4 _030_
rlabel metal1 s 12558 5100 12558 5100 4 _031_
rlabel metal2 s 6578 5304 6578 5304 4 _032_
rlabel metal2 s 13294 3808 13294 3808 4 _033_
rlabel metal1 s 1610 13158 1610 13158 4 _034_
rlabel metal3 s 8809 1564 8809 1564 4 _035_
rlabel metal3 s 6233 12716 6233 12716 4 _036_
rlabel metal3 s 10741 13668 10741 13668 4 _037_
rlabel metal1 s 13662 13192 13662 13192 4 _038_
rlabel metal1 s 12558 6630 12558 6630 4 _039_
rlabel metal2 s 13846 7276 13846 7276 4 _040_
rlabel metal3 s 4232 7956 4232 7956 4 _041_
rlabel metal2 s 11730 8296 11730 8296 4 _042_
rlabel metal1 s 7682 10982 7682 10982 4 _043_
rlabel metal1 s 8602 2414 8602 2414 4 _044_
rlabel metal1 s 2254 4760 2254 4760 4 _045_
rlabel metal1 s 12604 14042 12604 14042 4 _046_
rlabel metal2 s 8786 14297 8786 14297 4 _047_
rlabel metal2 s 6026 14586 6026 14586 4 _048_
rlabel metal3 s 14214 15555 14214 15555 4 _049_
rlabel metal2 s 2530 2159 2530 2159 4 _050_
rlabel metal2 s 13938 11458 13938 11458 4 _051_
rlabel metal4 s 1012 9860 1012 9860 4 _052_
rlabel metal2 s 10166 9010 10166 9010 4 _053_
rlabel metal2 s 14398 4335 14398 4335 4 _054_
rlabel metal2 s 13478 7650 13478 7650 4 _055_
rlabel metal1 s 9062 4794 9062 4794 4 _056_
rlabel metal1 s 4823 12138 4823 12138 4 _057_
rlabel metal1 s 7820 5882 7820 5882 4 _058_
rlabel metal3 s 6463 15436 6463 15436 4 _059_
rlabel metal1 s 12098 5746 12098 5746 4 _060_
rlabel metal2 s 6854 10234 6854 10234 4 _061_
rlabel metal1 s 2162 3978 2162 3978 4 _062_
rlabel metal4 s 3979 13124 3979 13124 4 _063_
rlabel metal2 s 2806 11526 2806 11526 4 _064_
rlabel metal2 s 2392 3876 2392 3876 4 _065_
rlabel metal1 s 2392 7854 2392 7854 4 _066_
rlabel metal1 s 10350 6358 10350 6358 4 _067_
rlabel metal1 s 13110 8942 13110 8942 4 _068_
rlabel metal4 s 644 6392 644 6392 4 _069_
rlabel metal2 s 6854 3519 6854 3519 4 _070_
rlabel metal1 s 10626 14790 10626 14790 4 _071_
rlabel metal1 s 1472 3706 1472 3706 4 _072_
rlabel metal2 s 9706 11424 9706 11424 4 _073_
rlabel metal1 s 2162 4624 2162 4624 4 _074_
rlabel metal1 s 4416 15470 4416 15470 4 _075_
rlabel metal1 s 8188 3502 8188 3502 4 _076_
rlabel metal2 s 13294 14178 13294 14178 4 _077_
rlabel metal1 s 13432 9350 13432 9350 4 _078_
rlabel metal2 s 13386 12036 13386 12036 4 _079_
rlabel metal1 s 4048 6766 4048 6766 4 _080_
rlabel metal2 s 13478 14127 13478 14127 4 _081_
rlabel metal1 s 2346 4556 2346 4556 4 _082_
rlabel metal1 s 2714 4624 2714 4624 4 _083_
rlabel metal1 s 2438 4726 2438 4726 4 _084_
rlabel metal1 s 13938 8398 13938 8398 4 _085_
rlabel metal1 s 13294 2856 13294 2856 4 _086_
rlabel metal2 s 2438 11832 2438 11832 4 _087_
rlabel metal2 s 2714 7105 2714 7105 4 _088_
rlabel metal2 s 1242 7412 1242 7412 4 _089_
rlabel metal1 s 9338 3468 9338 3468 4 _090_
rlabel metal1 s 14536 10438 14536 10438 4 _091_
rlabel metal2 s 13018 4097 13018 4097 4 _092_
rlabel metal1 s 10810 3162 10810 3162 4 _093_
rlabel metal3 s 4991 13804 4991 13804 4 _094_
rlabel metal1 s 9154 13940 9154 13940 4 _095_
rlabel metal2 s 14306 4199 14306 4199 4 _096_
rlabel metal2 s 14766 5321 14766 5321 4 _097_
rlabel metal3 s 14122 3621 14122 3621 4 _098_
rlabel metal1 s 8510 2890 8510 2890 4 _099_
rlabel metal1 s 13938 13974 13938 13974 4 _100_
rlabel metal1 s 15042 13838 15042 13838 4 _101_
rlabel metal1 s 13846 2992 13846 2992 4 _102_
rlabel metal1 s 1886 13226 1886 13226 4 _103_
rlabel metal1 s 14030 2992 14030 2992 4 _104_
rlabel metal3 s 4761 13940 4761 13940 4 _105_
rlabel metal1 s 10488 13498 10488 13498 4 _106_
rlabel metal2 s 8510 14484 8510 14484 4 _107_
rlabel metal2 s 4002 11305 4002 11305 4 _108_
rlabel metal2 s 2990 5729 2990 5729 4 _109_
rlabel metal2 s 1610 14535 1610 14535 4 _110_
rlabel metal2 s 1886 11339 1886 11339 4 _111_
rlabel metal3 s 1495 13940 1495 13940 4 _112_
rlabel metal1 s 3404 3026 3404 3026 4 _113_
rlabel metal1 s 1610 14960 1610 14960 4 _114_
rlabel metal2 s 13386 5338 13386 5338 4 _115_
rlabel metal1 s 14030 5576 14030 5576 4 _116_
rlabel metal2 s 14122 7089 14122 7089 4 _117_
rlabel metal2 s 10534 10642 10534 10642 4 _118_
rlabel metal1 s 7206 10710 7206 10710 4 _119_
rlabel metal1 s 4370 9452 4370 9452 4 _120_
rlabel metal2 s 5750 11441 5750 11441 4 _121_
rlabel metal2 s 6026 5253 6026 5253 4 _122_
rlabel metal1 s 9246 12682 9246 12682 4 _123_
rlabel metal2 s 10350 15130 10350 15130 4 _124_
rlabel metal1 s 7130 3536 7130 3536 4 _125_
rlabel metal1 s 3036 5882 3036 5882 4 _126_
rlabel metal1 s 10948 5542 10948 5542 4 _127_
rlabel metal2 s 6026 6936 6026 6936 4 _128_
rlabel metal4 s 5635 13804 5635 13804 4 _129_
rlabel metal1 s 11362 6256 11362 6256 4 _130_
rlabel metal2 s 7222 7718 7222 7718 4 _131_
rlabel metal2 s 11569 4590 11569 4590 4 _132_
rlabel metal2 s 8602 6919 8602 6919 4 _133_
rlabel metal1 s 9338 13736 9338 13736 4 _134_
rlabel metal1 s 11868 6290 11868 6290 4 _135_
rlabel metal1 s 7038 14926 7038 14926 4 _136_
rlabel metal1 s 14306 7514 14306 7514 4 _137_
rlabel metal1 s 10442 14042 10442 14042 4 _138_
rlabel metal1 s 14536 8262 14536 8262 4 _139_
rlabel metal2 s 12466 8806 12466 8806 4 _140_
rlabel metal1 s 13294 12818 13294 12818 4 _141_
rlabel metal1 s 4646 5712 4646 5712 4 _142_
rlabel metal2 s 10258 8364 10258 8364 4 _143_
rlabel metal2 s 5934 5372 5934 5372 4 _144_
rlabel metal1 s 5436 5338 5436 5338 4 _145_
rlabel metal1 s 6026 10642 6026 10642 4 _146_
rlabel metal1 s 7038 6290 7038 6290 4 _147_
rlabel metal2 s 7314 6460 7314 6460 4 _148_
rlabel metal1 s 7130 7242 7130 7242 4 _149_
rlabel metal1 s 6578 7480 6578 7480 4 _150_
rlabel metal2 s 13294 12682 13294 12682 4 _151_
rlabel metal1 s 13424 12070 13424 12070 4 _152_
rlabel metal3 s 12788 11152 12788 11152 4 _153_
rlabel metal2 s 9614 4709 9614 4709 4 _154_
rlabel metal2 s 1978 14178 1978 14178 4 _155_
rlabel metal2 s 9522 5287 9522 5287 4 _156_
rlabel metal2 s 4278 12954 4278 12954 4 _157_
rlabel metal1 s 5428 4590 5428 4590 4 _158_
rlabel metal2 s 9568 11764 9568 11764 4 _159_
rlabel metal2 s 10166 2142 10166 2142 4 _160_
rlabel metal1 s 14168 15130 14168 15130 4 _161_
rlabel metal3 s 1579 4420 1579 4420 4 clk
rlabel metal1 s 8694 12886 8694 12886 4 clknet_0_clk
rlabel metal2 s 5842 3536 5842 3536 4 clknet_2_0__leaf_clk
rlabel metal1 s 9430 8908 9430 8908 4 clknet_2_1__leaf_clk
rlabel metal2 s 4370 14127 4370 14127 4 clknet_2_2__leaf_clk
rlabel metal1 s 9844 12614 9844 12614 4 clknet_2_3__leaf_clk
rlabel metal1 s 2576 3706 2576 3706 4 decoder.digit\[0\]
rlabel metal1 s 8970 12240 8970 12240 4 decoder.digit\[1\]
rlabel metal2 s 2254 7616 2254 7616 4 decoder.digit\[2\]
rlabel metal1 s 2668 9486 2668 9486 4 decoder.digit\[3\]
rlabel metal1 s 4002 14008 4002 14008 4 net1
rlabel metal3 s 14490 8789 14490 8789 4 net10
rlabel metal3 s 14490 9877 14490 9877 4 net11
rlabel metal2 s 14490 10999 14490 10999 4 net12
rlabel metal3 s 14490 12053 14490 12053 4 net13
rlabel metal2 s 14122 13039 14122 13039 4 net14
rlabel metal3 s 14490 14229 14490 14229 4 net15
rlabel metal3 s 13938 15317 13938 15317 4 net16
rlabel metal1 s 2990 5610 2990 5610 4 net2
rlabel metal1 s 13662 2414 13662 2414 4 net3
rlabel metal4 s 1771 13804 1771 13804 4 net4
rlabel metal2 s 12926 4845 12926 4845 4 net5
rlabel metal1 s 14628 12614 14628 12614 4 net6
rlabel metal2 s 13938 6035 13938 6035 4 net7
rlabel metal2 s 14306 6970 14306 6970 4 net8
rlabel metal2 s 14490 15691 14490 15691 4 net9
rlabel metal1 s 2254 10676 2254 10676 4 one_second_counter\[0\]
rlabel metal1 s 9200 13158 9200 13158 4 one_second_counter\[10\]
rlabel metal1 s 12834 10200 12834 10200 4 one_second_counter\[11\]
rlabel metal2 s 2438 15232 2438 15232 4 one_second_counter\[12\]
rlabel metal1 s 2024 14790 2024 14790 4 one_second_counter\[13\]
rlabel metal1 s 12742 15436 12742 15436 4 one_second_counter\[14\]
rlabel metal1 s 5888 7854 5888 7854 4 one_second_counter\[15\]
rlabel metal1 s 4830 7922 4830 7922 4 one_second_counter\[16\]
rlabel metal1 s 3726 6766 3726 6766 4 one_second_counter\[17\]
rlabel metal2 s 4290 6766 4290 6766 4 one_second_counter\[18\]
rlabel metal2 s 8878 11050 8878 11050 4 one_second_counter\[19\]
rlabel metal2 s 5750 7344 5750 7344 4 one_second_counter\[1\]
rlabel metal1 s 10166 2346 10166 2346 4 one_second_counter\[20\]
rlabel metal2 s 9614 2074 9614 2074 4 one_second_counter\[21\]
rlabel metal1 s 6578 2584 6578 2584 4 one_second_counter\[22\]
rlabel metal1 s 10350 2482 10350 2482 4 one_second_counter\[23\]
rlabel metal1 s 8694 13294 8694 13294 4 one_second_counter\[24\]
rlabel metal1 s 10396 4794 10396 4794 4 one_second_counter\[25\]
rlabel metal1 s 8786 9894 8786 9894 4 one_second_counter\[26\]
rlabel metal1 s 10166 7378 10166 7378 4 one_second_counter\[2\]
rlabel metal2 s 11362 6273 11362 6273 4 one_second_counter\[3\]
rlabel metal1 s 8234 4658 8234 4658 4 one_second_counter\[4\]
rlabel metal1 s 12604 2550 12604 2550 4 one_second_counter\[5\]
rlabel metal1 s 9246 9520 9246 9520 4 one_second_counter\[6\]
rlabel metal2 s 9062 13260 9062 13260 4 one_second_counter\[7\]
rlabel metal1 s 13202 13872 13202 13872 4 one_second_counter\[8\]
rlabel metal1 s 7268 7174 7268 7174 4 one_second_counter\[9\]
rlabel metal1 s 10902 15130 10902 15130 4 one_second_enable
rlabel metal3 s 1050 13396 1050 13396 4 rst
rlabel metal2 s 13662 1717 13662 1717 4 seg0
rlabel metal3 s 13938 2261 13938 2261 4 seg1
rlabel metal2 s 13938 3791 13938 3791 4 seg2
rlabel metal3 s 13938 4437 13938 4437 4 seg3
rlabel metal2 s 14490 5151 14490 5151 4 seg4
rlabel metal2 s 14214 6885 14214 6885 4 seg5
rlabel metal3 s 14490 7701 14490 7701 4 seg6
flabel metal5 s 1056 13676 14860 13996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8676 14860 8996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3676 14860 3996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 12604 2128 12924 15824 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7604 2128 7924 15824 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2604 2128 2924 15824 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 13016 14860 13336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 8016 14860 8336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3016 14860 3336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 11944 2128 12264 15824 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 6944 2128 7264 15824 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1944 2128 2264 15824 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 15200 8712 16000 8832 0 FreeSans 600 0 0 0 an0
port 3 nsew
flabel metal3 s 15200 9800 16000 9920 0 FreeSans 600 0 0 0 an1
port 4 nsew
flabel metal3 s 15200 10888 16000 11008 0 FreeSans 600 0 0 0 an2
port 5 nsew
flabel metal3 s 15200 11976 16000 12096 0 FreeSans 600 0 0 0 an3
port 6 nsew
flabel metal3 s 15200 13064 16000 13184 0 FreeSans 600 0 0 0 an4
port 7 nsew
flabel metal3 s 15200 14152 16000 14272 0 FreeSans 600 0 0 0 an5
port 8 nsew
flabel metal3 s 15200 15240 16000 15360 0 FreeSans 600 0 0 0 an6
port 9 nsew
flabel metal3 s 15200 16328 16000 16448 0 FreeSans 600 0 0 0 an7
port 10 nsew
flabel metal3 s 0 4360 800 4480 0 FreeSans 600 0 0 0 clk
port 11 nsew
flabel metal3 s 0 13336 800 13456 0 FreeSans 600 0 0 0 rst
port 12 nsew
flabel metal3 s 15200 1096 16000 1216 0 FreeSans 600 0 0 0 seg0
port 13 nsew
flabel metal3 s 15200 2184 16000 2304 0 FreeSans 600 0 0 0 seg1
port 14 nsew
flabel metal3 s 15200 3272 16000 3392 0 FreeSans 600 0 0 0 seg2
port 15 nsew
flabel metal3 s 15200 4360 16000 4480 0 FreeSans 600 0 0 0 seg3
port 16 nsew
flabel metal3 s 15200 5448 16000 5568 0 FreeSans 600 0 0 0 seg4
port 17 nsew
flabel metal3 s 15200 6536 16000 6656 0 FreeSans 600 0 0 0 seg5
port 18 nsew
flabel metal3 s 15200 7624 16000 7744 0 FreeSans 600 0 0 0 seg6
port 19 nsew
<< properties >>
string FIXED_BBOX 0 0 16000 18000
<< end >>
