VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO project4
  CLASS BLOCK ;
  FOREIGN project4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END A1[4]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.168500 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.921000 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END A2[4]
  PIN A3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END A3[0]
  PIN A3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END A3[1]
  PIN A3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END A3[2]
  PIN A3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END A3[3]
  PIN A3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END A3[4]
  PIN ALU_result[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END ALU_result[0]
  PIN ALU_result[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 163.240 400.000 163.840 ;
    END
  END ALU_result[10]
  PIN ALU_result[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 268.640 400.000 269.240 ;
    END
  END ALU_result[11]
  PIN ALU_result[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 200.640 400.000 201.240 ;
    END
  END ALU_result[12]
  PIN ALU_result[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.040 400.000 204.640 ;
    END
  END ALU_result[13]
  PIN ALU_result[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END ALU_result[14]
  PIN ALU_result[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 231.240 400.000 231.840 ;
    END
  END ALU_result[15]
  PIN ALU_result[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 210.840 400.000 211.440 ;
    END
  END ALU_result[16]
  PIN ALU_result[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.240 400.000 214.840 ;
    END
  END ALU_result[17]
  PIN ALU_result[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 217.640 400.000 218.240 ;
    END
  END ALU_result[18]
  PIN ALU_result[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 400.000 238.640 ;
    END
  END ALU_result[19]
  PIN ALU_result[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.040 400.000 187.640 ;
    END
  END ALU_result[1]
  PIN ALU_result[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 224.440 400.000 225.040 ;
    END
  END ALU_result[20]
  PIN ALU_result[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 234.640 400.000 235.240 ;
    END
  END ALU_result[21]
  PIN ALU_result[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.040 400.000 221.640 ;
    END
  END ALU_result[22]
  PIN ALU_result[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 265.240 400.000 265.840 ;
    END
  END ALU_result[23]
  PIN ALU_result[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 227.840 400.000 228.440 ;
    END
  END ALU_result[24]
  PIN ALU_result[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 244.840 400.000 245.440 ;
    END
  END ALU_result[25]
  PIN ALU_result[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 241.440 400.000 242.040 ;
    END
  END ALU_result[26]
  PIN ALU_result[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 261.840 400.000 262.440 ;
    END
  END ALU_result[27]
  PIN ALU_result[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.040 400.000 255.640 ;
    END
  END ALU_result[28]
  PIN ALU_result[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 251.640 400.000 252.240 ;
    END
  END ALU_result[29]
  PIN ALU_result[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.240 400.000 180.840 ;
    END
  END ALU_result[2]
  PIN ALU_result[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 258.440 400.000 259.040 ;
    END
  END ALU_result[30]
  PIN ALU_result[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.240 400.000 248.840 ;
    END
  END ALU_result[31]
  PIN ALU_result[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 190.440 400.000 191.040 ;
    END
  END ALU_result[3]
  PIN ALU_result[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 166.640 400.000 167.240 ;
    END
  END ALU_result[4]
  PIN ALU_result[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.840 400.000 194.440 ;
    END
  END ALU_result[5]
  PIN ALU_result[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 400.000 170.640 ;
    END
  END ALU_result[6]
  PIN ALU_result[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.840 400.000 177.440 ;
    END
  END ALU_result[7]
  PIN ALU_result[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 207.440 400.000 208.040 ;
    END
  END ALU_result[8]
  PIN ALU_result[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.840 400.000 160.440 ;
    END
  END ALU_result[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 10.640 39.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.020 10.640 64.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.020 10.640 89.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 113.020 10.640 114.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.020 10.640 139.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 163.020 10.640 164.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 10.640 189.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 213.020 10.640 214.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 238.020 10.640 239.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 263.020 10.640 264.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 288.020 10.640 289.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 313.020 10.640 314.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 338.020 10.640 339.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 363.020 10.640 364.620 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 388.020 10.640 389.620 389.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.380 394.460 19.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.380 394.460 44.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.380 394.460 69.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 93.380 394.460 94.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 118.380 394.460 119.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 143.380 394.460 144.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 168.380 394.460 169.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 193.380 394.460 194.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 218.380 394.460 219.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 243.380 394.460 244.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 268.380 394.460 269.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 293.380 394.460 294.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 318.380 394.460 319.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 343.380 394.460 344.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 368.380 394.460 369.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.720 10.640 61.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.720 10.640 86.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 109.720 10.640 111.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.720 10.640 136.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.720 10.640 161.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 10.640 186.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.720 10.640 211.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.720 10.640 236.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 259.720 10.640 261.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.720 10.640 286.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 309.720 10.640 311.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.720 10.640 336.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 359.720 10.640 361.320 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.720 10.640 386.320 389.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 394.460 16.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.080 394.460 41.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 65.080 394.460 66.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 90.080 394.460 91.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 115.080 394.460 116.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 140.080 394.460 141.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 165.080 394.460 166.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 190.080 394.460 191.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 215.080 394.460 216.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 240.080 394.460 241.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 265.080 394.460 266.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 290.080 394.460 291.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 315.080 394.460 316.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 340.080 394.460 341.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 365.080 394.460 366.680 ;
    END
  END VPWR
  PIN WD3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END WD3[0]
  PIN WD3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END WD3[10]
  PIN WD3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END WD3[11]
  PIN WD3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END WD3[12]
  PIN WD3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END WD3[13]
  PIN WD3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END WD3[14]
  PIN WD3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END WD3[15]
  PIN WD3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END WD3[16]
  PIN WD3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END WD3[17]
  PIN WD3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END WD3[18]
  PIN WD3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END WD3[19]
  PIN WD3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END WD3[1]
  PIN WD3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 396.000 228.990 400.000 ;
    END
  END WD3[20]
  PIN WD3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 396.000 142.050 400.000 ;
    END
  END WD3[21]
  PIN WD3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 396.000 225.770 400.000 ;
    END
  END WD3[22]
  PIN WD3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 161.090 396.000 161.370 400.000 ;
    END
  END WD3[23]
  PIN WD3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 396.000 190.350 400.000 ;
    END
  END WD3[24]
  PIN WD3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 396.000 222.550 400.000 ;
    END
  END WD3[25]
  PIN WD3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 396.000 174.250 400.000 ;
    END
  END WD3[26]
  PIN WD3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 396.000 158.150 400.000 ;
    END
  END WD3[27]
  PIN WD3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 396.000 154.930 400.000 ;
    END
  END WD3[28]
  PIN WD3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 231.930 396.000 232.210 400.000 ;
    END
  END WD3[29]
  PIN WD3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END WD3[2]
  PIN WD3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END WD3[30]
  PIN WD3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END WD3[31]
  PIN WD3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END WD3[3]
  PIN WD3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END WD3[4]
  PIN WD3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END WD3[5]
  PIN WD3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END WD3[6]
  PIN WD3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END WD3[7]
  PIN WD3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.840 400.000 143.440 ;
    END
  END WD3[8]
  PIN WD3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END WD3[9]
  PIN WE3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END WE3
  PIN opcode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 183.640 400.000 184.240 ;
    END
  END opcode[0]
  PIN opcode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 173.440 400.000 174.040 ;
    END
  END opcode[1]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 394.410 389.150 ;
      LAYER li1 ;
        RECT 5.520 10.795 394.220 389.045 ;
      LAYER met1 ;
        RECT 4.210 10.640 394.220 389.200 ;
      LAYER met2 ;
        RECT 4.230 395.720 141.490 396.000 ;
        RECT 142.330 395.720 154.370 396.000 ;
        RECT 155.210 395.720 157.590 396.000 ;
        RECT 158.430 395.720 160.810 396.000 ;
        RECT 161.650 395.720 173.690 396.000 ;
        RECT 174.530 395.720 189.790 396.000 ;
        RECT 190.630 395.720 221.990 396.000 ;
        RECT 222.830 395.720 225.210 396.000 ;
        RECT 226.050 395.720 228.430 396.000 ;
        RECT 229.270 395.720 231.650 396.000 ;
        RECT 232.490 395.720 392.750 396.000 ;
        RECT 4.230 4.280 392.750 395.720 ;
        RECT 4.230 3.670 38.450 4.280 ;
        RECT 39.290 3.670 89.970 4.280 ;
        RECT 90.810 3.670 138.270 4.280 ;
        RECT 139.110 3.670 144.710 4.280 ;
        RECT 145.550 3.670 147.930 4.280 ;
        RECT 148.770 3.670 151.150 4.280 ;
        RECT 151.990 3.670 157.590 4.280 ;
        RECT 158.430 3.670 160.810 4.280 ;
        RECT 161.650 3.670 164.030 4.280 ;
        RECT 164.870 3.670 167.250 4.280 ;
        RECT 168.090 3.670 176.910 4.280 ;
        RECT 177.750 3.670 186.570 4.280 ;
        RECT 187.410 3.670 212.330 4.280 ;
        RECT 213.170 3.670 218.770 4.280 ;
        RECT 219.610 3.670 225.210 4.280 ;
        RECT 226.050 3.670 241.310 4.280 ;
        RECT 242.150 3.670 244.530 4.280 ;
        RECT 245.370 3.670 250.970 4.280 ;
        RECT 251.810 3.670 267.070 4.280 ;
        RECT 267.910 3.670 276.730 4.280 ;
        RECT 277.570 3.670 308.930 4.280 ;
        RECT 309.770 3.670 312.150 4.280 ;
        RECT 312.990 3.670 315.370 4.280 ;
        RECT 316.210 3.670 318.590 4.280 ;
        RECT 319.430 3.670 392.750 4.280 ;
      LAYER met3 ;
        RECT 3.990 269.640 396.000 389.125 ;
        RECT 3.990 268.240 395.600 269.640 ;
        RECT 3.990 266.240 396.000 268.240 ;
        RECT 3.990 264.840 395.600 266.240 ;
        RECT 3.990 262.840 396.000 264.840 ;
        RECT 3.990 261.440 395.600 262.840 ;
        RECT 3.990 259.440 396.000 261.440 ;
        RECT 3.990 258.040 395.600 259.440 ;
        RECT 3.990 256.040 396.000 258.040 ;
        RECT 4.400 254.640 395.600 256.040 ;
        RECT 3.990 252.640 396.000 254.640 ;
        RECT 3.990 251.240 395.600 252.640 ;
        RECT 3.990 249.240 396.000 251.240 ;
        RECT 3.990 247.840 395.600 249.240 ;
        RECT 3.990 245.840 396.000 247.840 ;
        RECT 3.990 244.440 395.600 245.840 ;
        RECT 3.990 242.440 396.000 244.440 ;
        RECT 3.990 241.040 395.600 242.440 ;
        RECT 3.990 239.040 396.000 241.040 ;
        RECT 3.990 237.640 395.600 239.040 ;
        RECT 3.990 235.640 396.000 237.640 ;
        RECT 4.400 234.240 395.600 235.640 ;
        RECT 3.990 232.240 396.000 234.240 ;
        RECT 3.990 230.840 395.600 232.240 ;
        RECT 3.990 228.840 396.000 230.840 ;
        RECT 4.400 227.440 395.600 228.840 ;
        RECT 3.990 225.440 396.000 227.440 ;
        RECT 4.400 224.040 395.600 225.440 ;
        RECT 3.990 222.040 396.000 224.040 ;
        RECT 4.400 220.640 395.600 222.040 ;
        RECT 3.990 218.640 396.000 220.640 ;
        RECT 4.400 217.240 395.600 218.640 ;
        RECT 3.990 215.240 396.000 217.240 ;
        RECT 4.400 213.840 395.600 215.240 ;
        RECT 3.990 211.840 396.000 213.840 ;
        RECT 4.400 210.440 395.600 211.840 ;
        RECT 3.990 208.440 396.000 210.440 ;
        RECT 4.400 207.040 395.600 208.440 ;
        RECT 3.990 205.040 396.000 207.040 ;
        RECT 4.400 203.640 395.600 205.040 ;
        RECT 3.990 201.640 396.000 203.640 ;
        RECT 3.990 200.240 395.600 201.640 ;
        RECT 3.990 198.240 396.000 200.240 ;
        RECT 3.990 196.840 395.600 198.240 ;
        RECT 3.990 194.840 396.000 196.840 ;
        RECT 3.990 193.440 395.600 194.840 ;
        RECT 3.990 191.440 396.000 193.440 ;
        RECT 4.400 190.040 395.600 191.440 ;
        RECT 3.990 188.040 396.000 190.040 ;
        RECT 3.990 186.640 395.600 188.040 ;
        RECT 3.990 184.640 396.000 186.640 ;
        RECT 3.990 183.240 395.600 184.640 ;
        RECT 3.990 181.240 396.000 183.240 ;
        RECT 3.990 179.840 395.600 181.240 ;
        RECT 3.990 177.840 396.000 179.840 ;
        RECT 4.400 176.440 395.600 177.840 ;
        RECT 3.990 174.440 396.000 176.440 ;
        RECT 3.990 173.040 395.600 174.440 ;
        RECT 3.990 171.040 396.000 173.040 ;
        RECT 3.990 169.640 395.600 171.040 ;
        RECT 3.990 167.640 396.000 169.640 ;
        RECT 4.400 166.240 395.600 167.640 ;
        RECT 3.990 164.240 396.000 166.240 ;
        RECT 3.990 162.840 395.600 164.240 ;
        RECT 3.990 160.840 396.000 162.840 ;
        RECT 3.990 159.440 395.600 160.840 ;
        RECT 3.990 157.440 396.000 159.440 ;
        RECT 3.990 156.040 395.600 157.440 ;
        RECT 3.990 150.640 396.000 156.040 ;
        RECT 4.400 149.240 396.000 150.640 ;
        RECT 3.990 143.840 396.000 149.240 ;
        RECT 3.990 142.440 395.600 143.840 ;
        RECT 3.990 10.715 396.000 142.440 ;
      LAYER met4 ;
        RECT 56.415 13.095 59.320 386.745 ;
        RECT 61.720 13.095 62.620 386.745 ;
        RECT 65.020 13.095 84.320 386.745 ;
        RECT 86.720 13.095 87.620 386.745 ;
        RECT 90.020 13.095 109.320 386.745 ;
        RECT 111.720 13.095 112.620 386.745 ;
        RECT 115.020 13.095 134.320 386.745 ;
        RECT 136.720 13.095 137.620 386.745 ;
        RECT 140.020 13.095 159.320 386.745 ;
        RECT 161.720 13.095 162.620 386.745 ;
        RECT 165.020 13.095 184.320 386.745 ;
        RECT 186.720 13.095 187.620 386.745 ;
        RECT 190.020 13.095 209.320 386.745 ;
        RECT 211.720 13.095 212.620 386.745 ;
        RECT 215.020 13.095 234.320 386.745 ;
        RECT 236.720 13.095 237.620 386.745 ;
        RECT 240.020 13.095 259.320 386.745 ;
        RECT 261.720 13.095 262.620 386.745 ;
        RECT 265.020 13.095 284.320 386.745 ;
        RECT 286.720 13.095 287.620 386.745 ;
        RECT 290.020 13.095 309.320 386.745 ;
        RECT 311.720 13.095 312.620 386.745 ;
        RECT 315.020 13.095 334.320 386.745 ;
        RECT 336.720 13.095 337.620 386.745 ;
        RECT 340.020 13.095 359.320 386.745 ;
        RECT 361.720 13.095 362.185 386.745 ;
      LAYER met5 ;
        RECT 146.860 82.500 241.380 84.100 ;
  END
END project4
END LIBRARY

