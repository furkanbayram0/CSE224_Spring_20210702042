* NGSPICE file created from project4.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

.subckt project4 A1[0] A1[1] A1[2] A1[3] A1[4] A2[0] A2[1] A2[2] A2[3] A2[4] A3[0]
+ A3[1] A3[2] A3[3] A3[4] ALU_result[0] ALU_result[10] ALU_result[11] ALU_result[12]
+ ALU_result[13] ALU_result[14] ALU_result[15] ALU_result[16] ALU_result[17] ALU_result[18]
+ ALU_result[19] ALU_result[1] ALU_result[20] ALU_result[21] ALU_result[22] ALU_result[23]
+ ALU_result[24] ALU_result[25] ALU_result[26] ALU_result[27] ALU_result[28] ALU_result[29]
+ ALU_result[2] ALU_result[30] ALU_result[31] ALU_result[3] ALU_result[4] ALU_result[5]
+ ALU_result[6] ALU_result[7] ALU_result[8] ALU_result[9] CLK VGND VPWR WD3[0] WD3[10]
+ WD3[11] WD3[12] WD3[13] WD3[14] WD3[15] WD3[16] WD3[17] WD3[18] WD3[19] WD3[1] WD3[20]
+ WD3[21] WD3[22] WD3[23] WD3[24] WD3[25] WD3[26] WD3[27] WD3[28] WD3[29] WD3[2] WD3[30]
+ WD3[31] WD3[3] WD3[4] WD3[5] WD3[6] WD3[7] WD3[8] WD3[9] WE3 opcode[0] opcode[1]
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7963_ RF.registers\[18\]\[29\] _3448_ _3938_ VGND VGND VPWR VPWR _3948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6914_ _3375_ VGND VGND VPWR VPWR _3376_ sky130_fd_sc_hd__clkbuf_8
X_7894_ _3911_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6845_ _3091_ _3302_ VGND VGND VPWR VPWR _3339_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9564_ clknet_leaf_16_CLK _0724_ VGND VGND VPWR VPWR RF.registers\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6776_ net13 net12 net11 VGND VGND VPWR VPWR _3302_ sky130_fd_sc_hd__or3b_2
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9495_ clknet_leaf_33_CLK _0655_ VGND VGND VPWR VPWR RF.registers\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5727_ _2062_ _2479_ VGND VGND VPWR VPWR _2480_ sky130_fd_sc_hd__nor2_1
X_8515_ _4240_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__clkbuf_1
X_8446_ _3003_ _3411_ VGND VGND VPWR VPWR _4204_ sky130_fd_sc_hd__nor2_2
XFILLER_0_115_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5658_ _2410_ _2412_ _2097_ VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4609_ _1254_ _1364_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_107_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8377_ _4167_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__clkbuf_1
X_5589_ _1799_ _2141_ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7328_ _3611_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7259_ _3060_ RF.registers\[29\]\[18\] _3566_ VGND VGND VPWR VPWR _3575_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_6_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_82_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4960_ _1655_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_82_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4891_ RF.registers\[28\]\[0\] RF.registers\[29\]\[0\] RF.registers\[30\]\[0\] RF.registers\[31\]\[0\]
+ net1 net2 VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6630_ _3079_ RF.registers\[15\]\[27\] _3217_ VGND VGND VPWR VPWR _3225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6561_ _3187_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8300_ _3009_ RF.registers\[13\]\[27\] _4119_ VGND VGND VPWR VPWR _4127_ sky130_fd_sc_hd__mux2_1
X_5512_ RF.registers\[0\]\[6\] RF.registers\[1\]\[6\] RF.registers\[2\]\[6\] RF.registers\[3\]\[6\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2268_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6492_ _3149_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9280_ clknet_leaf_74_CLK _0440_ VGND VGND VPWR VPWR RF.registers\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8231_ _4090_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5443_ RF.registers\[16\]\[10\] RF.registers\[17\]\[10\] RF.registers\[18\]\[10\]
+ RF.registers\[19\]\[10\] _2050_ _2052_ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8162_ RF.registers\[24\]\[26\] _3442_ _4047_ VGND VGND VPWR VPWR _4054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5374_ _2128_ _2129_ _2044_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7113_ net23 VGND VGND VPWR VPWR _3493_ sky130_fd_sc_hd__buf_2
X_4325_ _1079_ _1080_ _1040_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__mux2_1
X_8093_ _4017_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_93_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7044_ net34 VGND VGND VPWR VPWR _3446_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8995_ clknet_leaf_75_CLK _0155_ VGND VGND VPWR VPWR RF.registers\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_7946_ _3939_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__clkbuf_1
X_7877_ _3134_ RF.registers\[23\]\[20\] _3902_ VGND VGND VPWR VPWR _3903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6828_ _3330_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6759_ _3293_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9547_ clknet_leaf_89_CLK _0707_ VGND VGND VPWR VPWR RF.registers\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9478_ clknet_leaf_62_CLK _0638_ VGND VGND VPWR VPWR RF.registers\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8429_ _4195_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5090_ RF.registers\[28\]\[17\] RF.registers\[29\]\[17\] RF.registers\[30\]\[17\]
+ RF.registers\[31\]\[17\] _1689_ _1693_ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7800_ RF.registers\[9\]\[16\] _3489_ _3855_ VGND VGND VPWR VPWR _3862_ sky130_fd_sc_hd__mux2_1
X_5992_ _2347_ _2622_ VGND VGND VPWR VPWR _2732_ sky130_fd_sc_hd__nor2_1
X_8780_ clknet_leaf_82_CLK _0964_ VGND VGND VPWR VPWR RF.registers\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_4943_ _1696_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__buf_4
X_7731_ _3825_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__clkbuf_1
X_7662_ RF.registers\[2\]\[15\] _3487_ _3783_ VGND VGND VPWR VPWR _3789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9401_ clknet_leaf_27_CLK _0561_ VGND VGND VPWR VPWR RF.registers\[24\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4874_ RF.registers\[4\]\[18\] RF.registers\[5\]\[18\] RF.registers\[6\]\[18\] RF.registers\[7\]\[18\]
+ _1173_ _1175_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__mux4_1
X_6613_ _3062_ RF.registers\[15\]\[19\] _3206_ VGND VGND VPWR VPWR _3216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7593_ _3752_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9332_ clknet_leaf_37_CLK _0492_ VGND VGND VPWR VPWR RF.registers\[21\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6544_ _3178_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6475_ net28 VGND VGND VPWR VPWR _3139_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_95_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9263_ clknet_leaf_5_CLK _0423_ VGND VGND VPWR VPWR RF.registers\[23\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8214_ _4081_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__clkbuf_1
X_5426_ RF.registers\[16\]\[11\] RF.registers\[17\]\[11\] RF.registers\[18\]\[11\]
+ RF.registers\[19\]\[11\] _1675_ _1692_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9194_ clknet_leaf_2_CLK _0354_ VGND VGND VPWR VPWR RF.registers\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8145_ RF.registers\[24\]\[18\] _3493_ _4036_ VGND VGND VPWR VPWR _4045_ sky130_fd_sc_hd__mux2_1
X_5357_ _1702_ VGND VGND VPWR VPWR _2113_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8076_ _4008_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__clkbuf_1
X_5288_ _1684_ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__buf_4
X_4308_ _1062_ _1063_ _1035_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__mux2_1
X_7027_ _3436_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8978_ clknet_leaf_42_CLK _0138_ VGND VGND VPWR VPWR RF.registers\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_7929_ _3930_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4590_ _1344_ _1345_ _1259_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6260_ _2984_ _2985_ VGND VGND VPWR VPWR _2986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5211_ RF.registers\[24\]\[27\] RF.registers\[25\]\[27\] RF.registers\[26\]\[27\]
+ RF.registers\[27\]\[27\] _1767_ _1768_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__mux4_1
X_6191_ _1996_ _2903_ _2919_ VGND VGND VPWR VPWR _2920_ sky130_fd_sc_hd__o21ba_1
X_5142_ _1897_ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_90_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5073_ _1824_ _1825_ _1826_ _1827_ _1713_ _1828_ VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__mux4_2
X_8901_ clknet_leaf_64_CLK _0061_ VGND VGND VPWR VPWR RF.registers\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8832_ clknet_leaf_70_CLK _1016_ VGND VGND VPWR VPWR RF.registers\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8763_ clknet_leaf_45_CLK _0947_ VGND VGND VPWR VPWR RF.registers\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_5975_ _2573_ _2591_ VGND VGND VPWR VPWR _2716_ sky130_fd_sc_hd__and2_1
X_8694_ clknet_leaf_33_CLK _0878_ VGND VGND VPWR VPWR RF.registers\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_4926_ RF.registers\[20\]\[23\] RF.registers\[21\]\[23\] RF.registers\[22\]\[23\]
+ RF.registers\[23\]\[23\] _1676_ _1681_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7714_ _3816_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__clkbuf_1
X_4857_ _1190_ _1612_ _1205_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7645_ RF.registers\[2\]\[7\] _3470_ _3772_ VGND VGND VPWR VPWR _3780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7576_ _3743_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9315_ clknet_leaf_76_CLK _0475_ VGND VGND VPWR VPWR RF.registers\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_4788_ RF.registers\[16\]\[10\] RF.registers\[17\]\[10\] RF.registers\[18\]\[10\]
+ RF.registers\[19\]\[10\] _1041_ _1043_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__mux4_1
X_6527_ RF.registers\[0\]\[11\] _3116_ _3168_ VGND VGND VPWR VPWR _3170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6458_ _3127_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__clkbuf_1
X_9246_ clknet_leaf_68_CLK _0406_ VGND VGND VPWR VPWR RF.registers\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6389_ _3079_ RF.registers\[22\]\[27\] _3065_ VGND VGND VPWR VPWR _3080_ sky130_fd_sc_hd__mux2_1
X_9177_ clknet_leaf_50_CLK _0337_ VGND VGND VPWR VPWR RF.registers\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xclkload90 clknet_leaf_35_CLK VGND VGND VPWR VPWR clkload90/Y sky130_fd_sc_hd__clkinv_1
X_5409_ RF.registers\[20\]\[12\] RF.registers\[21\]\[12\] RF.registers\[22\]\[12\]
+ RF.registers\[23\]\[12\] _2113_ _2114_ VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8128_ _4024_ VGND VGND VPWR VPWR _4036_ sky130_fd_sc_hd__buf_4
XFILLER_0_11_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8059_ _3999_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5760_ _2481_ _2484_ _2480_ VGND VGND VPWR VPWR _2512_ sky130_fd_sc_hd__a21o_1
X_5691_ _2441_ _2444_ _2040_ VGND VGND VPWR VPWR _2445_ sky130_fd_sc_hd__mux2_1
X_4711_ _1465_ _1466_ _1036_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7430_ _3666_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_1
X_4642_ _1392_ _1394_ _1397_ _1078_ _1057_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4573_ _1189_ _1328_ _1078_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__a21o_1
X_7361_ _3025_ RF.registers\[26\]\[1\] _3628_ VGND VGND VPWR VPWR _3630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6312_ _3027_ RF.registers\[22\]\[2\] _3023_ VGND VGND VPWR VPWR _3028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7292_ _3025_ RF.registers\[31\]\[1\] _3591_ VGND VGND VPWR VPWR _3593_ sky130_fd_sc_hd__mux2_1
X_9100_ clknet_leaf_3_CLK _0260_ VGND VGND VPWR VPWR RF.registers\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6243_ _2420_ _2968_ _2501_ VGND VGND VPWR VPWR _2969_ sky130_fd_sc_hd__mux2_1
X_9031_ clknet_leaf_57_CLK _0191_ VGND VGND VPWR VPWR RF.registers\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6174_ _1996_ _2903_ VGND VGND VPWR VPWR _2904_ sky130_fd_sc_hd__xor2_2
X_5125_ _1720_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5056_ RF.registers\[8\]\[18\] RF.registers\[9\]\[18\] RF.registers\[10\]\[18\] RF.registers\[11\]\[18\]
+ _1689_ _1693_ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8815_ clknet_leaf_84_CLK _0999_ VGND VGND VPWR VPWR RF.registers\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5958_ _2104_ _2696_ _2700_ VGND VGND VPWR VPWR _2701_ sky130_fd_sc_hd__o21a_1
X_8746_ clknet_leaf_87_CLK _0930_ VGND VGND VPWR VPWR RF.registers\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_4909_ _1664_ _1060_ _1084_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5889_ _2246_ _2616_ _2634_ VGND VGND VPWR VPWR _2635_ sky130_fd_sc_hd__a21oi_1
X_8677_ clknet_leaf_79_CLK _0861_ VGND VGND VPWR VPWR RF.registers\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7628_ _3770_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7559_ _3087_ RF.registers\[27\]\[31\] _3699_ VGND VGND VPWR VPWR _3734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9229_ clknet_leaf_12_CLK _0389_ VGND VGND VPWR VPWR RF.registers\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 _1735_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6930_ _3384_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6861_ RF.registers\[5\]\[7\] _3107_ _3340_ VGND VGND VPWR VPWR _3348_ sky130_fd_sc_hd__mux2_1
X_8600_ clknet_leaf_39_CLK _0784_ VGND VGND VPWR VPWR RF.registers\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5812_ _2559_ _2560_ VGND VGND VPWR VPWR _2561_ sky130_fd_sc_hd__or2b_1
XFILLER_0_57_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9580_ clknet_leaf_10_CLK _0740_ VGND VGND VPWR VPWR RF.registers\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6792_ _3311_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5743_ _2040_ _2335_ VGND VGND VPWR VPWR _2495_ sky130_fd_sc_hd__nor2_1
X_8531_ RF.registers\[10\]\[8\] net44 _4244_ VGND VGND VPWR VPWR _4249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5674_ _1168_ _2230_ VGND VGND VPWR VPWR _2428_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8462_ RF.registers\[11\]\[7\] net43 _4205_ VGND VGND VPWR VPWR _4213_ sky130_fd_sc_hd__mux2_1
X_4625_ RF.registers\[12\]\[24\] RF.registers\[13\]\[24\] RF.registers\[14\]\[24\]
+ RF.registers\[15\]\[24\] _1351_ _1352_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7413_ _3077_ RF.registers\[26\]\[26\] _3650_ VGND VGND VPWR VPWR _3657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8393_ _4176_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4556_ RF.registers\[0\]\[27\] RF.registers\[1\]\[27\] RF.registers\[2\]\[27\] RF.registers\[3\]\[27\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__mux4_1
X_7344_ _3077_ RF.registers\[31\]\[26\] _3613_ VGND VGND VPWR VPWR _3620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7275_ _3583_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
X_4487_ RF.registers\[28\]\[20\] RF.registers\[29\]\[20\] RF.registers\[30\]\[20\]
+ RF.registers\[31\]\[20\] _1207_ _1208_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9014_ clknet_leaf_32_CLK _0174_ VGND VGND VPWR VPWR RF.registers\[31\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6226_ _2951_ _2952_ VGND VGND VPWR VPWR _2953_ sky130_fd_sc_hd__or2b_1
X_6157_ _1447_ _1384_ _2871_ _2741_ VGND VGND VPWR VPWR _2888_ sky130_fd_sc_hd__a31o_1
X_5108_ RF.registers\[20\]\[16\] RF.registers\[21\]\[16\] RF.registers\[22\]\[16\]
+ RF.registers\[23\]\[16\] _1705_ _1708_ VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6088_ _2040_ _2797_ VGND VGND VPWR VPWR _2823_ sky130_fd_sc_hd__nor2_1
X_5039_ RF.registers\[0\]\[20\] RF.registers\[1\]\[20\] RF.registers\[2\]\[20\] RF.registers\[3\]\[20\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8729_ clknet_leaf_34_CLK _0913_ VGND VGND VPWR VPWR RF.registers\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput64 net64 VGND VGND VPWR VPWR ALU_result[23] sky130_fd_sc_hd__buf_1
Xoutput53 net53 VGND VGND VPWR VPWR ALU_result[13] sky130_fd_sc_hd__buf_1
Xoutput75 net75 VGND VGND VPWR VPWR ALU_result[4] sky130_fd_sc_hd__buf_1
XFILLER_0_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4410_ _1057_ _1153_ _1157_ _1161_ _1165_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a32o_2
XFILLER_0_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5390_ RF.registers\[16\]\[13\] RF.registers\[17\]\[13\] RF.registers\[18\]\[13\]
+ RF.registers\[19\]\[13\] _1673_ _1690_ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4341_ _1095_ _1096_ _1040_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7060_ _3457_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
X_4272_ A2[1] VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__buf_4
X_6011_ _2730_ _2740_ _2750_ _2621_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__o22a_1
XFILLER_0_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7962_ _3947_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__clkbuf_1
X_6913_ _3155_ _3302_ VGND VGND VPWR VPWR _3375_ sky130_fd_sc_hd__nor2_2
X_7893_ _3011_ RF.registers\[23\]\[28\] _3902_ VGND VGND VPWR VPWR _3911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6844_ _3338_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9563_ clknet_leaf_45_CLK _0723_ VGND VGND VPWR VPWR RF.registers\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6775_ _3301_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9494_ clknet_leaf_47_CLK _0654_ VGND VGND VPWR VPWR RF.registers\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5726_ _2039_ _2478_ VGND VGND VPWR VPWR _2479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8514_ RF.registers\[10\]\[0\] net14 _3007_ VGND VGND VPWR VPWR _4240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8445_ _4203_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5657_ _1166_ _2411_ _1145_ VGND VGND VPWR VPWR _2412_ sky130_fd_sc_hd__o21ai_1
X_4608_ _1362_ _1363_ _1190_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__mux2_1
X_8376_ RF.registers\[16\]\[31\] _3452_ _4132_ VGND VGND VPWR VPWR _4167_ sky130_fd_sc_hd__mux2_1
X_5588_ _2341_ _2342_ VGND VGND VPWR VPWR _2343_ sky130_fd_sc_hd__and2b_1
X_4539_ RF.registers\[12\]\[26\] RF.registers\[13\]\[26\] RF.registers\[14\]\[26\]
+ RF.registers\[15\]\[26\] _1172_ _1279_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__mux4_1
X_7327_ _3060_ RF.registers\[31\]\[18\] _3602_ VGND VGND VPWR VPWR _3611_ sky130_fd_sc_hd__mux2_1
X_7258_ _3574_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6209_ _2875_ _2892_ VGND VGND VPWR VPWR _2937_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_129_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7189_ RF.registers\[7\]\[18\] _3493_ _3528_ VGND VGND VPWR VPWR _3537_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4890_ _1643_ _1644_ _1645_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6560_ RF.registers\[0\]\[27\] _3009_ _3179_ VGND VGND VPWR VPWR _3187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5511_ RF.registers\[4\]\[6\] RF.registers\[5\]\[6\] RF.registers\[6\]\[6\] RF.registers\[7\]\[6\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2267_ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6491_ RF.registers\[17\]\[28\] _3011_ _3135_ VGND VGND VPWR VPWR _3149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8230_ RF.registers\[1\]\[26\] _3442_ _4083_ VGND VGND VPWR VPWR _4090_ sky130_fd_sc_hd__mux2_1
X_5442_ RF.registers\[20\]\[10\] RF.registers\[21\]\[10\] RF.registers\[22\]\[10\]
+ RF.registers\[23\]\[10\] _2050_ _2052_ VGND VGND VPWR VPWR _2198_ sky130_fd_sc_hd__mux4_1
X_8161_ _4053_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5373_ RF.registers\[24\]\[14\] RF.registers\[25\]\[14\] RF.registers\[26\]\[14\]
+ RF.registers\[27\]\[14\] _1674_ _1691_ VGND VGND VPWR VPWR _2129_ sky130_fd_sc_hd__mux4_1
X_8092_ RF.registers\[20\]\[25\] _3508_ _4011_ VGND VGND VPWR VPWR _4017_ sky130_fd_sc_hd__mux2_1
X_7112_ _3492_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4324_ RF.registers\[0\]\[5\] RF.registers\[1\]\[5\] RF.registers\[2\]\[5\] RF.registers\[3\]\[5\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__mux4_1
X_7043_ _3445_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8994_ clknet_leaf_93_CLK _0154_ VGND VGND VPWR VPWR RF.registers\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_124_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7945_ RF.registers\[18\]\[20\] _3497_ _3938_ VGND VGND VPWR VPWR _3939_ sky130_fd_sc_hd__mux2_1
X_7876_ _3879_ VGND VGND VPWR VPWR _3902_ sky130_fd_sc_hd__buf_4
X_6827_ RF.registers\[6\]\[23\] _3141_ _3326_ VGND VGND VPWR VPWR _3330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9546_ clknet_leaf_85_CLK _0706_ VGND VGND VPWR VPWR RF.registers\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6758_ _3071_ RF.registers\[14\]\[23\] _3289_ VGND VGND VPWR VPWR _3293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6689_ _3256_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__clkbuf_1
X_5709_ _2460_ _2461_ _2252_ VGND VGND VPWR VPWR _2462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9477_ clknet_leaf_63_CLK _0637_ VGND VGND VPWR VPWR RF.registers\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8428_ RF.registers\[12\]\[23\] _3504_ _4191_ VGND VGND VPWR VPWR _4195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8359_ _4158_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5991_ _1111_ _2335_ VGND VGND VPWR VPWR _2731_ sky130_fd_sc_hd__nor2_2
X_4942_ _1687_ _1695_ _1697_ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7730_ _3054_ RF.registers\[30\]\[15\] _3819_ VGND VGND VPWR VPWR _3825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7661_ _3788_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_1
X_9400_ clknet_leaf_38_CLK _0560_ VGND VGND VPWR VPWR RF.registers\[24\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_4873_ _1214_ _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__nand2_1
X_6612_ _3215_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7592_ _3052_ RF.registers\[28\]\[14\] _3747_ VGND VGND VPWR VPWR _3752_ sky130_fd_sc_hd__mux2_1
X_9331_ clknet_leaf_30_CLK _0491_ VGND VGND VPWR VPWR RF.registers\[21\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6543_ RF.registers\[0\]\[19\] _3132_ _3168_ VGND VGND VPWR VPWR _3178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6474_ _3138_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9262_ clknet_leaf_21_CLK _0422_ VGND VGND VPWR VPWR RF.registers\[23\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8213_ RF.registers\[1\]\[18\] _3493_ _4072_ VGND VGND VPWR VPWR _4081_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5425_ RF.registers\[28\]\[11\] RF.registers\[29\]\[11\] RF.registers\[30\]\[11\]
+ RF.registers\[31\]\[11\] _1675_ _1692_ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9193_ clknet_leaf_1_CLK _0353_ VGND VGND VPWR VPWR RF.registers\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8144_ _4044_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__clkbuf_1
X_5356_ _1712_ _2111_ VGND VGND VPWR VPWR _2112_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8075_ RF.registers\[20\]\[17\] _3491_ _4000_ VGND VGND VPWR VPWR _4008_ sky130_fd_sc_hd__mux2_1
X_5287_ RF.registers\[16\]\[3\] RF.registers\[17\]\[3\] RF.registers\[18\]\[3\] RF.registers\[19\]\[3\]
+ _1674_ _1691_ VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__mux4_1
X_4307_ RF.registers\[16\]\[5\] RF.registers\[17\]\[5\] RF.registers\[18\]\[5\] RF.registers\[19\]\[5\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__mux4_1
X_7026_ RF.registers\[3\]\[20\] _3134_ _3435_ VGND VGND VPWR VPWR _3436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8977_ clknet_leaf_19_CLK _0137_ VGND VGND VPWR VPWR RF.registers\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7928_ RF.registers\[18\]\[12\] _3481_ _3927_ VGND VGND VPWR VPWR _3930_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7859_ _3893_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9529_ clknet_leaf_34_CLK _0689_ VGND VGND VPWR VPWR RF.registers\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5210_ RF.registers\[28\]\[27\] RF.registers\[29\]\[27\] RF.registers\[30\]\[27\]
+ RF.registers\[31\]\[27\] _1767_ _1768_ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__mux4_1
XFILLER_0_122_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6190_ _2875_ _2885_ _2892_ _2904_ _2890_ VGND VGND VPWR VPWR _2919_ sky130_fd_sc_hd__o311a_1
X_5141_ _1693_ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_90_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5072_ _1716_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8900_ clknet_leaf_95_CLK _0060_ VGND VGND VPWR VPWR RF.registers\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8831_ clknet_leaf_66_CLK _1015_ VGND VGND VPWR VPWR RF.registers\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8762_ clknet_leaf_36_CLK _0946_ VGND VGND VPWR VPWR RF.registers\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5974_ _2707_ _2709_ _2715_ _2621_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__o22a_1
X_7713_ _3037_ RF.registers\[30\]\[7\] _3808_ VGND VGND VPWR VPWR _3816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8693_ clknet_leaf_29_CLK _0877_ VGND VGND VPWR VPWR RF.registers\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_4925_ _1680_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4856_ RF.registers\[0\]\[19\] RF.registers\[1\]\[19\] RF.registers\[2\]\[19\] RF.registers\[3\]\[19\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7644_ _3779_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7575_ _3035_ RF.registers\[28\]\[6\] _3736_ VGND VGND VPWR VPWR _3743_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9314_ clknet_leaf_91_CLK _0474_ VGND VGND VPWR VPWR RF.registers\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_4787_ RF.registers\[20\]\[10\] RF.registers\[21\]\[10\] RF.registers\[22\]\[10\]
+ RF.registers\[23\]\[10\] _1041_ _1043_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__mux4_1
X_6526_ _3169_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload80 clknet_leaf_53_CLK VGND VGND VPWR VPWR clkload80/Y sky130_fd_sc_hd__inv_6
X_9245_ clknet_leaf_15_CLK _0405_ VGND VGND VPWR VPWR RF.registers\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6457_ RF.registers\[17\]\[16\] _3126_ _3114_ VGND VGND VPWR VPWR _3127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6388_ net33 VGND VGND VPWR VPWR _3079_ sky130_fd_sc_hd__clkbuf_2
Xclkload91 clknet_leaf_36_CLK VGND VGND VPWR VPWR clkload91/Y sky130_fd_sc_hd__clkinvlp_4
X_9176_ clknet_leaf_39_CLK _0336_ VGND VGND VPWR VPWR RF.registers\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5408_ RF.registers\[16\]\[12\] RF.registers\[17\]\[12\] RF.registers\[18\]\[12\]
+ RF.registers\[19\]\[12\] _2113_ _2114_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__mux4_1
X_8127_ _4035_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__clkbuf_1
X_5339_ _2093_ _2094_ net3 VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__mux2_1
X_8058_ RF.registers\[20\]\[9\] _3474_ _3989_ VGND VGND VPWR VPWR _3999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7009_ RF.registers\[3\]\[12\] _3118_ _3424_ VGND VGND VPWR VPWR _3427_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5690_ _2442_ _2443_ _2252_ VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4710_ RF.registers\[16\]\[13\] RF.registers\[17\]\[13\] RF.registers\[18\]\[13\]
+ RF.registers\[19\]\[13\] _1027_ _1029_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4641_ _1395_ _1396_ _1040_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4572_ RF.registers\[12\]\[31\] RF.registers\[13\]\[31\] RF.registers\[14\]\[31\]
+ RF.registers\[15\]\[31\] _1324_ _1325_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7360_ _3629_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
X_7291_ _3592_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
X_6311_ net36 VGND VGND VPWR VPWR _3027_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6242_ _2498_ _2967_ _2327_ VGND VGND VPWR VPWR _2968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9030_ clknet_leaf_64_CLK _0190_ VGND VGND VPWR VPWR RF.registers\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6173_ _1298_ _2902_ VGND VGND VPWR VPWR _2903_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5124_ _1804_ _1878_ _1879_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5055_ _1807_ _1810_ _1697_ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8814_ clknet_leaf_56_CLK _0998_ VGND VGND VPWR VPWR RF.registers\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5957_ _2104_ _2699_ VGND VGND VPWR VPWR _2700_ sky130_fd_sc_hd__nand2_1
X_8745_ clknet_leaf_87_CLK _0929_ VGND VGND VPWR VPWR RF.registers\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4908_ net47 VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8676_ clknet_leaf_89_CLK _0860_ VGND VGND VPWR VPWR RF.registers\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7627_ _3087_ RF.registers\[28\]\[31\] _3735_ VGND VGND VPWR VPWR _3770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5888_ _2229_ _2597_ _2616_ _2246_ VGND VGND VPWR VPWR _2634_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4839_ _1593_ _1594_ _1287_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7558_ _3733_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
X_7489_ _3085_ RF.registers\[25\]\[30\] _3663_ VGND VGND VPWR VPWR _3697_ sky130_fd_sc_hd__mux2_1
X_6509_ _3160_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9228_ clknet_leaf_10_CLK _0388_ VGND VGND VPWR VPWR RF.registers\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_112_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9159_ clknet_leaf_59_CLK _0319_ VGND VGND VPWR VPWR RF.registers\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_6 _1754_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6860_ _3347_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5811_ _2286_ _2558_ VGND VGND VPWR VPWR _2560_ sky130_fd_sc_hd__or2_1
X_6791_ RF.registers\[6\]\[6\] _3105_ _3304_ VGND VGND VPWR VPWR _3311_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5742_ _2105_ _2491_ _2493_ VGND VGND VPWR VPWR _2494_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8530_ _4248_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5673_ _2424_ _2425_ _2426_ VGND VGND VPWR VPWR _2427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8461_ _4212_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__clkbuf_1
X_7412_ _3656_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__clkbuf_1
X_4624_ RF.registers\[8\]\[24\] RF.registers\[9\]\[24\] RF.registers\[10\]\[24\] RF.registers\[11\]\[24\]
+ _1351_ _1352_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8392_ RF.registers\[12\]\[6\] _3468_ _4169_ VGND VGND VPWR VPWR _4176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7343_ _3619_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
X_4555_ RF.registers\[4\]\[27\] RF.registers\[5\]\[27\] RF.registers\[6\]\[27\] RF.registers\[7\]\[27\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_633 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7274_ _3075_ RF.registers\[29\]\[25\] _3577_ VGND VGND VPWR VPWR _3583_ sky130_fd_sc_hd__mux2_1
X_9013_ clknet_leaf_25_CLK _0173_ VGND VGND VPWR VPWR RF.registers\[31\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4486_ _1240_ _1241_ _1211_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6225_ _1942_ _2950_ VGND VGND VPWR VPWR _2952_ sky130_fd_sc_hd__or2_1
X_6156_ _2875_ _2885_ VGND VGND VPWR VPWR _2887_ sky130_fd_sc_hd__or2_1
X_5107_ RF.registers\[16\]\[16\] RF.registers\[17\]\[16\] RF.registers\[18\]\[16\]
+ RF.registers\[19\]\[16\] _1705_ _1708_ VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6087_ _2753_ _2821_ _1126_ VGND VGND VPWR VPWR _2822_ sky130_fd_sc_hd__mux2_1
X_5038_ RF.registers\[4\]\[20\] RF.registers\[5\]\[20\] RF.registers\[6\]\[20\] RF.registers\[7\]\[20\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8728_ clknet_leaf_39_CLK _0912_ VGND VGND VPWR VPWR RF.registers\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6989_ _3416_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8659_ clknet_leaf_51_CLK _0843_ VGND VGND VPWR VPWR RF.registers\[0\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput65 net65 VGND VGND VPWR VPWR ALU_result[24] sky130_fd_sc_hd__buf_1
Xoutput54 net54 VGND VGND VPWR VPWR ALU_result[14] sky130_fd_sc_hd__buf_1
Xoutput76 net76 VGND VGND VPWR VPWR ALU_result[5] sky130_fd_sc_hd__buf_1
XFILLER_0_86_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4340_ RF.registers\[24\]\[3\] RF.registers\[25\]\[3\] RF.registers\[26\]\[3\] RF.registers\[27\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4271_ _1026_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6010_ _2744_ _2749_ VGND VGND VPWR VPWR _2750_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7961_ RF.registers\[18\]\[28\] _3446_ _3938_ VGND VGND VPWR VPWR _3947_ sky130_fd_sc_hd__mux2_1
X_7892_ _3910_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__clkbuf_1
X_6912_ _3374_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6843_ RF.registers\[6\]\[31\] _3017_ _3303_ VGND VGND VPWR VPWR _3338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9562_ clknet_leaf_35_CLK _0722_ VGND VGND VPWR VPWR RF.registers\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6774_ _3087_ RF.registers\[14\]\[31\] _3266_ VGND VGND VPWR VPWR _3301_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9493_ clknet_leaf_28_CLK _0653_ VGND VGND VPWR VPWR RF.registers\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_8513_ _4239_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5725_ _1125_ _1145_ _1167_ _2411_ VGND VGND VPWR VPWR _2478_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8444_ RF.registers\[12\]\[31\] net38 _4168_ VGND VGND VPWR VPWR _4203_ sky130_fd_sc_hd__mux2_1
X_5656_ _2409_ VGND VGND VPWR VPWR _2411_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4607_ RF.registers\[12\]\[25\] RF.registers\[13\]\[25\] RF.registers\[14\]\[25\]
+ RF.registers\[15\]\[25\] _1360_ _1361_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_98_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8375_ _4166_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__clkbuf_1
X_5587_ _1667_ _2124_ VGND VGND VPWR VPWR _2342_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4538_ RF.registers\[8\]\[26\] RF.registers\[9\]\[26\] RF.registers\[10\]\[26\] RF.registers\[11\]\[26\]
+ _1172_ _1279_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__mux4_1
X_7326_ _3610_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4469_ RF.registers\[28\]\[28\] RF.registers\[29\]\[28\] RF.registers\[30\]\[28\]
+ RF.registers\[31\]\[28\] _1220_ _1222_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__mux4_1
X_7257_ _3058_ RF.registers\[29\]\[17\] _3566_ VGND VGND VPWR VPWR _3574_ sky130_fd_sc_hd__mux2_1
X_6208_ _2893_ _2935_ VGND VGND VPWR VPWR _2936_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7188_ _3536_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
X_6139_ _1512_ _2835_ _1635_ _2658_ VGND VGND VPWR VPWR _2871_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_51_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5510_ _1699_ _2265_ VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__nand2_1
X_6490_ _3148_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5441_ _2195_ _2196_ _1711_ VGND VGND VPWR VPWR _2197_ sky130_fd_sc_hd__mux2_1
X_8160_ RF.registers\[24\]\[25\] _3508_ _4047_ VGND VGND VPWR VPWR _4053_ sky130_fd_sc_hd__mux2_1
X_5372_ RF.registers\[28\]\[14\] RF.registers\[29\]\[14\] RF.registers\[30\]\[14\]
+ RF.registers\[31\]\[14\] _1674_ _1691_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__mux4_1
X_8091_ _4016_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7111_ RF.registers\[19\]\[17\] _3491_ _3477_ VGND VGND VPWR VPWR _3492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4323_ RF.registers\[4\]\[5\] RF.registers\[5\]\[5\] RF.registers\[6\]\[5\] RF.registers\[7\]\[5\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__mux4_1
X_7042_ RF.registers\[3\]\[27\] _3444_ _3435_ VGND VGND VPWR VPWR _3445_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8993_ clknet_leaf_97_CLK _0153_ VGND VGND VPWR VPWR RF.registers\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7944_ _3915_ VGND VGND VPWR VPWR _3938_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7875_ _3901_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__clkbuf_1
X_6826_ _3329_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6757_ _3292_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9545_ clknet_leaf_88_CLK _0705_ VGND VGND VPWR VPWR RF.registers\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5708_ _2346_ _2351_ _2327_ VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__mux2_1
X_6688_ RF.registers\[8\]\[22\] _3139_ _3253_ VGND VGND VPWR VPWR _3256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9476_ clknet_leaf_95_CLK _0636_ VGND VGND VPWR VPWR RF.registers\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8427_ _4194_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__clkbuf_1
X_5639_ _1168_ _1755_ VGND VGND VPWR VPWR _2394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8358_ RF.registers\[16\]\[22\] _3502_ _4155_ VGND VGND VPWR VPWR _4158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7309_ _3601_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
X_8289_ _4121_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5990_ _2041_ _2102_ VGND VGND VPWR VPWR _2730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4941_ _1696_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4872_ _1626_ _1627_ _1189_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__mux2_1
X_7660_ RF.registers\[2\]\[14\] _3485_ _3783_ VGND VGND VPWR VPWR _3788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6611_ _3060_ RF.registers\[15\]\[18\] _3206_ VGND VGND VPWR VPWR _3215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9330_ clknet_leaf_41_CLK _0490_ VGND VGND VPWR VPWR RF.registers\[21\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7591_ _3751_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6542_ _3177_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_65_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_92_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6473_ RF.registers\[17\]\[21\] _3137_ _3135_ VGND VGND VPWR VPWR _3138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9261_ clknet_leaf_8_CLK _0421_ VGND VGND VPWR VPWR RF.registers\[23\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8212_ _4080_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__clkbuf_1
X_9192_ clknet_leaf_0_CLK _0352_ VGND VGND VPWR VPWR RF.registers\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5424_ RF.registers\[24\]\[11\] RF.registers\[25\]\[11\] RF.registers\[26\]\[11\]
+ RF.registers\[27\]\[11\] _1675_ _1692_ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8143_ RF.registers\[24\]\[17\] _3491_ _4036_ VGND VGND VPWR VPWR _4044_ sky130_fd_sc_hd__mux2_1
X_5355_ RF.registers\[8\]\[15\] RF.registers\[9\]\[15\] RF.registers\[10\]\[15\] RF.registers\[11\]\[15\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_7_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8074_ _4007_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4306_ RF.registers\[20\]\[5\] RF.registers\[21\]\[5\] RF.registers\[22\]\[5\] RF.registers\[23\]\[5\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__mux4_1
X_5286_ RF.registers\[20\]\[3\] RF.registers\[21\]\[3\] RF.registers\[22\]\[3\] RF.registers\[23\]\[3\]
+ _1674_ _1691_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7025_ _3412_ VGND VGND VPWR VPWR _3435_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_74_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8976_ clknet_leaf_6_CLK _0136_ VGND VGND VPWR VPWR RF.registers\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_7927_ _3929_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7858_ _3116_ RF.registers\[23\]\[11\] _3891_ VGND VGND VPWR VPWR _3893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6809_ _3320_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7789_ _3856_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9528_ clknet_leaf_39_CLK _0688_ VGND VGND VPWR VPWR RF.registers\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_83_CLK sky130_fd_sc_hd__clkbuf_8
X_9459_ clknet_leaf_30_CLK _0619_ VGND VGND VPWR VPWR RF.registers\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_74_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_12_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5140_ _1895_ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_90_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5071_ RF.registers\[20\]\[19\] RF.registers\[21\]\[19\] RF.registers\[22\]\[19\]
+ RF.registers\[23\]\[19\] _1676_ _1681_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8830_ clknet_leaf_67_CLK _1014_ VGND VGND VPWR VPWR RF.registers\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8761_ clknet_leaf_32_CLK _0945_ VGND VGND VPWR VPWR RF.registers\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5973_ _2712_ _2714_ VGND VGND VPWR VPWR _2715_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7712_ _3815_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4924_ _1679_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__buf_4
XFILLER_0_118_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8692_ clknet_leaf_43_CLK _0876_ VGND VGND VPWR VPWR RF.registers\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4855_ _1211_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7643_ RF.registers\[2\]\[6\] _3468_ _3772_ VGND VGND VPWR VPWR _3779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4786_ _1025_ _1533_ _1541_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__o21ai_2
X_7574_ _3742_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_65_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_65_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9313_ clknet_leaf_93_CLK _0473_ VGND VGND VPWR VPWR RF.registers\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6525_ RF.registers\[0\]\[10\] _3113_ _3168_ VGND VGND VPWR VPWR _3169_ sky130_fd_sc_hd__mux2_1
X_9244_ clknet_leaf_16_CLK _0404_ VGND VGND VPWR VPWR RF.registers\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload70 clknet_leaf_27_CLK VGND VGND VPWR VPWR clkload70/Y sky130_fd_sc_hd__bufinv_16
X_6456_ net21 VGND VGND VPWR VPWR _3126_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9175_ clknet_leaf_49_CLK _0335_ VGND VGND VPWR VPWR RF.registers\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload92 clknet_leaf_47_CLK VGND VGND VPWR VPWR clkload92/Y sky130_fd_sc_hd__clkinv_1
X_6387_ _3078_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__clkbuf_1
Xclkload81 clknet_leaf_54_CLK VGND VGND VPWR VPWR clkload81/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5407_ RF.registers\[28\]\[12\] RF.registers\[29\]\[12\] RF.registers\[30\]\[12\]
+ RF.registers\[31\]\[12\] _1703_ _1706_ VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__mux4_1
X_8126_ RF.registers\[24\]\[9\] _3474_ _4025_ VGND VGND VPWR VPWR _4035_ sky130_fd_sc_hd__mux2_1
X_5338_ RF.registers\[12\]\[1\] RF.registers\[13\]\[1\] RF.registers\[14\]\[1\] RF.registers\[15\]\[1\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _2094_ sky130_fd_sc_hd__mux4_1
X_8057_ _3998_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__clkbuf_1
X_5269_ RF.registers\[12\]\[24\] RF.registers\[13\]\[24\] RF.registers\[14\]\[24\]
+ RF.registers\[15\]\[24\] _1881_ _1883_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__mux4_1
X_7008_ _3426_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8959_ clknet_leaf_72_CLK _0119_ VGND VGND VPWR VPWR RF.registers\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_56_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_47_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_47_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4640_ RF.registers\[0\]\[6\] RF.registers\[1\]\[6\] RF.registers\[2\]\[6\] RF.registers\[3\]\[6\]
+ _1072_ _1073_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4571_ _1178_ _1326_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__and2_1
X_6310_ _3026_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7290_ _3019_ RF.registers\[31\]\[0\] _3591_ VGND VGND VPWR VPWR _3592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6241_ _2547_ VGND VGND VPWR VPWR _2967_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6172_ _1447_ _2901_ _2871_ _2741_ VGND VGND VPWR VPWR _2902_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5123_ _1126_ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5054_ _1808_ _1809_ _1739_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8813_ clknet_leaf_58_CLK _0997_ VGND VGND VPWR VPWR RF.registers\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5956_ _2610_ _2698_ _2251_ VGND VGND VPWR VPWR _2699_ sky130_fd_sc_hd__mux2_1
X_8744_ clknet_leaf_88_CLK _0928_ VGND VGND VPWR VPWR RF.registers\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5887_ _2210_ _2632_ VGND VGND VPWR VPWR _2633_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4907_ _1148_ _1662_ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__nand2_1
X_8675_ clknet_leaf_76_CLK _0859_ VGND VGND VPWR VPWR RF.registers\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_38_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_38_CLK sky130_fd_sc_hd__clkbuf_8
X_7626_ _3769_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__clkbuf_1
X_4838_ RF.registers\[12\]\[17\] RF.registers\[13\]\[17\] RF.registers\[14\]\[17\]
+ RF.registers\[15\]\[17\] _1191_ _1279_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_134_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7557_ _3085_ RF.registers\[27\]\[30\] _3699_ VGND VGND VPWR VPWR _3733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4769_ RF.registers\[0\]\[8\] RF.registers\[1\]\[8\] RF.registers\[2\]\[8\] RF.registers\[3\]\[8\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__mux4_1
X_7488_ _3696_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
X_6508_ RF.registers\[0\]\[2\] _3097_ _3157_ VGND VGND VPWR VPWR _3160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9227_ clknet_leaf_89_CLK _0387_ VGND VGND VPWR VPWR RF.registers\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6439_ RF.registers\[17\]\[10\] _3113_ _3114_ VGND VGND VPWR VPWR _3115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9158_ clknet_leaf_61_CLK _0318_ VGND VGND VPWR VPWR RF.registers\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_112_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8109_ _4026_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__clkbuf_1
X_9089_ clknet_leaf_97_CLK _0249_ VGND VGND VPWR VPWR RF.registers\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_29_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_7 _1811_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5810_ _2286_ _2558_ VGND VGND VPWR VPWR _2559_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6790_ _3310_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5741_ _2250_ _2255_ _2492_ _2373_ VGND VGND VPWR VPWR _2493_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8460_ RF.registers\[11\]\[6\] net42 _4205_ VGND VGND VPWR VPWR _4212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7411_ _3075_ RF.registers\[26\]\[25\] _3650_ VGND VGND VPWR VPWR _3656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5672_ _1879_ VGND VGND VPWR VPWR _2426_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4623_ _1214_ _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8391_ _4175_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__clkbuf_1
X_7342_ _3075_ RF.registers\[31\]\[25\] _3613_ VGND VGND VPWR VPWR _3619_ sky130_fd_sc_hd__mux2_1
X_4554_ _1254_ _1309_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7273_ _3582_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9012_ clknet_leaf_22_CLK _0172_ VGND VGND VPWR VPWR RF.registers\[31\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_4485_ RF.registers\[16\]\[20\] RF.registers\[17\]\[20\] RF.registers\[18\]\[20\]
+ RF.registers\[19\]\[20\] _1207_ _1208_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__mux4_1
X_6224_ _1942_ _2950_ VGND VGND VPWR VPWR _2951_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6155_ _2863_ _2870_ _2886_ _2408_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__o22a_1
XFILLER_0_0_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6086_ _2790_ _2820_ _1146_ VGND VGND VPWR VPWR _2821_ sky130_fd_sc_hd__mux2_1
X_5106_ RF.registers\[28\]\[16\] RF.registers\[29\]\[16\] RF.registers\[30\]\[16\]
+ RF.registers\[31\]\[16\] _1720_ _1723_ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__mux4_1
X_5037_ _1712_ _1792_ _1716_ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8727_ clknet_leaf_50_CLK _0911_ VGND VGND VPWR VPWR RF.registers\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6988_ RF.registers\[3\]\[2\] _3097_ _3413_ VGND VGND VPWR VPWR _3416_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5939_ _2504_ _2671_ _2682_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8658_ clknet_leaf_54_CLK _0842_ VGND VGND VPWR VPWR RF.registers\[0\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7609_ _3069_ RF.registers\[28\]\[22\] _3758_ VGND VGND VPWR VPWR _3761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8589_ clknet_leaf_8_CLK _0773_ VGND VGND VPWR VPWR RF.registers\[22\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput66 net66 VGND VGND VPWR VPWR ALU_result[25] sky130_fd_sc_hd__buf_1
Xoutput55 net55 VGND VGND VPWR VPWR ALU_result[15] sky130_fd_sc_hd__buf_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput77 net77 VGND VGND VPWR VPWR ALU_result[6] sky130_fd_sc_hd__buf_1
XFILLER_0_86_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4270_ A2[0] VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_9_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_9_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7960_ _3946_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__clkbuf_1
X_7891_ _3009_ RF.registers\[23\]\[27\] _3902_ VGND VGND VPWR VPWR _3910_ sky130_fd_sc_hd__mux2_1
X_6911_ RF.registers\[5\]\[31\] _3017_ _3339_ VGND VGND VPWR VPWR _3374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6842_ _3337_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9561_ clknet_leaf_30_CLK _0721_ VGND VGND VPWR VPWR RF.registers\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6773_ _3300_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9492_ clknet_leaf_17_CLK _0652_ VGND VGND VPWR VPWR RF.registers\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8512_ RF.registers\[11\]\[31\] net38 _4204_ VGND VGND VPWR VPWR _4239_ sky130_fd_sc_hd__mux2_1
X_5724_ _2468_ _2476_ VGND VGND VPWR VPWR _2477_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8443_ _4202_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__clkbuf_1
X_5655_ _1145_ _1166_ _2409_ VGND VGND VPWR VPWR _2410_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4606_ RF.registers\[8\]\[25\] RF.registers\[9\]\[25\] RF.registers\[10\]\[25\] RF.registers\[11\]\[25\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8374_ RF.registers\[16\]\[30\] _3450_ _4132_ VGND VGND VPWR VPWR _4166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5586_ _1758_ _1874_ _1839_ VGND VGND VPWR VPWR _2341_ sky130_fd_sc_hd__o21a_1
X_7325_ _3058_ RF.registers\[31\]\[17\] _3602_ VGND VGND VPWR VPWR _3610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4537_ _1198_ _1292_ _1071_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4468_ _1218_ _1223_ _1178_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__mux2_1
X_7256_ _3573_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6207_ _2904_ _2918_ VGND VGND VPWR VPWR _2935_ sky130_fd_sc_hd__nand2_1
X_7187_ RF.registers\[7\]\[17\] _3491_ _3528_ VGND VGND VPWR VPWR _3536_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _2504_ _2865_ _2869_ VGND VGND VPWR VPWR _2870_ sky130_fd_sc_hd__or3_1
X_4399_ RF.registers\[24\]\[0\] RF.registers\[25\]\[0\] RF.registers\[26\]\[0\] RF.registers\[27\]\[0\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_51_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _1256_ _2804_ VGND VGND VPWR VPWR _2805_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_3_4__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5440_ RF.registers\[28\]\[10\] RF.registers\[29\]\[10\] RF.registers\[30\]\[10\]
+ RF.registers\[31\]\[10\] _1674_ _1691_ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_112_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5371_ _2125_ _2126_ _2044_ VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__mux2_1
X_8090_ RF.registers\[20\]\[24\] _3506_ _4011_ VGND VGND VPWR VPWR _4016_ sky130_fd_sc_hd__mux2_1
X_7110_ net22 VGND VGND VPWR VPWR _3491_ sky130_fd_sc_hd__clkbuf_4
X_4322_ _1050_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__buf_6
X_7041_ net33 VGND VGND VPWR VPWR _3444_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_93_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8992_ clknet_leaf_69_CLK _0152_ VGND VGND VPWR VPWR RF.registers\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_121_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7943_ _3937_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_124_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7874_ _3132_ RF.registers\[23\]\[19\] _3891_ VGND VGND VPWR VPWR _3901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6825_ RF.registers\[6\]\[22\] _3139_ _3326_ VGND VGND VPWR VPWR _3329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6756_ _3069_ RF.registers\[14\]\[22\] _3289_ VGND VGND VPWR VPWR _3292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9544_ clknet_leaf_88_CLK _0704_ VGND VGND VPWR VPWR RF.registers\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5707_ _2402_ _2343_ _2327_ VGND VGND VPWR VPWR _2460_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6687_ _3255_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9475_ clknet_leaf_75_CLK _0635_ VGND VGND VPWR VPWR RF.registers\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_8426_ RF.registers\[12\]\[22\] _3502_ _4191_ VGND VGND VPWR VPWR _4194_ sky130_fd_sc_hd__mux2_1
X_5638_ _2391_ _2392_ VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__nor2_1
X_8357_ _4157_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__clkbuf_1
X_5569_ _1839_ _2324_ VGND VGND VPWR VPWR _2325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7308_ _3041_ RF.registers\[31\]\[9\] _3591_ VGND VGND VPWR VPWR _3601_ sky130_fd_sc_hd__mux2_1
X_8288_ _3137_ RF.registers\[13\]\[21\] _4119_ VGND VGND VPWR VPWR _4121_ sky130_fd_sc_hd__mux2_1
X_7239_ _3564_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4940_ net4 VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__clkbuf_8
X_4871_ RF.registers\[12\]\[18\] RF.registers\[13\]\[18\] RF.registers\[14\]\[18\]
+ RF.registers\[15\]\[18\] _1192_ _1195_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6610_ _3214_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7590_ _3050_ RF.registers\[28\]\[13\] _3747_ VGND VGND VPWR VPWR _3751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6541_ RF.registers\[0\]\[18\] _3130_ _3168_ VGND VGND VPWR VPWR _3177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6472_ net27 VGND VGND VPWR VPWR _3137_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_95_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9260_ clknet_leaf_3_CLK _0420_ VGND VGND VPWR VPWR RF.registers\[23\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5423_ _2143_ _2177_ _2178_ VGND VGND VPWR VPWR _2179_ sky130_fd_sc_hd__mux2_1
X_8211_ RF.registers\[1\]\[17\] _3491_ _4072_ VGND VGND VPWR VPWR _4080_ sky130_fd_sc_hd__mux2_1
X_9191_ clknet_leaf_58_CLK _0351_ VGND VGND VPWR VPWR RF.registers\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_8142_ _4043_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__clkbuf_1
X_5354_ _2106_ _2107_ _2108_ _2109_ _1685_ _1696_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__mux4_2
XFILLER_0_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4305_ A2[1] VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__buf_4
X_8073_ RF.registers\[20\]\[16\] _3489_ _4000_ VGND VGND VPWR VPWR _4007_ sky130_fd_sc_hd__mux2_1
X_5285_ _1880_ _2038_ _2040_ VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7024_ _3434_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8975_ clknet_leaf_6_CLK _0135_ VGND VGND VPWR VPWR RF.registers\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7926_ RF.registers\[18\]\[11\] _3479_ _3927_ VGND VGND VPWR VPWR _3929_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7857_ _3892_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__clkbuf_1
X_6808_ RF.registers\[6\]\[14\] _3122_ _3315_ VGND VGND VPWR VPWR _3320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7788_ RF.registers\[9\]\[10\] _3476_ _3855_ VGND VGND VPWR VPWR _3856_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9527_ clknet_leaf_49_CLK _0687_ VGND VGND VPWR VPWR RF.registers\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6739_ _3052_ RF.registers\[14\]\[14\] _3278_ VGND VGND VPWR VPWR _3283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9458_ clknet_leaf_43_CLK _0618_ VGND VGND VPWR VPWR RF.registers\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8409_ RF.registers\[12\]\[14\] _3485_ _4180_ VGND VGND VPWR VPWR _4185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9389_ clknet_leaf_4_CLK _0549_ VGND VGND VPWR VPWR RF.registers\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5070_ RF.registers\[16\]\[19\] RF.registers\[17\]\[19\] RF.registers\[18\]\[19\]
+ RF.registers\[19\]\[19\] _1676_ _1681_ VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8760_ clknet_leaf_38_CLK _0944_ VGND VGND VPWR VPWR RF.registers\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5972_ _2669_ _2689_ _2713_ VGND VGND VPWR VPWR _2714_ sky130_fd_sc_hd__o21ai_1
X_7711_ _3035_ RF.registers\[30\]\[6\] _3808_ VGND VGND VPWR VPWR _3815_ sky130_fd_sc_hd__mux2_1
X_4923_ _1678_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__buf_4
X_8691_ clknet_leaf_30_CLK _0875_ VGND VGND VPWR VPWR RF.registers\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4854_ RF.registers\[4\]\[19\] RF.registers\[5\]\[19\] RF.registers\[6\]\[19\] RF.registers\[7\]\[19\]
+ _1173_ _1175_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__mux4_1
X_7642_ _3778_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7573_ _3033_ RF.registers\[28\]\[5\] _3736_ VGND VGND VPWR VPWR _3742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4785_ _1535_ _1537_ _1540_ _1088_ net8 VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6524_ _3156_ VGND VGND VPWR VPWR _3168_ sky130_fd_sc_hd__buf_4
X_9312_ clknet_leaf_73_CLK _0472_ VGND VGND VPWR VPWR RF.registers\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9243_ clknet_leaf_45_CLK _0403_ VGND VGND VPWR VPWR RF.registers\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload71 clknet_leaf_28_CLK VGND VGND VPWR VPWR clkload71/Y sky130_fd_sc_hd__clkinv_4
Xclkload60 clknet_leaf_16_CLK VGND VGND VPWR VPWR clkload60/Y sky130_fd_sc_hd__clkinv_4
X_6455_ _3125_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9174_ clknet_leaf_48_CLK _0334_ VGND VGND VPWR VPWR RF.registers\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
Xclkload93 clknet_leaf_48_CLK VGND VGND VPWR VPWR clkload93/Y sky130_fd_sc_hd__clkinvlp_2
XTAP_TAPCELL_ROW_132_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6386_ _3077_ RF.registers\[22\]\[26\] _3065_ VGND VGND VPWR VPWR _3078_ sky130_fd_sc_hd__mux2_1
Xclkload82 clknet_leaf_55_CLK VGND VGND VPWR VPWR clkload82/Y sky130_fd_sc_hd__inv_8
X_5406_ RF.registers\[24\]\[12\] RF.registers\[25\]\[12\] RF.registers\[26\]\[12\]
+ RF.registers\[27\]\[12\] _2113_ _2114_ VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__mux4_1
X_5337_ RF.registers\[8\]\[1\] RF.registers\[9\]\[1\] RF.registers\[10\]\[1\] RF.registers\[11\]\[1\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__mux4_1
X_8125_ _4034_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__clkbuf_1
X_5268_ _2020_ _2023_ _1766_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__mux2_1
X_8056_ RF.registers\[20\]\[8\] _3472_ _3989_ VGND VGND VPWR VPWR _3998_ sky130_fd_sc_hd__mux2_1
X_7007_ RF.registers\[3\]\[11\] _3116_ _3424_ VGND VGND VPWR VPWR _3426_ sky130_fd_sc_hd__mux2_1
X_5199_ RF.registers\[12\]\[28\] RF.registers\[13\]\[28\] RF.registers\[14\]\[28\]
+ RF.registers\[15\]\[28\] _1896_ _1898_ VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8958_ clknet_leaf_68_CLK _0118_ VGND VGND VPWR VPWR RF.registers\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7909_ RF.registers\[18\]\[3\] _3462_ _3916_ VGND VGND VPWR VPWR _3920_ sky130_fd_sc_hd__mux2_1
X_8889_ clknet_leaf_49_CLK _0049_ VGND VGND VPWR VPWR RF.registers\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4570_ RF.registers\[8\]\[31\] RF.registers\[9\]\[31\] RF.registers\[10\]\[31\] RF.registers\[11\]\[31\]
+ _1324_ _1325_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6240_ _2442_ _2942_ VGND VGND VPWR VPWR _2966_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6171_ _1385_ VGND VGND VPWR VPWR _2901_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5122_ _1841_ _1876_ _1877_ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__mux2_1
X_5053_ RF.registers\[24\]\[18\] RF.registers\[25\]\[18\] RF.registers\[26\]\[18\]
+ RF.registers\[27\]\[18\] _1734_ _1735_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8812_ clknet_leaf_83_CLK _0996_ VGND VGND VPWR VPWR RF.registers\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5955_ _2649_ _2697_ _1803_ VGND VGND VPWR VPWR _2698_ sky130_fd_sc_hd__mux2_1
X_8743_ clknet_leaf_81_CLK _0927_ VGND VGND VPWR VPWR RF.registers\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4906_ _1169_ _1661_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__and2_1
X_5886_ _1558_ _2631_ VGND VGND VPWR VPWR _2632_ sky130_fd_sc_hd__xnor2_1
X_8674_ clknet_leaf_91_CLK _0858_ VGND VGND VPWR VPWR RF.registers\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7625_ _3085_ RF.registers\[28\]\[30\] _3735_ VGND VGND VPWR VPWR _3769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4837_ RF.registers\[8\]\[17\] RF.registers\[9\]\[17\] RF.registers\[10\]\[17\] RF.registers\[11\]\[17\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_134_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7556_ _3732_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
X_4768_ RF.registers\[4\]\[8\] RF.registers\[5\]\[8\] RF.registers\[6\]\[8\] RF.registers\[7\]\[8\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7487_ _3083_ RF.registers\[25\]\[29\] _3686_ VGND VGND VPWR VPWR _3696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4699_ _1451_ _1454_ _1071_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__mux2_1
X_6507_ _3159_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__clkbuf_1
X_6438_ _3092_ VGND VGND VPWR VPWR _3114_ sky130_fd_sc_hd__buf_4
X_9226_ clknet_leaf_85_CLK _0386_ VGND VGND VPWR VPWR RF.registers\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9157_ clknet_leaf_81_CLK _0317_ VGND VGND VPWR VPWR RF.registers\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_112_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6369_ _3066_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__clkbuf_1
X_8108_ RF.registers\[24\]\[0\] _3454_ _4025_ VGND VGND VPWR VPWR _4026_ sky130_fd_sc_hd__mux2_1
X_9088_ clknet_leaf_74_CLK _0248_ VGND VGND VPWR VPWR RF.registers\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8039_ _3988_ VGND VGND VPWR VPWR _3989_ sky130_fd_sc_hd__buf_6
XFILLER_0_98_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_8 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5740_ _2336_ _2328_ VGND VGND VPWR VPWR _2492_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7410_ _3655_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5671_ _2177_ _2213_ _2363_ VGND VGND VPWR VPWR _2425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4622_ _1376_ _1377_ _1199_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8390_ RF.registers\[12\]\[5\] _3466_ _4169_ VGND VGND VPWR VPWR _4175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7341_ _3618_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
X_4553_ _1307_ _1308_ _1199_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7272_ _3073_ RF.registers\[29\]\[24\] _3577_ VGND VGND VPWR VPWR _3582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4484_ RF.registers\[20\]\[20\] RF.registers\[21\]\[20\] RF.registers\[22\]\[20\]
+ RF.registers\[23\]\[20\] _1207_ _1208_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__mux4_1
X_9011_ clknet_leaf_25_CLK _0171_ VGND VGND VPWR VPWR RF.registers\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6223_ _1217_ _2949_ VGND VGND VPWR VPWR _2950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6154_ _2884_ _2885_ VGND VGND VPWR VPWR _2886_ sky130_fd_sc_hd__nor2_1
X_6085_ _2398_ _2395_ VGND VGND VPWR VPWR _2820_ sky130_fd_sc_hd__nor2_1
X_5105_ RF.registers\[24\]\[16\] RF.registers\[25\]\[16\] RF.registers\[26\]\[16\]
+ RF.registers\[27\]\[16\] _1705_ _1708_ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__mux4_1
X_5036_ RF.registers\[12\]\[20\] RF.registers\[13\]\[20\] RF.registers\[14\]\[20\]
+ RF.registers\[15\]\[20\] _1719_ _1722_ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6987_ _3415_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8726_ clknet_leaf_46_CLK _0910_ VGND VGND VPWR VPWR RF.registers\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_5938_ _1087_ _2678_ _2681_ VGND VGND VPWR VPWR _2682_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8657_ clknet_leaf_55_CLK _0841_ VGND VGND VPWR VPWR RF.registers\[0\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5869_ _1542_ _2615_ VGND VGND VPWR VPWR _2616_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7608_ _3760_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8588_ clknet_leaf_3_CLK _0772_ VGND VGND VPWR VPWR RF.registers\[22\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_7539_ _3067_ RF.registers\[27\]\[21\] _3722_ VGND VGND VPWR VPWR _3724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9209_ clknet_leaf_26_CLK _0369_ VGND VGND VPWR VPWR RF.registers\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_56_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput67 net67 VGND VGND VPWR VPWR ALU_result[26] sky130_fd_sc_hd__buf_1
Xoutput56 net56 VGND VGND VPWR VPWR ALU_result[16] sky130_fd_sc_hd__buf_1
XFILLER_0_31_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput78 net78 VGND VGND VPWR VPWR ALU_result[7] sky130_fd_sc_hd__buf_1
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7890_ _3909_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6910_ _3373_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__clkbuf_1
X_6841_ RF.registers\[6\]\[30\] _3015_ _3303_ VGND VGND VPWR VPWR _3337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9560_ clknet_leaf_39_CLK _0720_ VGND VGND VPWR VPWR RF.registers\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8511_ _4238_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__clkbuf_1
X_6772_ _3085_ RF.registers\[14\]\[30\] _3266_ VGND VGND VPWR VPWR _3300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9491_ clknet_leaf_27_CLK _0651_ VGND VGND VPWR VPWR RF.registers\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5723_ _2471_ _2475_ _2040_ VGND VGND VPWR VPWR _2476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8442_ RF.registers\[12\]\[30\] net37 _4168_ VGND VGND VPWR VPWR _4202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5654_ _1664_ net48 VGND VGND VPWR VPWR _2409_ sky130_fd_sc_hd__nor2_1
X_4605_ _1352_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__clkbuf_4
X_8373_ _4165_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7324_ _3609_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
X_5585_ _2178_ _2339_ VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4536_ RF.registers\[0\]\[26\] RF.registers\[1\]\[26\] RF.registers\[2\]\[26\] RF.registers\[3\]\[26\]
+ _1291_ _1194_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4467_ RF.registers\[16\]\[28\] RF.registers\[17\]\[28\] RF.registers\[18\]\[28\]
+ RF.registers\[19\]\[28\] _1220_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__mux4_1
X_7255_ _3056_ RF.registers\[29\]\[16\] _3566_ VGND VGND VPWR VPWR _3573_ sky130_fd_sc_hd__mux2_1
X_6206_ _2932_ _2933_ VGND VGND VPWR VPWR _2934_ sky130_fd_sc_hd__nor2_1
X_7186_ _3535_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_4398_ RF.registers\[28\]\[0\] RF.registers\[29\]\[0\] RF.registers\[30\]\[0\] RF.registers\[31\]\[0\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_129_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6137_ _2104_ _2736_ _2868_ _1086_ VGND VGND VPWR VPWR _2869_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_51_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _1512_ _1635_ _2658_ _2536_ VGND VGND VPWR VPWR _2804_ sky130_fd_sc_hd__a31o_1
X_5019_ RF.registers\[0\]\[21\] RF.registers\[1\]\[21\] RF.registers\[2\]\[21\] RF.registers\[3\]\[21\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8709_ clknet_leaf_59_CLK _0893_ VGND VGND VPWR VPWR RF.registers\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5370_ RF.registers\[16\]\[14\] RF.registers\[17\]\[14\] RF.registers\[18\]\[14\]
+ RF.registers\[19\]\[14\] _1674_ _1691_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4321_ _1071_ _1076_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__nand2_1
X_7040_ _3443_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8991_ clknet_leaf_72_CLK _0151_ VGND VGND VPWR VPWR RF.registers\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_7942_ RF.registers\[18\]\[19\] _3495_ _3927_ VGND VGND VPWR VPWR _3937_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7873_ _3900_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6824_ _3328_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6755_ _3291_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9543_ clknet_leaf_59_CLK _0703_ VGND VGND VPWR VPWR RF.registers\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5706_ _1128_ _2458_ _2421_ VGND VGND VPWR VPWR _2459_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9474_ clknet_leaf_76_CLK _0634_ VGND VGND VPWR VPWR RF.registers\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8425_ _4193_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__clkbuf_1
X_6686_ RF.registers\[8\]\[21\] _3137_ _3253_ VGND VGND VPWR VPWR _3255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5637_ _1799_ _1732_ VGND VGND VPWR VPWR _2392_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8356_ RF.registers\[16\]\[21\] _3500_ _4155_ VGND VGND VPWR VPWR _4157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5568_ _1842_ _2323_ VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4519_ _1273_ _1274_ _1211_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__mux2_1
X_8287_ _4120_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__clkbuf_1
X_7307_ _3600_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5499_ _2254_ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__buf_2
X_7238_ _3039_ RF.registers\[29\]\[8\] _3555_ VGND VGND VPWR VPWR _3564_ sky130_fd_sc_hd__mux2_1
X_7169_ _3526_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4870_ RF.registers\[8\]\[18\] RF.registers\[9\]\[18\] RF.registers\[10\]\[18\] RF.registers\[11\]\[18\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6540_ _3176_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6471_ _3136_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5422_ _1877_ VGND VGND VPWR VPWR _2178_ sky130_fd_sc_hd__clkbuf_4
X_8210_ _4079_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9190_ clknet_leaf_63_CLK _0350_ VGND VGND VPWR VPWR RF.registers\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8141_ RF.registers\[24\]\[16\] _3489_ _4036_ VGND VGND VPWR VPWR _4043_ sky130_fd_sc_hd__mux2_1
X_5353_ RF.registers\[24\]\[15\] RF.registers\[25\]\[15\] RF.registers\[26\]\[15\]
+ RF.registers\[27\]\[15\] _1782_ _1680_ VGND VGND VPWR VPWR _2109_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4304_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5284_ _2039_ VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__buf_2
X_8072_ _4006_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__clkbuf_1
X_7023_ RF.registers\[3\]\[19\] _3132_ _3424_ VGND VGND VPWR VPWR _3434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8974_ clknet_leaf_20_CLK _0134_ VGND VGND VPWR VPWR RF.registers\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7925_ _3928_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7856_ _3113_ RF.registers\[23\]\[10\] _3891_ VGND VGND VPWR VPWR _3892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6807_ _3319_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__clkbuf_1
X_9526_ clknet_leaf_47_CLK _0686_ VGND VGND VPWR VPWR RF.registers\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4999_ _1639_ _1754_ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__and2b_1
X_7787_ _3843_ VGND VGND VPWR VPWR _3855_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_137_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6738_ _3282_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9457_ clknet_leaf_13_CLK _0617_ VGND VGND VPWR VPWR RF.registers\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6669_ RF.registers\[8\]\[13\] _3120_ _3242_ VGND VGND VPWR VPWR _3246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8408_ _4184_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__clkbuf_1
X_9388_ clknet_leaf_3_CLK _0548_ VGND VGND VPWR VPWR RF.registers\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8339_ RF.registers\[16\]\[13\] _3483_ _4144_ VGND VGND VPWR VPWR _4148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5971_ _2661_ _2688_ _2687_ VGND VGND VPWR VPWR _2713_ sky130_fd_sc_hd__o21ba_1
X_8690_ clknet_leaf_43_CLK _0874_ VGND VGND VPWR VPWR RF.registers\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4922_ _1677_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__clkbuf_4
X_7710_ _3814_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7641_ RF.registers\[2\]\[5\] _3466_ _3772_ VGND VGND VPWR VPWR _3778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4853_ _1605_ _1608_ _1187_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7572_ _3741_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4784_ _1538_ _1539_ _1107_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9311_ clknet_leaf_71_CLK _0471_ VGND VGND VPWR VPWR RF.registers\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6523_ _3167_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_119_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9242_ clknet_leaf_35_CLK _0402_ VGND VGND VPWR VPWR RF.registers\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6454_ RF.registers\[17\]\[15\] _3124_ _3114_ VGND VGND VPWR VPWR _3125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload61 clknet_leaf_19_CLK VGND VGND VPWR VPWR clkload61/Y sky130_fd_sc_hd__inv_6
X_5405_ _2144_ _2160_ _1800_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_82_CLK VGND VGND VPWR VPWR clkload50/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_132_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9173_ clknet_leaf_44_CLK _0333_ VGND VGND VPWR VPWR RF.registers\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload72 clknet_leaf_37_CLK VGND VGND VPWR VPWR clkload72/Y sky130_fd_sc_hd__clkinv_4
X_6385_ net32 VGND VGND VPWR VPWR _3077_ sky130_fd_sc_hd__clkbuf_2
Xclkload83 clknet_leaf_56_CLK VGND VGND VPWR VPWR clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_0_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5336_ net3 _2091_ _1655_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__o21a_1
X_8124_ RF.registers\[24\]\[8\] _3472_ _4025_ VGND VGND VPWR VPWR _4034_ sky130_fd_sc_hd__mux2_1
X_5267_ _2021_ _2022_ _1745_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__mux2_1
X_8055_ _3997_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__clkbuf_1
X_7006_ _3425_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
X_5198_ RF.registers\[8\]\[28\] RF.registers\[9\]\[28\] RF.registers\[10\]\[28\] RF.registers\[11\]\[28\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__mux4_1
X_8957_ clknet_leaf_15_CLK _0117_ VGND VGND VPWR VPWR RF.registers\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7908_ _3919_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8888_ clknet_leaf_39_CLK _0048_ VGND VGND VPWR VPWR RF.registers\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7839_ _3097_ RF.registers\[23\]\[2\] _3880_ VGND VGND VPWR VPWR _3883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload0 clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9509_ clknet_leaf_80_CLK _0669_ VGND VGND VPWR VPWR RF.registers\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6170_ _2621_ _2894_ _2900_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__o21a_1
XFILLER_0_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5121_ _1145_ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5052_ RF.registers\[28\]\[18\] RF.registers\[29\]\[18\] RF.registers\[30\]\[18\]
+ RF.registers\[31\]\[18\] _1734_ _1735_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8811_ clknet_leaf_82_CLK _0995_ VGND VGND VPWR VPWR RF.registers\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8742_ clknet_leaf_59_CLK _0926_ VGND VGND VPWR VPWR RF.registers\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_5954_ _2345_ _2349_ VGND VGND VPWR VPWR _2697_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_101_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4905_ _1639_ _1660_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__nor2_1
X_5885_ _2630_ _1416_ _2593_ _2594_ _2595_ VGND VGND VPWR VPWR _2631_ sky130_fd_sc_hd__o41a_1
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8673_ clknet_leaf_95_CLK _0857_ VGND VGND VPWR VPWR RF.registers\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7624_ _3768_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__clkbuf_1
X_4836_ _1588_ _1589_ _1590_ _1591_ _1287_ _1078_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_134_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7555_ _3083_ RF.registers\[27\]\[29\] _3722_ VGND VGND VPWR VPWR _3732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6506_ RF.registers\[0\]\[1\] _3095_ _3157_ VGND VGND VPWR VPWR _3159_ sky130_fd_sc_hd__mux2_1
X_4767_ _1047_ _1522_ _1037_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7486_ _3695_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
X_4698_ _1452_ _1453_ _1036_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__mux2_1
X_6437_ net15 VGND VGND VPWR VPWR _3113_ sky130_fd_sc_hd__buf_2
X_9225_ clknet_leaf_87_CLK _0385_ VGND VGND VPWR VPWR RF.registers\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6368_ _3064_ RF.registers\[22\]\[20\] _3065_ VGND VGND VPWR VPWR _3066_ sky130_fd_sc_hd__mux2_1
X_9156_ clknet_leaf_90_CLK _0316_ VGND VGND VPWR VPWR RF.registers\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8107_ _4024_ VGND VGND VPWR VPWR _4025_ sky130_fd_sc_hd__buf_6
X_5319_ net3 _2074_ _1655_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__a21o_1
X_6299_ RF.registers\[10\]\[31\] _3017_ _3007_ VGND VGND VPWR VPWR _3018_ sky130_fd_sc_hd__mux2_1
X_9087_ clknet_leaf_73_CLK _0247_ VGND VGND VPWR VPWR RF.registers\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8038_ _3987_ _3155_ VGND VGND VPWR VPWR _3988_ sky130_fd_sc_hd__nor2_2
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 _1942_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5670_ _2423_ _2143_ _1147_ VGND VGND VPWR VPWR _2424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4621_ RF.registers\[0\]\[24\] RF.registers\[1\]\[24\] RF.registers\[2\]\[24\] RF.registers\[3\]\[24\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7340_ _3073_ RF.registers\[31\]\[24\] _3613_ VGND VGND VPWR VPWR _3618_ sky130_fd_sc_hd__mux2_1
X_4552_ RF.registers\[8\]\[27\] RF.registers\[9\]\[27\] RF.registers\[10\]\[27\] RF.registers\[11\]\[27\]
+ _1267_ _1268_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7271_ _3581_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
X_4483_ _1215_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6222_ _1237_ _2741_ _2930_ VGND VGND VPWR VPWR _2949_ sky130_fd_sc_hd__o21ba_1
X_9010_ clknet_leaf_42_CLK _0170_ VGND VGND VPWR VPWR RF.registers\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6153_ _2879_ _2883_ _2877_ VGND VGND VPWR VPWR _2885_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6084_ _2795_ _2798_ _2803_ _2819_ _2408_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__o32a_1
X_5104_ _1168_ _1859_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__or2_1
X_5035_ _1686_ _1790_ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6986_ RF.registers\[3\]\[1\] _3095_ _3413_ VGND VGND VPWR VPWR _3415_ sky130_fd_sc_hd__mux2_1
X_8725_ clknet_leaf_34_CLK _0909_ VGND VGND VPWR VPWR RF.registers\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_5937_ _2491_ _2591_ _2680_ VGND VGND VPWR VPWR _2681_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_0_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8656_ clknet_leaf_55_CLK _0840_ VGND VGND VPWR VPWR RF.registers\[0\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_7607_ _3067_ RF.registers\[28\]\[21\] _3758_ VGND VGND VPWR VPWR _3760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5868_ _1528_ _1416_ _2593_ _2594_ _2595_ VGND VGND VPWR VPWR _2615_ sky130_fd_sc_hd__o41a_1
X_4819_ RF.registers\[28\]\[16\] RF.registers\[29\]\[16\] RF.registers\[30\]\[16\]
+ RF.registers\[31\]\[16\] _1291_ _1174_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__mux4_1
X_5799_ _2546_ _2548_ _2501_ VGND VGND VPWR VPWR _2549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8587_ clknet_leaf_98_CLK _0771_ VGND VGND VPWR VPWR RF.registers\[22\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_7538_ _3723_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7469_ _3064_ RF.registers\[25\]\[20\] _3686_ VGND VGND VPWR VPWR _3687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9208_ clknet_leaf_38_CLK _0368_ VGND VGND VPWR VPWR RF.registers\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_56_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput57 net57 VGND VGND VPWR VPWR ALU_result[17] sky130_fd_sc_hd__buf_1
X_9139_ clknet_leaf_28_CLK _0299_ VGND VGND VPWR VPWR RF.registers\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xoutput68 net68 VGND VGND VPWR VPWR ALU_result[27] sky130_fd_sc_hd__buf_1
Xoutput79 net79 VGND VGND VPWR VPWR ALU_result[8] sky130_fd_sc_hd__buf_1
XFILLER_0_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6840_ _3336_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6771_ _3299_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8510_ RF.registers\[11\]\[30\] net37 _4204_ VGND VGND VPWR VPWR _4238_ sky130_fd_sc_hd__mux2_1
X_5722_ _2472_ _2474_ _2251_ VGND VGND VPWR VPWR _2475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9490_ clknet_leaf_42_CLK _0650_ VGND VGND VPWR VPWR RF.registers\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8441_ _4201_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__clkbuf_1
X_5653_ _2333_ VGND VGND VPWR VPWR _2408_ sky130_fd_sc_hd__buf_2
XFILLER_0_33_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4604_ _1351_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__buf_4
X_8372_ RF.registers\[16\]\[29\] _3448_ _4155_ VGND VGND VPWR VPWR _4165_ sky130_fd_sc_hd__mux2_1
X_5584_ _1799_ _2098_ _2338_ VGND VGND VPWR VPWR _2339_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7323_ _3056_ RF.registers\[31\]\[16\] _3602_ VGND VGND VPWR VPWR _3609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4535_ _1290_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4466_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__clkbuf_4
X_7254_ _3572_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6205_ _1958_ _2931_ VGND VGND VPWR VPWR _2933_ sky130_fd_sc_hd__and2_1
X_7185_ RF.registers\[7\]\[16\] _3489_ _3528_ VGND VGND VPWR VPWR _3535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4397_ _1088_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6136_ _2254_ _2801_ _2867_ _2336_ VGND VGND VPWR VPWR _2868_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6067_ _2799_ _2731_ _2802_ _2496_ VGND VGND VPWR VPWR _2803_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5018_ RF.registers\[4\]\[21\] RF.registers\[5\]\[21\] RF.registers\[6\]\[21\] RF.registers\[7\]\[21\]
+ _1705_ _1708_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6969_ RF.registers\[4\]\[26\] _3002_ _3398_ VGND VGND VPWR VPWR _3405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8708_ clknet_leaf_90_CLK _0892_ VGND VGND VPWR VPWR RF.registers\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8639_ clknet_leaf_66_CLK _0823_ VGND VGND VPWR VPWR RF.registers\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4320_ _1074_ _1075_ _1048_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8990_ clknet_leaf_69_CLK _0150_ VGND VGND VPWR VPWR RF.registers\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7941_ _3936_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7872_ _3130_ RF.registers\[23\]\[18\] _3891_ VGND VGND VPWR VPWR _3900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6823_ RF.registers\[6\]\[21\] _3137_ _3326_ VGND VGND VPWR VPWR _3328_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6754_ _3067_ RF.registers\[14\]\[21\] _3289_ VGND VGND VPWR VPWR _3291_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_95_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_95_CLK sky130_fd_sc_hd__clkbuf_8
X_9542_ clknet_leaf_60_CLK _0702_ VGND VGND VPWR VPWR RF.registers\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6685_ _3254_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5705_ _2455_ _2457_ _1146_ VGND VGND VPWR VPWR _2458_ sky130_fd_sc_hd__mux2_1
X_9473_ clknet_leaf_93_CLK _0633_ VGND VGND VPWR VPWR RF.registers\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8424_ RF.registers\[12\]\[21\] _3500_ _4191_ VGND VGND VPWR VPWR _4193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5636_ _1667_ _2034_ VGND VGND VPWR VPWR _2391_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8355_ _4156_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5567_ _1728_ _2314_ _2318_ _2322_ VGND VGND VPWR VPWR _2323_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4518_ RF.registers\[0\]\[21\] RF.registers\[1\]\[21\] RF.registers\[2\]\[21\] RF.registers\[3\]\[21\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__mux4_1
X_8286_ _3134_ RF.registers\[13\]\[20\] _4119_ VGND VGND VPWR VPWR _4120_ sky130_fd_sc_hd__mux2_1
X_5498_ _2039_ _1126_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__or2_2
X_7306_ _3039_ RF.registers\[31\]\[8\] _3591_ VGND VGND VPWR VPWR _3600_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4449_ _1078_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__buf_4
X_7237_ _3563_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7168_ RF.registers\[7\]\[8\] _3472_ _3517_ VGND VGND VPWR VPWR _3526_ sky130_fd_sc_hd__mux2_1
X_6119_ _1446_ _2741_ _2836_ VGND VGND VPWR VPWR _2852_ sky130_fd_sc_hd__o21ai_1
X_7099_ RF.registers\[19\]\[13\] _3483_ _3477_ VGND VGND VPWR VPWR _3484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_86_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_86_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_40_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_10_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_77_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_77_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6470_ RF.registers\[17\]\[20\] _3134_ _3135_ VGND VGND VPWR VPWR _3136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5421_ _2161_ _2176_ VGND VGND VPWR VPWR _2177_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8140_ _4042_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__clkbuf_1
X_5352_ RF.registers\[28\]\[15\] RF.registers\[29\]\[15\] RF.registers\[30\]\[15\]
+ RF.registers\[31\]\[15\] _1782_ _1680_ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8071_ RF.registers\[20\]\[15\] _3487_ _4000_ VGND VGND VPWR VPWR _4006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4303_ _1025_ _1039_ _1058_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__o21ai_2
X_7022_ _3433_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
X_5283_ _1171_ _1094_ _1098_ _1102_ _1109_ VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8973_ clknet_leaf_2_CLK _0133_ VGND VGND VPWR VPWR RF.registers\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_7924_ RF.registers\[18\]\[10\] _3476_ _3927_ VGND VGND VPWR VPWR _3928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7855_ _3879_ VGND VGND VPWR VPWR _3891_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_68_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_68_CLK sky130_fd_sc_hd__clkbuf_8
X_6806_ RF.registers\[6\]\[13\] _3120_ _3315_ VGND VGND VPWR VPWR _3319_ sky130_fd_sc_hd__mux2_1
X_9525_ clknet_leaf_36_CLK _0685_ VGND VGND VPWR VPWR RF.registers\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_4998_ _1671_ _1744_ _1749_ _1753_ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__o22a_1
X_7786_ _3854_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6737_ _3050_ RF.registers\[14\]\[13\] _3278_ VGND VGND VPWR VPWR _3282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9456_ clknet_leaf_13_CLK _0616_ VGND VGND VPWR VPWR RF.registers\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6668_ _3245_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5619_ _2255_ _2364_ _2371_ _2373_ VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__o211a_1
X_9387_ clknet_leaf_0_CLK _0547_ VGND VGND VPWR VPWR RF.registers\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8407_ RF.registers\[12\]\[13\] _3483_ _4180_ VGND VGND VPWR VPWR _4184_ sky130_fd_sc_hd__mux2_1
X_6599_ _3048_ RF.registers\[15\]\[12\] _3206_ VGND VGND VPWR VPWR _3209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8338_ _4147_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8269_ _3118_ RF.registers\[13\]\[12\] _4108_ VGND VGND VPWR VPWR _4111_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_61_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_59_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_59_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5970_ _2140_ _2711_ VGND VGND VPWR VPWR _2712_ sky130_fd_sc_hd__xnor2_1
X_4921_ net2 VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4852_ _1606_ _1607_ _1178_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__mux2_1
X_7640_ _3777_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7571_ _3031_ RF.registers\[28\]\[4\] _3736_ VGND VGND VPWR VPWR _3741_ sky130_fd_sc_hd__mux2_1
X_4783_ RF.registers\[0\]\[9\] RF.registers\[1\]\[9\] RF.registers\[2\]\[9\] RF.registers\[3\]\[9\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9310_ clknet_leaf_68_CLK _0470_ VGND VGND VPWR VPWR RF.registers\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6522_ RF.registers\[0\]\[9\] _3111_ _3157_ VGND VGND VPWR VPWR _3167_ sky130_fd_sc_hd__mux2_1
X_9241_ clknet_leaf_34_CLK _0401_ VGND VGND VPWR VPWR RF.registers\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6453_ net20 VGND VGND VPWR VPWR _3124_ sky130_fd_sc_hd__buf_2
XFILLER_0_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9172_ clknet_leaf_44_CLK _0332_ VGND VGND VPWR VPWR RF.registers\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xclkload62 clknet_leaf_20_CLK VGND VGND VPWR VPWR clkload62/Y sky130_fd_sc_hd__inv_8
Xclkload51 clknet_leaf_83_CLK VGND VGND VPWR VPWR clkload51/Y sky130_fd_sc_hd__clkinv_4
X_5404_ _1640_ _2151_ _2159_ VGND VGND VPWR VPWR _2160_ sky130_fd_sc_hd__o21a_2
Xclkload40 clknet_leaf_78_CLK VGND VGND VPWR VPWR clkload40/Y sky130_fd_sc_hd__clkinvlp_2
X_6384_ _3076_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_132_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload84 clknet_leaf_29_CLK VGND VGND VPWR VPWR clkload84/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_113_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload73 clknet_leaf_40_CLK VGND VGND VPWR VPWR clkload73/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8123_ _4033_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__clkbuf_1
X_5335_ RF.registers\[0\]\[1\] RF.registers\[1\]\[1\] RF.registers\[2\]\[1\] RF.registers\[3\]\[1\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2091_ sky130_fd_sc_hd__mux4_1
X_5266_ RF.registers\[24\]\[24\] RF.registers\[25\]\[24\] RF.registers\[26\]\[24\]
+ RF.registers\[27\]\[24\] _1918_ _1919_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8054_ RF.registers\[20\]\[7\] _3470_ _3989_ VGND VGND VPWR VPWR _3997_ sky130_fd_sc_hd__mux2_1
X_7005_ RF.registers\[3\]\[10\] _3113_ _3424_ VGND VGND VPWR VPWR _3425_ sky130_fd_sc_hd__mux2_1
X_5197_ _1901_ _1952_ _1766_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__a21o_1
X_8956_ clknet_leaf_37_CLK _0116_ VGND VGND VPWR VPWR RF.registers\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7907_ RF.registers\[18\]\[2\] _3460_ _3916_ VGND VGND VPWR VPWR _3919_ sky130_fd_sc_hd__mux2_1
X_8887_ clknet_leaf_49_CLK _0047_ VGND VGND VPWR VPWR RF.registers\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7838_ _3882_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7769_ RF.registers\[9\]\[1\] _3458_ _3844_ VGND VGND VPWR VPWR _3846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9508_ clknet_leaf_89_CLK _0668_ VGND VGND VPWR VPWR RF.registers\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload1 clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_8
XFILLER_0_116_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9439_ clknet_leaf_65_CLK _0599_ VGND VGND VPWR VPWR RF.registers\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5120_ _1860_ _1875_ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__nand2_1
X_5051_ _1805_ _1806_ _1739_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8810_ clknet_leaf_83_CLK _0994_ VGND VGND VPWR VPWR RF.registers\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8741_ clknet_leaf_80_CLK _0925_ VGND VGND VPWR VPWR RF.registers\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5953_ _2340_ _2608_ _1879_ VGND VGND VPWR VPWR _2696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5884_ _1528_ _1542_ VGND VGND VPWR VPWR _2630_ sky130_fd_sc_hd__or2b_1
X_8672_ clknet_leaf_73_CLK _0856_ VGND VGND VPWR VPWR RF.registers\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_4904_ _1640_ _1650_ _1654_ _1659_ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7623_ _3083_ RF.registers\[28\]\[29\] _3758_ VGND VGND VPWR VPWR _3768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4835_ RF.registers\[20\]\[17\] RF.registers\[21\]\[17\] RF.registers\[22\]\[17\]
+ RF.registers\[23\]\[17\] _1291_ _1194_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7554_ _3731_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4766_ RF.registers\[8\]\[8\] RF.registers\[9\]\[8\] RF.registers\[10\]\[8\] RF.registers\[11\]\[8\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6505_ _3158_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__clkbuf_1
X_7485_ _3081_ RF.registers\[25\]\[28\] _3686_ VGND VGND VPWR VPWR _3695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4697_ RF.registers\[24\]\[12\] RF.registers\[25\]\[12\] RF.registers\[26\]\[12\]
+ RF.registers\[27\]\[12\] _1219_ _1221_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6436_ _3112_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9224_ clknet_leaf_88_CLK _0384_ VGND VGND VPWR VPWR RF.registers\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6367_ _3022_ VGND VGND VPWR VPWR _3065_ sky130_fd_sc_hd__buf_4
X_9155_ clknet_leaf_75_CLK _0315_ VGND VGND VPWR VPWR RF.registers\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8106_ _3155_ _3626_ VGND VGND VPWR VPWR _4024_ sky130_fd_sc_hd__nor2b_4
X_5318_ RF.registers\[12\]\[2\] RF.registers\[13\]\[2\] RF.registers\[14\]\[2\] RF.registers\[15\]\[2\]
+ _1673_ _1690_ VGND VGND VPWR VPWR _2074_ sky130_fd_sc_hd__mux4_1
X_6298_ net38 VGND VGND VPWR VPWR _3017_ sky130_fd_sc_hd__buf_2
X_9086_ clknet_leaf_69_CLK _0246_ VGND VGND VPWR VPWR RF.registers\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_5249_ _2003_ _2004_ _1726_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__mux2_1
X_8037_ _3021_ VGND VGND VPWR VPWR _3987_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8939_ clknet_leaf_90_CLK _0099_ VGND VGND VPWR VPWR RF.registers\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4620_ RF.registers\[4\]\[24\] RF.registers\[5\]\[24\] RF.registers\[6\]\[24\] RF.registers\[7\]\[24\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4551_ RF.registers\[12\]\[27\] RF.registers\[13\]\[27\] RF.registers\[14\]\[27\]
+ RF.registers\[15\]\[27\] _1267_ _1268_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_116_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7270_ _3071_ RF.registers\[29\]\[23\] _3577_ VGND VGND VPWR VPWR _3581_ sky130_fd_sc_hd__mux2_1
X_4482_ _1217_ _1237_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nand2_1
X_6221_ _2421_ _2941_ _2943_ _2948_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__o22a_1
X_6152_ _2877_ _2879_ _2883_ VGND VGND VPWR VPWR _2884_ sky130_fd_sc_hd__and3_1
X_5103_ _1842_ _1858_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_111_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _2808_ _2818_ VGND VGND VPWR VPWR _2819_ sky130_fd_sc_hd__xnor2_1
X_5034_ RF.registers\[8\]\[20\] RF.registers\[9\]\[20\] RF.registers\[10\]\[20\] RF.registers\[11\]\[20\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_127_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6985_ _3414_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
X_8724_ clknet_leaf_44_CLK _0908_ VGND VGND VPWR VPWR RF.registers\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5936_ _2486_ _2588_ _2679_ _1962_ _2333_ VGND VGND VPWR VPWR _2680_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8655_ clknet_leaf_57_CLK _0839_ VGND VGND VPWR VPWR RF.registers\[0\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7606_ _3759_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__clkbuf_1
X_5867_ _1087_ _2613_ VGND VGND VPWR VPWR _2614_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4818_ RF.registers\[24\]\[16\] RF.registers\[25\]\[16\] RF.registers\[26\]\[16\]
+ RF.registers\[27\]\[16\] _1291_ _1194_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__mux4_1
X_5798_ _2499_ _2547_ _2347_ VGND VGND VPWR VPWR _2548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8586_ clknet_leaf_9_CLK _0770_ VGND VGND VPWR VPWR RF.registers\[22\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7537_ _3064_ RF.registers\[27\]\[20\] _3722_ VGND VGND VPWR VPWR _3723_ sky130_fd_sc_hd__mux2_1
X_4749_ _1503_ _1504_ _1190_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7468_ _3663_ VGND VGND VPWR VPWR _3686_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9207_ clknet_leaf_31_CLK _0367_ VGND VGND VPWR VPWR RF.registers\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6419_ net40 VGND VGND VPWR VPWR _3101_ sky130_fd_sc_hd__buf_2
Xoutput58 net58 VGND VGND VPWR VPWR ALU_result[18] sky130_fd_sc_hd__buf_1
X_7399_ _3649_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__clkbuf_1
X_9138_ clknet_leaf_42_CLK _0298_ VGND VGND VPWR VPWR RF.registers\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xoutput69 net69 VGND VGND VPWR VPWR ALU_result[28] sky130_fd_sc_hd__buf_1
X_9069_ clknet_leaf_3_CLK _0229_ VGND VGND VPWR VPWR RF.registers\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6770_ _3083_ RF.registers\[14\]\[29\] _3289_ VGND VGND VPWR VPWR _3299_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5721_ _2473_ _2385_ _1146_ VGND VGND VPWR VPWR _2474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8440_ RF.registers\[12\]\[29\] net35 _4191_ VGND VGND VPWR VPWR _4201_ sky130_fd_sc_hd__mux2_1
X_5652_ _1666_ _2406_ VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__or2_1
X_4603_ _1355_ _1358_ _1214_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__mux2_1
X_8371_ _4164_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__clkbuf_1
X_5583_ _1167_ _1661_ VGND VGND VPWR VPWR _2338_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7322_ _3608_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
X_4534_ _1065_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7253_ _3054_ RF.registers\[29\]\[15\] _3566_ VGND VGND VPWR VPWR _3572_ sky130_fd_sc_hd__mux2_1
X_4465_ _1053_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6204_ _1958_ _2931_ VGND VGND VPWR VPWR _2932_ sky130_fd_sc_hd__nor2_1
X_7184_ _3534_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
X_4396_ _1150_ _1151_ _1035_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _2847_ _2866_ _1147_ VGND VGND VPWR VPWR _2867_ sky130_fd_sc_hd__mux2_1
X_6066_ _2735_ _2801_ _2252_ VGND VGND VPWR VPWR _2802_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _1717_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6968_ _3404_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8707_ clknet_leaf_78_CLK _0891_ VGND VGND VPWR VPWR RF.registers\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6899_ RF.registers\[5\]\[25\] _3145_ _3362_ VGND VGND VPWR VPWR _3368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5919_ _2661_ _2662_ VGND VGND VPWR VPWR _2663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8638_ clknet_leaf_67_CLK _0822_ VGND VGND VPWR VPWR RF.registers\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8569_ clknet_leaf_34_CLK _0753_ VGND VGND VPWR VPWR RF.registers\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7940_ RF.registers\[18\]\[18\] _3493_ _3927_ VGND VGND VPWR VPWR _3936_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7871_ _3899_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6822_ _3327_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6753_ _3290_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9541_ clknet_leaf_80_CLK _0701_ VGND VGND VPWR VPWR RF.registers\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6684_ RF.registers\[8\]\[20\] _3134_ _3253_ VGND VGND VPWR VPWR _3254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5704_ _2456_ VGND VGND VPWR VPWR _2457_ sky130_fd_sc_hd__inv_2
X_9472_ clknet_leaf_70_CLK _0632_ VGND VGND VPWR VPWR RF.registers\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8423_ _4192_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__clkbuf_1
X_5635_ _2382_ _2389_ _2251_ VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8354_ RF.registers\[16\]\[20\] _3497_ _4155_ VGND VGND VPWR VPWR _4156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5566_ _1696_ _2321_ _1670_ VGND VGND VPWR VPWR _2322_ sky130_fd_sc_hd__o21ai_1
X_4517_ RF.registers\[4\]\[21\] RF.registers\[5\]\[21\] RF.registers\[6\]\[21\] RF.registers\[7\]\[21\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__mux4_1
X_8285_ _4096_ VGND VGND VPWR VPWR _4119_ sky130_fd_sc_hd__buf_4
X_5497_ _2179_ _2250_ _2252_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__mux2_1
X_7305_ _3599_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
X_4448_ RF.registers\[8\]\[29\] RF.registers\[9\]\[29\] RF.registers\[10\]\[29\] RF.registers\[11\]\[29\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7236_ _3037_ RF.registers\[29\]\[7\] _3555_ VGND VGND VPWR VPWR _3563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4379_ _1131_ _1134_ _1037_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__mux2_1
X_7167_ _3525_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_6118_ _2408_ _2845_ _2846_ _2851_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__o22a_1
X_7098_ net18 VGND VGND VPWR VPWR _3483_ sky130_fd_sc_hd__buf_2
X_6049_ _1820_ _2768_ VGND VGND VPWR VPWR _2786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5420_ _1758_ _2175_ _1800_ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5351_ RF.registers\[16\]\[15\] RF.registers\[17\]\[15\] RF.registers\[18\]\[15\]
+ RF.registers\[19\]\[15\] _1782_ _1680_ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5282_ _1962_ _2037_ _1879_ VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4302_ _1046_ _1051_ _1056_ _1038_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8070_ _4005_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__clkbuf_1
X_7021_ RF.registers\[3\]\[18\] _3130_ _3424_ VGND VGND VPWR VPWR _3433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8972_ clknet_leaf_2_CLK _0132_ VGND VGND VPWR VPWR RF.registers\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7923_ _3915_ VGND VGND VPWR VPWR _3927_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7854_ _3890_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6805_ _3318_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__clkbuf_1
X_7785_ RF.registers\[9\]\[9\] _3474_ _3844_ VGND VGND VPWR VPWR _3854_ sky130_fd_sc_hd__mux2_1
X_4997_ _1717_ _1752_ _1729_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__a21o_1
X_9524_ clknet_leaf_44_CLK _0684_ VGND VGND VPWR VPWR RF.registers\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6736_ _3281_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_137_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9455_ clknet_leaf_11_CLK _0615_ VGND VGND VPWR VPWR RF.registers\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6667_ RF.registers\[8\]\[12\] _3118_ _3242_ VGND VGND VPWR VPWR _3245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5618_ _2372_ VGND VGND VPWR VPWR _2373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9386_ clknet_leaf_8_CLK _0546_ VGND VGND VPWR VPWR RF.registers\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6598_ _3208_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__clkbuf_1
X_8406_ _4183_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__clkbuf_1
X_8337_ RF.registers\[16\]\[12\] _3481_ _4144_ VGND VGND VPWR VPWR _4147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5549_ _1728_ _2296_ _2300_ _2304_ VGND VGND VPWR VPWR _2305_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_112_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8268_ _4110_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__clkbuf_1
X_7219_ net13 net12 net11 VGND VGND VPWR VPWR _3553_ sky130_fd_sc_hd__and3_4
X_8199_ RF.registers\[1\]\[11\] _3479_ _4072_ VGND VGND VPWR VPWR _4074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _1675_ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4851_ RF.registers\[24\]\[19\] RF.registers\[25\]\[19\] RF.registers\[26\]\[19\]
+ RF.registers\[27\]\[19\] _1220_ _1222_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_103_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4782_ RF.registers\[4\]\[9\] RF.registers\[5\]\[9\] RF.registers\[6\]\[9\] RF.registers\[7\]\[9\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__mux4_1
X_7570_ _3740_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6521_ _3166_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_119_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9240_ clknet_leaf_39_CLK _0400_ VGND VGND VPWR VPWR RF.registers\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6452_ _3123_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__clkbuf_1
X_9171_ clknet_leaf_50_CLK _0331_ VGND VGND VPWR VPWR RF.registers\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xclkload52 clknet_leaf_5_CLK VGND VGND VPWR VPWR clkload52/Y sky130_fd_sc_hd__clkinv_4
Xclkload30 clknet_leaf_67_CLK VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__clkinvlp_2
X_5403_ _2153_ _2155_ _2158_ net4 net5 VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__a221o_1
Xclkload41 clknet_leaf_79_CLK VGND VGND VPWR VPWR clkload41/Y sky130_fd_sc_hd__inv_6
X_6383_ _3075_ RF.registers\[22\]\[25\] _3065_ VGND VGND VPWR VPWR _3076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload85 clknet_leaf_30_CLK VGND VGND VPWR VPWR clkload85/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload74 clknet_leaf_41_CLK VGND VGND VPWR VPWR clkload74/Y sky130_fd_sc_hd__inv_6
Xclkload63 clknet_leaf_21_CLK VGND VGND VPWR VPWR clkload63/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8122_ RF.registers\[24\]\[7\] _3470_ _4025_ VGND VGND VPWR VPWR _4033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5334_ _1645_ _2089_ VGND VGND VPWR VPWR _2090_ sky130_fd_sc_hd__or2_1
X_5265_ RF.registers\[28\]\[24\] RF.registers\[29\]\[24\] RF.registers\[30\]\[24\]
+ RF.registers\[31\]\[24\] _1918_ _1919_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__mux4_1
X_8053_ _3996_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__clkbuf_1
X_5196_ RF.registers\[0\]\[28\] RF.registers\[1\]\[28\] RF.registers\[2\]\[28\] RF.registers\[3\]\[28\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__mux4_1
X_7004_ _3412_ VGND VGND VPWR VPWR _3424_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8955_ clknet_leaf_45_CLK _0115_ VGND VGND VPWR VPWR RF.registers\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_48_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8886_ clknet_leaf_48_CLK _0046_ VGND VGND VPWR VPWR RF.registers\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7906_ _3918_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7837_ _3095_ RF.registers\[23\]\[1\] _3880_ VGND VGND VPWR VPWR _3882_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7768_ _3845_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6719_ _3272_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__clkbuf_1
X_7699_ _3019_ RF.registers\[30\]\[0\] _3808_ VGND VGND VPWR VPWR _3809_ sky130_fd_sc_hd__mux2_1
X_9507_ clknet_leaf_77_CLK _0667_ VGND VGND VPWR VPWR RF.registers\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload2 clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9438_ clknet_leaf_67_CLK _0598_ VGND VGND VPWR VPWR RF.registers\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9369_ clknet_leaf_31_CLK _0529_ VGND VGND VPWR VPWR RF.registers\[20\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5050_ RF.registers\[16\]\[18\] RF.registers\[17\]\[18\] RF.registers\[18\]\[18\]
+ RF.registers\[19\]\[18\] _1719_ _1722_ VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5952_ _2503_ _2693_ _2694_ VGND VGND VPWR VPWR _2695_ sky130_fd_sc_hd__or3_1
X_8740_ clknet_leaf_89_CLK _0924_ VGND VGND VPWR VPWR RF.registers\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4903_ _1655_ _1658_ net5 VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_36_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5883_ _2427_ _2591_ _2628_ _2504_ VGND VGND VPWR VPWR _2629_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8671_ clknet_leaf_64_CLK _0855_ VGND VGND VPWR VPWR RF.registers\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7622_ _3767_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4834_ RF.registers\[16\]\[17\] RF.registers\[17\]\[17\] RF.registers\[18\]\[17\]
+ RF.registers\[19\]\[17\] _1291_ _1194_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__mux4_1
X_7553_ _3081_ RF.registers\[27\]\[28\] _3722_ VGND VGND VPWR VPWR _3731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4765_ _1107_ _1520_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_134_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6504_ RF.registers\[0\]\[0\] _3089_ _3157_ VGND VGND VPWR VPWR _3158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7484_ _3694_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9223_ clknet_leaf_59_CLK _0383_ VGND VGND VPWR VPWR RF.registers\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_4696_ RF.registers\[28\]\[12\] RF.registers\[29\]\[12\] RF.registers\[30\]\[12\]
+ RF.registers\[31\]\[12\] _1219_ _1221_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__mux4_1
X_6435_ RF.registers\[17\]\[9\] _3111_ _3093_ VGND VGND VPWR VPWR _3112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6366_ net26 VGND VGND VPWR VPWR _3064_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_58_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9154_ clknet_leaf_91_CLK _0314_ VGND VGND VPWR VPWR RF.registers\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8105_ _4023_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__clkbuf_1
X_9085_ clknet_leaf_19_CLK _0245_ VGND VGND VPWR VPWR RF.registers\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5317_ _1684_ _2072_ VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__and2_1
X_6297_ _3016_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__clkbuf_1
X_8036_ _3986_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__clkbuf_1
X_5248_ RF.registers\[24\]\[25\] RF.registers\[25\]\[25\] RF.registers\[26\]\[25\]
+ RF.registers\[27\]\[25\] _1822_ _1823_ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5179_ _1889_ _1934_ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8938_ clknet_leaf_82_CLK _0098_ VGND VGND VPWR VPWR RF.registers\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_119_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8869_ clknet_leaf_81_CLK _0029_ VGND VGND VPWR VPWR RF.registers\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_128_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_137_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4550_ _1302_ _1305_ _1187_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4481_ _1171_ _1228_ _1236_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a21oi_2
X_6220_ _1060_ _2678_ _2737_ _2947_ VGND VGND VPWR VPWR _2948_ sky130_fd_sc_hd__o22a_1
X_6151_ _2812_ _2878_ _2882_ VGND VGND VPWR VPWR _2883_ sky130_fd_sc_hd__o21a_1
X_5102_ _1672_ _1849_ _1853_ _1857_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_57_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _2812_ _2817_ VGND VGND VPWR VPWR _2818_ sky130_fd_sc_hd__nand2_1
X_5033_ _1785_ _1788_ _1699_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__mux2_1
X_6984_ RF.registers\[3\]\[0\] _3089_ _3413_ VGND VGND VPWR VPWR _3414_ sky130_fd_sc_hd__mux2_1
X_8723_ clknet_leaf_36_CLK _0907_ VGND VGND VPWR VPWR RF.registers\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5935_ _1666_ _2039_ _2251_ VGND VGND VPWR VPWR _2679_ sky130_fd_sc_hd__or3b_1
X_8654_ clknet_leaf_40_CLK _0838_ VGND VGND VPWR VPWR RF.registers\[0\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5866_ _2340_ _2487_ _2612_ _2530_ VGND VGND VPWR VPWR _2613_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7605_ _3064_ RF.registers\[28\]\[20\] _3758_ VGND VGND VPWR VPWR _3759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4817_ _1528_ _1542_ _1558_ _1572_ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__and4b_1
XFILLER_0_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5797_ _1669_ _2272_ _2325_ VGND VGND VPWR VPWR _2547_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8585_ clknet_leaf_1_CLK _0769_ VGND VGND VPWR VPWR RF.registers\[22\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_7536_ _3699_ VGND VGND VPWR VPWR _3722_ sky130_fd_sc_hd__clkbuf_8
X_4748_ RF.registers\[12\]\[15\] RF.registers\[13\]\[15\] RF.registers\[14\]\[15\]
+ RF.registers\[15\]\[15\] _1201_ _1203_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4679_ RF.registers\[24\]\[22\] RF.registers\[25\]\[22\] RF.registers\[26\]\[22\]
+ RF.registers\[27\]\[22\] _1182_ _1184_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__mux4_1
X_7467_ _3685_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9206_ clknet_leaf_32_CLK _0366_ VGND VGND VPWR VPWR RF.registers\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6418_ _3100_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__clkbuf_1
X_7398_ _3062_ RF.registers\[26\]\[19\] _3639_ VGND VGND VPWR VPWR _3649_ sky130_fd_sc_hd__mux2_1
X_9137_ clknet_leaf_6_CLK _0297_ VGND VGND VPWR VPWR RF.registers\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xoutput59 net59 VGND VGND VPWR VPWR ALU_result[19] sky130_fd_sc_hd__buf_1
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6349_ _3052_ RF.registers\[22\]\[14\] _3044_ VGND VGND VPWR VPWR _3053_ sky130_fd_sc_hd__mux2_1
X_9068_ clknet_leaf_3_CLK _0228_ VGND VGND VPWR VPWR RF.registers\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8019_ _3141_ RF.registers\[21\]\[23\] _3974_ VGND VGND VPWR VPWR _3978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5720_ _2381_ VGND VGND VPWR VPWR _2473_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5651_ _2390_ _2405_ _2104_ VGND VGND VPWR VPWR _2406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4602_ _1356_ _1357_ _1199_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__mux2_1
X_8370_ RF.registers\[16\]\[28\] _3446_ _4155_ VGND VGND VPWR VPWR _4164_ sky130_fd_sc_hd__mux2_1
X_5582_ _2336_ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__buf_2
X_4533_ _1287_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__and2_1
X_7321_ _3054_ RF.registers\[31\]\[15\] _3602_ VGND VGND VPWR VPWR _3608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7252_ _3571_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6203_ _1237_ _2930_ VGND VGND VPWR VPWR _2931_ sky130_fd_sc_hd__xnor2_1
X_4464_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7183_ RF.registers\[7\]\[15\] _3487_ _3528_ VGND VGND VPWR VPWR _3534_ sky130_fd_sc_hd__mux2_1
X_4395_ RF.registers\[16\]\[0\] RF.registers\[17\]\[0\] RF.registers\[18\]\[0\] RF.registers\[19\]\[0\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_129_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6134_ _1669_ _1732_ _2035_ VGND VGND VPWR VPWR _2866_ sky130_fd_sc_hd__a21oi_1
X_6065_ _2777_ _2800_ _1147_ VGND VGND VPWR VPWR _2801_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _1766_ _1771_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6967_ RF.registers\[4\]\[25\] _3145_ _3398_ VGND VGND VPWR VPWR _3404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5918_ _2175_ _2659_ _2660_ VGND VGND VPWR VPWR _2662_ sky130_fd_sc_hd__nand3_1
X_8706_ clknet_leaf_90_CLK _0890_ VGND VGND VPWR VPWR RF.registers\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6898_ _3367_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_66_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8637_ clknet_leaf_18_CLK _0821_ VGND VGND VPWR VPWR RF.registers\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5849_ _1528_ _2596_ VGND VGND VPWR VPWR _2597_ sky130_fd_sc_hd__xor2_2
XFILLER_0_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8568_ clknet_leaf_14_CLK _0752_ VGND VGND VPWR VPWR RF.registers\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7519_ _3713_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
X_8499_ _4232_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7870_ _3128_ RF.registers\[23\]\[17\] _3891_ VGND VGND VPWR VPWR _3899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6821_ RF.registers\[6\]\[20\] _3134_ _3326_ VGND VGND VPWR VPWR _3327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9540_ clknet_leaf_88_CLK _0700_ VGND VGND VPWR VPWR RF.registers\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6752_ _3064_ RF.registers\[14\]\[20\] _3289_ VGND VGND VPWR VPWR _3290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6683_ _3230_ VGND VGND VPWR VPWR _3253_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5703_ _2368_ _2367_ VGND VGND VPWR VPWR _2456_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9471_ clknet_leaf_64_CLK _0631_ VGND VGND VPWR VPWR RF.registers\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8422_ RF.registers\[12\]\[20\] _3497_ _4191_ VGND VGND VPWR VPWR _4192_ sky130_fd_sc_hd__mux2_1
X_5634_ _2388_ VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8353_ _4132_ VGND VGND VPWR VPWR _4155_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5565_ _2319_ _2320_ _2044_ VGND VGND VPWR VPWR _2321_ sky130_fd_sc_hd__mux2_1
X_7304_ _3037_ RF.registers\[31\]\[7\] _3591_ VGND VGND VPWR VPWR _3599_ sky130_fd_sc_hd__mux2_1
X_4516_ _1214_ _1271_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__nand2_1
X_5496_ _2251_ VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__clkbuf_4
X_8284_ _4118_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4447_ _1202_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__clkbuf_8
X_7235_ _3562_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7166_ RF.registers\[7\]\[7\] _3470_ _3517_ VGND VGND VPWR VPWR _3525_ sky130_fd_sc_hd__mux2_1
X_6117_ _2549_ _2823_ _2731_ _2705_ _2850_ VGND VGND VPWR VPWR _2851_ sky130_fd_sc_hd__a221o_1
X_4378_ _1132_ _1133_ _1035_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__mux2_1
X_7097_ _3482_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
X_6048_ _1820_ _2768_ VGND VGND VPWR VPWR _2785_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7999_ _3967_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5350_ RF.registers\[20\]\[15\] RF.registers\[21\]\[15\] RF.registers\[22\]\[15\]
+ RF.registers\[23\]\[15\] _1734_ _1680_ VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5281_ _1999_ _2036_ _1877_ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__mux2_1
X_4301_ net8 VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__buf_4
X_7020_ _3432_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8971_ clknet_leaf_0_CLK _0131_ VGND VGND VPWR VPWR RF.registers\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7922_ _3926_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__clkbuf_1
X_7853_ _3111_ RF.registers\[23\]\[9\] _3880_ VGND VGND VPWR VPWR _3890_ sky130_fd_sc_hd__mux2_1
X_4996_ _1750_ _1751_ _1739_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__mux2_1
X_7784_ _3853_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__clkbuf_1
X_6804_ RF.registers\[6\]\[12\] _3118_ _3315_ VGND VGND VPWR VPWR _3318_ sky130_fd_sc_hd__mux2_1
X_9523_ clknet_leaf_30_CLK _0683_ VGND VGND VPWR VPWR RF.registers\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6735_ _3048_ RF.registers\[14\]\[12\] _3278_ VGND VGND VPWR VPWR _3281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9454_ clknet_leaf_14_CLK _0614_ VGND VGND VPWR VPWR RF.registers\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6666_ _3244_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5617_ _1060_ _2101_ VGND VGND VPWR VPWR _2372_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9385_ clknet_leaf_9_CLK _0545_ VGND VGND VPWR VPWR RF.registers\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6597_ _3046_ RF.registers\[15\]\[11\] _3206_ VGND VGND VPWR VPWR _3208_ sky130_fd_sc_hd__mux2_1
X_8405_ RF.registers\[12\]\[12\] _3481_ _4180_ VGND VGND VPWR VPWR _4183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5548_ _1696_ _2303_ _1670_ VGND VGND VPWR VPWR _2304_ sky130_fd_sc_hd__o21ai_1
X_8336_ _4146_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__clkbuf_1
X_8267_ _3116_ RF.registers\[13\]\[11\] _4108_ VGND VGND VPWR VPWR _4110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7218_ net10 net9 net46 VGND VGND VPWR VPWR _3552_ sky130_fd_sc_hd__and3b_4
X_5479_ RF.registers\[16\]\[9\] RF.registers\[17\]\[9\] RF.registers\[18\]\[9\] RF.registers\[19\]\[9\]
+ _1675_ _1692_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8198_ _4073_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__clkbuf_1
X_7149_ _3515_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_100_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4850_ RF.registers\[28\]\[19\] RF.registers\[29\]\[19\] RF.registers\[30\]\[19\]
+ RF.registers\[31\]\[19\] _1220_ _1222_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4781_ _1040_ _1536_ _1037_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__o21a_1
X_6520_ RF.registers\[0\]\[8\] _3109_ _3157_ VGND VGND VPWR VPWR _3166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload20 clknet_leaf_9_CLK VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__clkinvlp_4
X_6451_ RF.registers\[17\]\[14\] _3122_ _3114_ VGND VGND VPWR VPWR _3123_ sky130_fd_sc_hd__mux2_1
X_6382_ net31 VGND VGND VPWR VPWR _3075_ sky130_fd_sc_hd__buf_2
X_9170_ clknet_leaf_54_CLK _0330_ VGND VGND VPWR VPWR RF.registers\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xclkload42 clknet_leaf_57_CLK VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__inv_6
Xclkload53 clknet_leaf_6_CLK VGND VGND VPWR VPWR clkload53/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload31 clknet_leaf_68_CLK VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5402_ _2156_ _2157_ net3 VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__mux2_1
Xclkload86 clknet_leaf_31_CLK VGND VGND VPWR VPWR clkload86/Y sky130_fd_sc_hd__clkinv_1
Xclkload75 clknet_leaf_42_CLK VGND VGND VPWR VPWR clkload75/Y sky130_fd_sc_hd__clkinvlp_2
Xclkload64 clknet_leaf_39_CLK VGND VGND VPWR VPWR clkload64/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8121_ _4032_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5333_ RF.registers\[4\]\[1\] RF.registers\[5\]\[1\] RF.registers\[6\]\[1\] RF.registers\[7\]\[1\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__mux4_1
X_5264_ _2018_ _2019_ _1901_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8052_ RF.registers\[20\]\[6\] _3468_ _3989_ VGND VGND VPWR VPWR _3996_ sky130_fd_sc_hd__mux2_1
X_5195_ _1889_ _1950_ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7003_ _3423_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
X_8954_ clknet_leaf_35_CLK _0114_ VGND VGND VPWR VPWR RF.registers\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8885_ clknet_leaf_51_CLK _0045_ VGND VGND VPWR VPWR RF.registers\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7905_ RF.registers\[18\]\[1\] _3458_ _3916_ VGND VGND VPWR VPWR _3918_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7836_ _3881_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7767_ RF.registers\[9\]\[0\] _3454_ _3844_ VGND VGND VPWR VPWR _3845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4979_ _1721_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload3 clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinvlp_4
X_7698_ _3807_ VGND VGND VPWR VPWR _3808_ sky130_fd_sc_hd__buf_6
X_9506_ clknet_leaf_91_CLK _0666_ VGND VGND VPWR VPWR RF.registers\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6718_ _3031_ RF.registers\[14\]\[4\] _3267_ VGND VGND VPWR VPWR _3272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9437_ clknet_leaf_16_CLK _0597_ VGND VGND VPWR VPWR RF.registers\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6649_ _3235_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9368_ clknet_leaf_39_CLK _0528_ VGND VGND VPWR VPWR RF.registers\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_76_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9299_ clknet_leaf_28_CLK _0459_ VGND VGND VPWR VPWR RF.registers\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_8319_ _4137_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5951_ _2522_ _2605_ _2591_ _2531_ VGND VGND VPWR VPWR _2694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8670_ clknet_leaf_69_CLK _0854_ VGND VGND VPWR VPWR RF.registers\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_4902_ _1656_ _1657_ _1645_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5882_ _2441_ _2588_ _2590_ _2444_ VGND VGND VPWR VPWR _2628_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7621_ _3081_ RF.registers\[28\]\[28\] _3758_ VGND VGND VPWR VPWR _3767_ sky130_fd_sc_hd__mux2_1
X_4833_ RF.registers\[28\]\[17\] RF.registers\[29\]\[17\] RF.registers\[30\]\[17\]
+ RF.registers\[31\]\[17\] _1191_ _1174_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7552_ _3730_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4764_ RF.registers\[12\]\[8\] RF.registers\[13\]\[8\] RF.registers\[14\]\[8\] RF.registers\[15\]\[8\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_134_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7483_ _3079_ RF.registers\[25\]\[27\] _3686_ VGND VGND VPWR VPWR _3694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6503_ _3156_ VGND VGND VPWR VPWR _3157_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9222_ clknet_leaf_61_CLK _0382_ VGND VGND VPWR VPWR RF.registers\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_4695_ _1449_ _1450_ _1036_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6434_ net45 VGND VGND VPWR VPWR _3111_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6365_ _3063_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9153_ clknet_leaf_73_CLK _0313_ VGND VGND VPWR VPWR RF.registers\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6296_ RF.registers\[10\]\[30\] _3015_ _3007_ VGND VGND VPWR VPWR _3016_ sky130_fd_sc_hd__mux2_1
X_9084_ clknet_leaf_23_CLK _0244_ VGND VGND VPWR VPWR RF.registers\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_8104_ RF.registers\[20\]\[31\] _3452_ _3988_ VGND VGND VPWR VPWR _4023_ sky130_fd_sc_hd__mux2_1
X_5316_ RF.registers\[8\]\[2\] RF.registers\[9\]\[2\] RF.registers\[10\]\[2\] RF.registers\[11\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__mux4_1
X_5247_ RF.registers\[28\]\[25\] RF.registers\[29\]\[25\] RF.registers\[30\]\[25\]
+ RF.registers\[31\]\[25\] _1822_ _1823_ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__mux4_1
X_8035_ _3017_ RF.registers\[21\]\[31\] _3951_ VGND VGND VPWR VPWR _3986_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5178_ RF.registers\[4\]\[29\] RF.registers\[5\]\[29\] RF.registers\[6\]\[29\] RF.registers\[7\]\[29\]
+ _1767_ _1768_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8937_ clknet_leaf_85_CLK _0097_ VGND VGND VPWR VPWR RF.registers\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8868_ clknet_leaf_90_CLK _0028_ VGND VGND VPWR VPWR RF.registers\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_7819_ RF.registers\[9\]\[25\] _3508_ _3866_ VGND VGND VPWR VPWR _3872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8799_ clknet_leaf_66_CLK _0983_ VGND VGND VPWR VPWR RF.registers\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4480_ _1230_ _1232_ _1235_ _1205_ _1215_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6150_ _2840_ _2843_ _2854_ _2880_ _2881_ VGND VGND VPWR VPWR _2882_ sky130_fd_sc_hd__o311a_1
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5101_ _1717_ _1856_ _1729_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _2814_ _2815_ _2748_ _2816_ VGND VGND VPWR VPWR _2817_ sky130_fd_sc_hd__a31o_1
X_5032_ _1786_ _1787_ _1739_ VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6983_ _3412_ VGND VGND VPWR VPWR _3413_ sky130_fd_sc_hd__clkbuf_8
X_8722_ clknet_leaf_54_CLK _0906_ VGND VGND VPWR VPWR RF.registers\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5934_ _2502_ _2677_ _2104_ VGND VGND VPWR VPWR _2678_ sky130_fd_sc_hd__mux2_1
X_5865_ _2426_ _2608_ _2611_ VGND VGND VPWR VPWR _2612_ sky130_fd_sc_hd__o21ai_1
X_8653_ clknet_leaf_57_CLK _0837_ VGND VGND VPWR VPWR RF.registers\[0\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_7604_ _3735_ VGND VGND VPWR VPWR _3758_ sky130_fd_sc_hd__buf_4
XFILLER_0_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4816_ _1025_ _1563_ _1567_ _1571_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5796_ _2363_ _1758_ _2331_ _2419_ VGND VGND VPWR VPWR _2546_ sky130_fd_sc_hd__o31ai_1
X_8584_ clknet_leaf_96_CLK _0768_ VGND VGND VPWR VPWR RF.registers\[22\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7535_ _3721_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
X_4747_ RF.registers\[8\]\[15\] RF.registers\[9\]\[15\] RF.registers\[10\]\[15\] RF.registers\[11\]\[15\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__mux4_1
X_4678_ RF.registers\[28\]\[22\] RF.registers\[29\]\[22\] RF.registers\[30\]\[22\]
+ RF.registers\[31\]\[22\] _1182_ _1184_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__mux4_1
X_7466_ _3062_ RF.registers\[25\]\[19\] _3675_ VGND VGND VPWR VPWR _3685_ sky130_fd_sc_hd__mux2_1
X_9205_ clknet_leaf_25_CLK _0365_ VGND VGND VPWR VPWR RF.registers\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7397_ _3648_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
X_6417_ RF.registers\[17\]\[3\] _3099_ _3093_ VGND VGND VPWR VPWR _3100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9136_ clknet_leaf_6_CLK _0296_ VGND VGND VPWR VPWR RF.registers\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
Xoutput49 net49 VGND VGND VPWR VPWR ALU_result[0] sky130_fd_sc_hd__buf_1
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6348_ net19 VGND VGND VPWR VPWR _3052_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6279_ net13 net11 net12 VGND VGND VPWR VPWR _3003_ sky130_fd_sc_hd__or3b_4
X_9067_ clknet_leaf_98_CLK _0227_ VGND VGND VPWR VPWR RF.registers\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_8018_ _3977_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_40_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5650_ _2404_ VGND VGND VPWR VPWR _2405_ sky130_fd_sc_hd__inv_2
X_4601_ RF.registers\[24\]\[25\] RF.registers\[25\]\[25\] RF.registers\[26\]\[25\]
+ RF.registers\[27\]\[25\] _1351_ _1352_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5581_ _1111_ _1126_ VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__nand2_2
XFILLER_0_53_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4532_ RF.registers\[4\]\[26\] RF.registers\[5\]\[26\] RF.registers\[6\]\[26\] RF.registers\[7\]\[26\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7320_ _3607_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4463_ _1089_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__buf_4
X_7251_ _3052_ RF.registers\[29\]\[14\] _3566_ VGND VGND VPWR VPWR _3571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6202_ _2595_ _2929_ VGND VGND VPWR VPWR _2930_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_31_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_55_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7182_ _3533_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_4394_ RF.registers\[20\]\[0\] RF.registers\[21\]\[0\] RF.registers\[22\]\[0\] RF.registers\[23\]\[0\]
+ _1149_ _1061_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6133_ _2038_ _2864_ VGND VGND VPWR VPWR _2865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6064_ _1840_ _1801_ VGND VGND VPWR VPWR _2800_ sky130_fd_sc_hd__and2b_1
X_5015_ _1769_ _1770_ _1713_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6966_ _3403_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_98_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_98_CLK sky130_fd_sc_hd__clkbuf_8
X_5917_ _2659_ _2660_ _2175_ VGND VGND VPWR VPWR _2661_ sky130_fd_sc_hd__a21o_1
X_8705_ clknet_leaf_91_CLK _0889_ VGND VGND VPWR VPWR RF.registers\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6897_ RF.registers\[5\]\[24\] _3143_ _3362_ VGND VGND VPWR VPWR _3367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8636_ clknet_leaf_23_CLK _0820_ VGND VGND VPWR VPWR RF.registers\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_5848_ _1416_ _2593_ _2594_ _2595_ VGND VGND VPWR VPWR _2596_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8567_ _4267_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5779_ _1111_ VGND VGND VPWR VPWR _2530_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7518_ _3046_ RF.registers\[27\]\[11\] _3711_ VGND VGND VPWR VPWR _3713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8498_ RF.registers\[11\]\[24\] net30 _4227_ VGND VGND VPWR VPWR _4232_ sky130_fd_sc_hd__mux2_1
X_7449_ _3676_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_22_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9119_ clknet_leaf_71_CLK _0279_ VGND VGND VPWR VPWR RF.registers\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_89_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_89_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_13_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6820_ _3303_ VGND VGND VPWR VPWR _3326_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6751_ _3266_ VGND VGND VPWR VPWR _3289_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6682_ _3252_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5702_ _2339_ VGND VGND VPWR VPWR _2455_ sky130_fd_sc_hd__inv_2
X_9470_ clknet_leaf_68_CLK _0630_ VGND VGND VPWR VPWR RF.registers\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8421_ _4168_ VGND VGND VPWR VPWR _4191_ sky130_fd_sc_hd__buf_4
X_5633_ _2385_ _2387_ _1145_ VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8352_ _4154_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__clkbuf_1
X_5564_ RF.registers\[0\]\[5\] RF.registers\[1\]\[5\] RF.registers\[2\]\[5\] RF.registers\[3\]\[5\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2320_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4515_ _1269_ _1270_ _1190_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7303_ _3598_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8283_ _3132_ RF.registers\[13\]\[19\] _4108_ VGND VGND VPWR VPWR _4118_ sky130_fd_sc_hd__mux2_1
X_5495_ _1125_ VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__clkbuf_4
X_4446_ _1029_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__clkbuf_4
X_7234_ _3035_ RF.registers\[29\]\[6\] _3555_ VGND VGND VPWR VPWR _3562_ sky130_fd_sc_hd__mux2_1
X_7165_ _3524_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_4377_ RF.registers\[24\]\[1\] RF.registers\[25\]\[1\] RF.registers\[26\]\[1\] RF.registers\[27\]\[1\]
+ _1041_ _1043_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6116_ _2495_ _2849_ _2503_ VGND VGND VPWR VPWR _2850_ sky130_fd_sc_hd__a21o_1
X_7096_ RF.registers\[19\]\[12\] _3481_ _3477_ VGND VGND VPWR VPWR _3482_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_13_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6047_ _1838_ _2783_ VGND VGND VPWR VPWR _2784_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_68_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ _3120_ RF.registers\[21\]\[13\] _3963_ VGND VGND VPWR VPWR _3967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6949_ _3394_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8619_ clknet_leaf_98_CLK _0803_ VGND VGND VPWR VPWR RF.registers\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_2_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5280_ _2017_ _2035_ VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__or2_1
X_4300_ _1054_ _1055_ _1047_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8970_ clknet_leaf_8_CLK _0130_ VGND VGND VPWR VPWR RF.registers\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7921_ RF.registers\[18\]\[9\] _3474_ _3916_ VGND VGND VPWR VPWR _3926_ sky130_fd_sc_hd__mux2_1
X_7852_ _3889_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__clkbuf_1
X_4995_ RF.registers\[0\]\[22\] RF.registers\[1\]\[22\] RF.registers\[2\]\[22\] RF.registers\[3\]\[22\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6803_ _3317_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__clkbuf_1
X_7783_ RF.registers\[9\]\[8\] _3472_ _3844_ VGND VGND VPWR VPWR _3853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9522_ clknet_leaf_43_CLK _0682_ VGND VGND VPWR VPWR RF.registers\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6734_ _3280_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9453_ clknet_leaf_10_CLK _0613_ VGND VGND VPWR VPWR RF.registers\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6665_ RF.registers\[8\]\[11\] _3116_ _3242_ VGND VGND VPWR VPWR _3244_ sky130_fd_sc_hd__mux2_1
X_8404_ _4182_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5616_ _2366_ _2367_ _2370_ _2336_ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__a211o_1
X_9384_ clknet_leaf_1_CLK _0544_ VGND VGND VPWR VPWR RF.registers\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6596_ _3207_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__clkbuf_1
X_5547_ _2301_ _2302_ _1738_ VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__mux2_1
X_8335_ RF.registers\[16\]\[11\] _3479_ _4144_ VGND VGND VPWR VPWR _4146_ sky130_fd_sc_hd__mux2_1
X_5478_ RF.registers\[20\]\[9\] RF.registers\[21\]\[9\] RF.registers\[22\]\[9\] RF.registers\[23\]\[9\]
+ _1675_ _1692_ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8266_ _4109_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4429_ RF.registers\[24\]\[29\] RF.registers\[25\]\[29\] RF.registers\[26\]\[29\]
+ RF.registers\[27\]\[29\] _1182_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__mux4_1
X_7217_ _3551_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8197_ RF.registers\[1\]\[10\] _3476_ _4072_ VGND VGND VPWR VPWR _4073_ sky130_fd_sc_hd__mux2_1
X_7148_ RF.registers\[19\]\[31\] _3452_ _3455_ VGND VGND VPWR VPWR _3515_ sky130_fd_sc_hd__mux2_1
X_7079_ net43 VGND VGND VPWR VPWR _3470_ sky130_fd_sc_hd__buf_2
XFILLER_0_138_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4780_ RF.registers\[12\]\[9\] RF.registers\[13\]\[9\] RF.registers\[14\]\[9\] RF.registers\[15\]\[9\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload10 clknet_leaf_92_CLK VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6450_ net19 VGND VGND VPWR VPWR _3122_ sky130_fd_sc_hd__buf_2
X_6381_ _3074_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__clkbuf_1
Xclkload43 clknet_leaf_58_CLK VGND VGND VPWR VPWR clkload43/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload21 clknet_leaf_10_CLK VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_11_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload32 clknet_leaf_69_CLK VGND VGND VPWR VPWR clkload32/X sky130_fd_sc_hd__clkbuf_4
X_5401_ RF.registers\[12\]\[13\] RF.registers\[13\]\[13\] RF.registers\[14\]\[13\]
+ RF.registers\[15\]\[13\] _1702_ _1678_ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__mux4_1
Xclkload87 clknet_leaf_32_CLK VGND VGND VPWR VPWR clkload87/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload65 clknet_leaf_17_CLK VGND VGND VPWR VPWR clkload65/Y sky130_fd_sc_hd__inv_8
Xclkload76 clknet_leaf_43_CLK VGND VGND VPWR VPWR clkload76/Y sky130_fd_sc_hd__clkinv_4
Xclkload54 clknet_leaf_7_CLK VGND VGND VPWR VPWR clkload54/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8120_ RF.registers\[24\]\[6\] _3468_ _4025_ VGND VGND VPWR VPWR _4032_ sky130_fd_sc_hd__mux2_1
X_5332_ _2084_ _2085_ _2086_ _2087_ net3 _1655_ VGND VGND VPWR VPWR _2088_ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5263_ RF.registers\[16\]\[24\] RF.registers\[17\]\[24\] RF.registers\[18\]\[24\]
+ RF.registers\[19\]\[24\] _1918_ _1919_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__mux4_1
X_8051_ _3995_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__clkbuf_1
X_5194_ RF.registers\[4\]\[28\] RF.registers\[5\]\[28\] RF.registers\[6\]\[28\] RF.registers\[7\]\[28\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7002_ RF.registers\[3\]\[9\] _3111_ _3413_ VGND VGND VPWR VPWR _3423_ sky130_fd_sc_hd__mux2_1
X_8953_ clknet_leaf_50_CLK _0113_ VGND VGND VPWR VPWR RF.registers\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8884_ clknet_leaf_53_CLK _0044_ VGND VGND VPWR VPWR RF.registers\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7904_ _3917_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7835_ _3089_ RF.registers\[23\]\[0\] _3880_ VGND VGND VPWR VPWR _3881_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7766_ _3843_ VGND VGND VPWR VPWR _3844_ sky130_fd_sc_hd__clkbuf_8
X_9505_ clknet_leaf_92_CLK _0665_ VGND VGND VPWR VPWR RF.registers\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4978_ _1733_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload4 clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_12
X_7697_ _3020_ _3553_ VGND VGND VPWR VPWR _3807_ sky130_fd_sc_hd__nand2_4
X_6717_ _3271_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9436_ clknet_leaf_37_CLK _0596_ VGND VGND VPWR VPWR RF.registers\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6648_ RF.registers\[8\]\[3\] _3099_ _3231_ VGND VGND VPWR VPWR _3235_ sky130_fd_sc_hd__mux2_1
X_9367_ clknet_leaf_32_CLK _0527_ VGND VGND VPWR VPWR RF.registers\[20\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8318_ RF.registers\[16\]\[3\] _3462_ _4133_ VGND VGND VPWR VPWR _4137_ sky130_fd_sc_hd__mux2_1
X_6579_ _3198_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9298_ clknet_leaf_42_CLK _0458_ VGND VGND VPWR VPWR RF.registers\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8249_ _4100_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5950_ _2692_ _2679_ VGND VGND VPWR VPWR _2693_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4901_ RF.registers\[0\]\[0\] RF.registers\[1\]\[0\] RF.registers\[2\]\[0\] RF.registers\[3\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_36_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7620_ _3766_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5881_ _2335_ _2626_ VGND VGND VPWR VPWR _2627_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4832_ RF.registers\[24\]\[17\] RF.registers\[25\]\[17\] RF.registers\[26\]\[17\]
+ RF.registers\[27\]\[17\] _1291_ _1194_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7551_ _3079_ RF.registers\[27\]\[27\] _3722_ VGND VGND VPWR VPWR _3730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4763_ _1515_ _1518_ _1037_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7482_ _3693_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__clkbuf_1
X_6502_ _3153_ _3155_ VGND VGND VPWR VPWR _3156_ sky130_fd_sc_hd__nor2_4
XFILLER_0_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4694_ RF.registers\[16\]\[12\] RF.registers\[17\]\[12\] RF.registers\[18\]\[12\]
+ RF.registers\[19\]\[12\] _1219_ _1221_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9221_ clknet_leaf_59_CLK _0381_ VGND VGND VPWR VPWR RF.registers\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6433_ _3110_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6364_ _3062_ RF.registers\[22\]\[19\] _3044_ VGND VGND VPWR VPWR _3063_ sky130_fd_sc_hd__mux2_1
X_9152_ clknet_leaf_70_CLK _0312_ VGND VGND VPWR VPWR RF.registers\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9083_ clknet_leaf_46_CLK _0243_ VGND VGND VPWR VPWR RF.registers\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_8103_ _4022_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__clkbuf_1
X_6295_ net37 VGND VGND VPWR VPWR _3015_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5315_ _2067_ _2070_ net4 VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__mux2_1
X_5246_ _2000_ _2001_ _1726_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__mux2_1
X_8034_ _3985_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5177_ _1929_ _1932_ _1700_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8936_ clknet_leaf_78_CLK _0096_ VGND VGND VPWR VPWR RF.registers\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8867_ clknet_leaf_75_CLK _0027_ VGND VGND VPWR VPWR RF.registers\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_7818_ _3871_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8798_ clknet_leaf_67_CLK _0982_ VGND VGND VPWR VPWR RF.registers\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7749_ _3073_ RF.registers\[30\]\[24\] _3830_ VGND VGND VPWR VPWR _3835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9419_ clknet_leaf_78_CLK _0579_ VGND VGND VPWR VPWR RF.registers\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6080_ _2770_ _2809_ VGND VGND VPWR VPWR _2816_ sky130_fd_sc_hd__or2_1
X_5100_ _1854_ _1855_ _1726_ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ RF.registers\[24\]\[20\] RF.registers\[25\]\[20\] RF.registers\[26\]\[20\]
+ RF.registers\[27\]\[20\] _1782_ _1680_ VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8721_ clknet_leaf_39_CLK _0905_ VGND VGND VPWR VPWR RF.registers\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6982_ _3153_ _3411_ VGND VGND VPWR VPWR _3412_ sky130_fd_sc_hd__nor2_4
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5933_ _2673_ _2676_ _2501_ VGND VGND VPWR VPWR _2677_ sky130_fd_sc_hd__mux2_1
X_5864_ _2252_ _2610_ VGND VGND VPWR VPWR _2611_ sky130_fd_sc_hd__nand2_1
X_8652_ clknet_leaf_83_CLK _0836_ VGND VGND VPWR VPWR RF.registers\[0\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_7603_ _3757_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
X_8583_ clknet_leaf_58_CLK _0767_ VGND VGND VPWR VPWR RF.registers\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4815_ _1088_ _1570_ net8 VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__a21oi_1
X_7534_ _3062_ RF.registers\[27\]\[19\] _3711_ VGND VGND VPWR VPWR _3721_ sky130_fd_sc_hd__mux2_1
X_5795_ _2539_ _2540_ _2543_ VGND VGND VPWR VPWR _2545_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4746_ _1498_ _1501_ _1187_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4677_ _1431_ _1432_ _1178_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__mux2_1
X_7465_ _3684_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9204_ clknet_leaf_23_CLK _0364_ VGND VGND VPWR VPWR RF.registers\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_7396_ _3060_ RF.registers\[26\]\[18\] _3639_ VGND VGND VPWR VPWR _3648_ sky130_fd_sc_hd__mux2_1
X_6416_ net39 VGND VGND VPWR VPWR _3099_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_73_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9135_ clknet_leaf_6_CLK _0295_ VGND VGND VPWR VPWR RF.registers\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6347_ _3051_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6278_ net32 VGND VGND VPWR VPWR _3002_ sky130_fd_sc_hd__buf_2
X_9066_ clknet_leaf_8_CLK _0226_ VGND VGND VPWR VPWR RF.registers\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8017_ _3139_ RF.registers\[21\]\[22\] _3974_ VGND VGND VPWR VPWR _3977_ sky130_fd_sc_hd__mux2_1
X_5229_ RF.registers\[24\]\[26\] RF.registers\[25\]\[26\] RF.registers\[26\]\[26\]
+ RF.registers\[27\]\[26\] _1881_ _1883_ VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__mux4_1
X_8919_ clknet_leaf_32_CLK _0079_ VGND VGND VPWR VPWR RF.registers\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4600_ RF.registers\[28\]\[25\] RF.registers\[29\]\[25\] RF.registers\[30\]\[25\]
+ RF.registers\[31\]\[25\] _1351_ _1352_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5580_ _1060_ _1085_ VGND VGND VPWR VPWR _2335_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_68_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4531_ _1048_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__buf_4
X_4462_ RF.registers\[20\]\[28\] RF.registers\[21\]\[28\] RF.registers\[22\]\[28\]
+ RF.registers\[23\]\[28\] _1182_ _1184_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__mux4_1
XFILLER_0_80_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7250_ _3570_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6201_ _1316_ _1385_ _2872_ VGND VGND VPWR VPWR _2929_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7181_ RF.registers\[7\]\[14\] _3485_ _3528_ VGND VGND VPWR VPWR _3533_ sky130_fd_sc_hd__mux2_1
X_4393_ A2[0] VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__buf_4
X_6132_ _2104_ _2373_ VGND VGND VPWR VPWR _2864_ sky130_fd_sc_hd__nand2_1
X_6063_ _2583_ _2733_ _2426_ VGND VGND VPWR VPWR _2799_ sky130_fd_sc_hd__mux2_1
X_5014_ RF.registers\[12\]\[21\] RF.registers\[13\]\[21\] RF.registers\[14\]\[21\]
+ RF.registers\[15\]\[21\] _1767_ _1768_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6965_ RF.registers\[4\]\[24\] _3143_ _3398_ VGND VGND VPWR VPWR _3403_ sky130_fd_sc_hd__mux2_1
X_5916_ _2536_ _2658_ _1464_ VGND VGND VPWR VPWR _2660_ sky130_fd_sc_hd__o21ai_1
X_8704_ clknet_leaf_71_CLK _0888_ VGND VGND VPWR VPWR RF.registers\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8635_ clknet_leaf_46_CLK _0819_ VGND VGND VPWR VPWR RF.registers\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6896_ _3366_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5847_ net47 _2503_ VGND VGND VPWR VPWR _2595_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8566_ RF.registers\[10\]\[25\] net31 _3006_ VGND VGND VPWR VPWR _4267_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_86_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5778_ _1666_ _2523_ _2528_ _2495_ VGND VGND VPWR VPWR _2529_ sky130_fd_sc_hd__a2bb2o_1
X_8497_ _4231_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7517_ _3712_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__clkbuf_1
X_4729_ _1481_ _1482_ _1483_ _1484_ _1189_ _1078_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__mux4_2
X_7448_ _3043_ RF.registers\[25\]\[10\] _3675_ VGND VGND VPWR VPWR _3676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7379_ _3627_ VGND VGND VPWR VPWR _3639_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9118_ clknet_leaf_68_CLK _0278_ VGND VGND VPWR VPWR RF.registers\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_9049_ clknet_leaf_26_CLK _0209_ VGND VGND VPWR VPWR RF.registers\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_95_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6750_ _3288_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5701_ _2422_ _2436_ _2446_ _2454_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__o31a_1
XFILLER_0_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6681_ RF.registers\[8\]\[19\] _3132_ _3242_ VGND VGND VPWR VPWR _3252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5632_ _1168_ _1997_ _2386_ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__o21ba_1
X_8420_ _4190_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8351_ RF.registers\[16\]\[19\] _3495_ _4144_ VGND VGND VPWR VPWR _4154_ sky130_fd_sc_hd__mux2_1
X_5563_ RF.registers\[4\]\[5\] RF.registers\[5\]\[5\] RF.registers\[6\]\[5\] RF.registers\[7\]\[5\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2319_ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4514_ RF.registers\[12\]\[21\] RF.registers\[13\]\[21\] RF.registers\[14\]\[21\]
+ RF.registers\[15\]\[21\] _1267_ _1268_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7302_ _3035_ RF.registers\[31\]\[6\] _3591_ VGND VGND VPWR VPWR _3598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8282_ _4117_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__clkbuf_1
X_5494_ _2213_ _2249_ _2178_ VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4445_ _1200_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7233_ _3561_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7164_ RF.registers\[7\]\[6\] _3468_ _3517_ VGND VGND VPWR VPWR _3524_ sky130_fd_sc_hd__mux2_1
X_4376_ RF.registers\[28\]\[1\] RF.registers\[29\]\[1\] RF.registers\[30\]\[1\] RF.registers\[31\]\[1\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__mux4_1
X_6115_ _2778_ _2848_ _1879_ VGND VGND VPWR VPWR _2849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7095_ net17 VGND VGND VPWR VPWR _3481_ sky130_fd_sc_hd__buf_2
X_6046_ _1618_ _2782_ VGND VGND VPWR VPWR _2783_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_68_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7997_ _3966_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ RF.registers\[4\]\[16\] _3126_ _3387_ VGND VGND VPWR VPWR _3394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6879_ _3357_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8618_ clknet_leaf_10_CLK _0802_ VGND VGND VPWR VPWR RF.registers\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8549_ _4258_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7920_ _3925_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__clkbuf_1
X_7851_ _3109_ RF.registers\[23\]\[8\] _3880_ VGND VGND VPWR VPWR _3889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6802_ RF.registers\[6\]\[11\] _3116_ _3315_ VGND VGND VPWR VPWR _3317_ sky130_fd_sc_hd__mux2_1
X_4994_ RF.registers\[4\]\[22\] RF.registers\[5\]\[22\] RF.registers\[6\]\[22\] RF.registers\[7\]\[22\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__mux4_1
X_7782_ _3852_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9521_ clknet_leaf_13_CLK _0681_ VGND VGND VPWR VPWR RF.registers\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6733_ _3046_ RF.registers\[14\]\[11\] _3278_ VGND VGND VPWR VPWR _3280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6664_ _3243_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__clkbuf_1
X_9452_ clknet_leaf_87_CLK _0612_ VGND VGND VPWR VPWR RF.registers\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5615_ _2363_ _2368_ _2369_ VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__and3b_1
X_8403_ RF.registers\[12\]\[11\] _3479_ _4180_ VGND VGND VPWR VPWR _4182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9383_ clknet_leaf_58_CLK _0543_ VGND VGND VPWR VPWR RF.registers\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6595_ _3043_ RF.registers\[15\]\[10\] _3206_ VGND VGND VPWR VPWR _3207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5546_ RF.registers\[0\]\[4\] RF.registers\[1\]\[4\] RF.registers\[2\]\[4\] RF.registers\[3\]\[4\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8334_ _4145_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__clkbuf_1
X_5477_ _2231_ _2232_ _1712_ VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__mux2_1
X_8265_ _3113_ RF.registers\[13\]\[10\] _4108_ VGND VGND VPWR VPWR _4109_ sky130_fd_sc_hd__mux2_1
X_7216_ RF.registers\[7\]\[31\] _3452_ _3516_ VGND VGND VPWR VPWR _3551_ sky130_fd_sc_hd__mux2_1
X_4428_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__buf_4
X_8196_ _4060_ VGND VGND VPWR VPWR _4072_ sky130_fd_sc_hd__buf_4
X_7147_ _3514_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4359_ RF.registers\[20\]\[2\] RF.registers\[21\]\[2\] RF.registers\[22\]\[2\] RF.registers\[23\]\[2\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__mux4_1
X_7078_ _3469_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
X_6029_ _1512_ _1602_ _2658_ _2536_ VGND VGND VPWR VPWR _2767_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6380_ _3073_ RF.registers\[22\]\[24\] _3065_ VGND VGND VPWR VPWR _3074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_3_5__leaf_CLK sky130_fd_sc_hd__clkbuf_16
Xclkload22 clknet_leaf_84_CLK VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_11_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload33 clknet_leaf_70_CLK VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__inv_6
Xclkload11 clknet_leaf_93_CLK VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__clkinvlp_2
X_5400_ RF.registers\[8\]\[13\] RF.registers\[9\]\[13\] RF.registers\[10\]\[13\] RF.registers\[11\]\[13\]
+ _1702_ _1678_ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__mux4_1
Xclkload44 clknet_leaf_60_CLK VGND VGND VPWR VPWR clkload44/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload77 clknet_leaf_44_CLK VGND VGND VPWR VPWR clkload77/X sky130_fd_sc_hd__clkbuf_4
Xclkload66 clknet_leaf_22_CLK VGND VGND VPWR VPWR clkload66/Y sky130_fd_sc_hd__inv_6
Xclkload55 clknet_leaf_11_CLK VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5331_ RF.registers\[20\]\[1\] RF.registers\[21\]\[1\] RF.registers\[22\]\[1\] RF.registers\[23\]\[1\]
+ _1673_ _1690_ VGND VGND VPWR VPWR _2087_ sky130_fd_sc_hd__mux4_1
Xclkload88 clknet_leaf_33_CLK VGND VGND VPWR VPWR clkload88/Y sky130_fd_sc_hd__clkinvlp_4
X_8050_ RF.registers\[20\]\[5\] _3466_ _3989_ VGND VGND VPWR VPWR _3995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5262_ RF.registers\[20\]\[24\] RF.registers\[21\]\[24\] RF.registers\[22\]\[24\]
+ RF.registers\[23\]\[24\] _1918_ _1919_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__mux4_1
X_7001_ _3422_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
X_5193_ _1945_ _1946_ _1947_ _1948_ _1889_ _1773_ VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__mux4_2
XFILLER_0_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8952_ clknet_leaf_40_CLK _0112_ VGND VGND VPWR VPWR RF.registers\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_50_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8883_ clknet_leaf_51_CLK _0043_ VGND VGND VPWR VPWR RF.registers\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7903_ RF.registers\[18\]\[0\] _3454_ _3916_ VGND VGND VPWR VPWR _3917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7834_ _3879_ VGND VGND VPWR VPWR _3880_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_19_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7765_ _3003_ _3091_ VGND VGND VPWR VPWR _3843_ sky130_fd_sc_hd__nor2_2
XFILLER_0_117_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9504_ clknet_leaf_73_CLK _0664_ VGND VGND VPWR VPWR RF.registers\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6716_ _3029_ RF.registers\[14\]\[3\] _3267_ VGND VGND VPWR VPWR _3271_ sky130_fd_sc_hd__mux2_1
X_4977_ _1702_ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload5 clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_8
X_7696_ _3806_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9435_ clknet_leaf_44_CLK _0595_ VGND VGND VPWR VPWR RF.registers\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6647_ _3234_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__clkbuf_1
X_9366_ clknet_leaf_48_CLK _0526_ VGND VGND VPWR VPWR RF.registers\[20\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6578_ _3027_ RF.registers\[15\]\[2\] _3195_ VGND VGND VPWR VPWR _3198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8317_ _4136_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5529_ _1828_ _2284_ _1728_ VGND VGND VPWR VPWR _2285_ sky130_fd_sc_hd__a21oi_1
X_9297_ clknet_leaf_19_CLK _0457_ VGND VGND VPWR VPWR RF.registers\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8248_ _3097_ RF.registers\[13\]\[2\] _4097_ VGND VGND VPWR VPWR _4100_ sky130_fd_sc_hd__mux2_1
X_8179_ _4063_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5880_ _2546_ _2570_ _2625_ _2105_ VGND VGND VPWR VPWR _2626_ sky130_fd_sc_hd__a22oi_2
X_4900_ RF.registers\[4\]\[0\] RF.registers\[5\]\[0\] RF.registers\[6\]\[0\] RF.registers\[7\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_36_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4831_ _1215_ _1578_ _1582_ _1586_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7550_ _3729_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4762_ _1516_ _1517_ _1035_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7481_ _3077_ RF.registers\[25\]\[26\] _3686_ VGND VGND VPWR VPWR _3693_ sky130_fd_sc_hd__mux2_1
X_6501_ _3154_ VGND VGND VPWR VPWR _3155_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4693_ RF.registers\[20\]\[12\] RF.registers\[21\]\[12\] RF.registers\[22\]\[12\]
+ RF.registers\[23\]\[12\] _1219_ _1221_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9220_ clknet_leaf_90_CLK _0380_ VGND VGND VPWR VPWR RF.registers\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6432_ RF.registers\[17\]\[8\] _3109_ _3093_ VGND VGND VPWR VPWR _3110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9151_ clknet_leaf_65_CLK _0311_ VGND VGND VPWR VPWR RF.registers\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_8102_ RF.registers\[20\]\[30\] _3450_ _3988_ VGND VGND VPWR VPWR _4022_ sky130_fd_sc_hd__mux2_1
X_6363_ net24 VGND VGND VPWR VPWR _3062_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6294_ _3014_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__clkbuf_1
X_9082_ clknet_leaf_25_CLK _0242_ VGND VGND VPWR VPWR RF.registers\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_58_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5314_ _2068_ _2069_ _1645_ VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__mux2_1
X_5245_ RF.registers\[16\]\[25\] RF.registers\[17\]\[25\] RF.registers\[18\]\[25\]
+ RF.registers\[19\]\[25\] _1822_ _1823_ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__mux4_1
X_8033_ _3015_ RF.registers\[21\]\[30\] _3951_ VGND VGND VPWR VPWR _3985_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5176_ _1930_ _1931_ _1726_ VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8935_ clknet_leaf_59_CLK _0095_ VGND VGND VPWR VPWR RF.registers\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8866_ clknet_leaf_91_CLK _0026_ VGND VGND VPWR VPWR RF.registers\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_7817_ RF.registers\[9\]\[24\] _3506_ _3866_ VGND VGND VPWR VPWR _3871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8797_ clknet_leaf_14_CLK _0981_ VGND VGND VPWR VPWR RF.registers\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_7748_ _3834_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7679_ RF.registers\[2\]\[23\] _3504_ _3794_ VGND VGND VPWR VPWR _3798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9418_ clknet_leaf_82_CLK _0578_ VGND VGND VPWR VPWR RF.registers\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9349_ clknet_leaf_62_CLK _0509_ VGND VGND VPWR VPWR RF.registers\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ RF.registers\[28\]\[20\] RF.registers\[29\]\[20\] RF.registers\[30\]\[20\]
+ RF.registers\[31\]\[20\] _1782_ _1680_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6981_ net10 net9 net46 VGND VGND VPWR VPWR _3411_ sky130_fd_sc_hd__nand3_4
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5932_ _2674_ _2675_ _1147_ VGND VGND VPWR VPWR _2676_ sky130_fd_sc_hd__mux2_1
X_8720_ clknet_leaf_84_CLK _0904_ VGND VGND VPWR VPWR RF.registers\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_124_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5863_ _2565_ _2609_ _1803_ VGND VGND VPWR VPWR _2610_ sky130_fd_sc_hd__mux2_1
X_8651_ clknet_leaf_78_CLK _0835_ VGND VGND VPWR VPWR RF.registers\[0\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_7602_ _3062_ RF.registers\[28\]\[19\] _3747_ VGND VGND VPWR VPWR _3757_ sky130_fd_sc_hd__mux2_1
X_5794_ _2539_ _2540_ _2543_ VGND VGND VPWR VPWR _2544_ sky130_fd_sc_hd__o21ai_1
X_4814_ _1568_ _1569_ _1107_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__mux2_1
X_8582_ clknet_leaf_62_CLK _0766_ VGND VGND VPWR VPWR RF.registers\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7533_ _3720_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
X_4745_ _1499_ _1500_ _1259_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4676_ RF.registers\[16\]\[22\] RF.registers\[17\]\[22\] RF.registers\[18\]\[22\]
+ RF.registers\[19\]\[22\] _1182_ _1184_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7464_ _3060_ RF.registers\[25\]\[18\] _3675_ VGND VGND VPWR VPWR _3684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9203_ clknet_leaf_25_CLK _0363_ VGND VGND VPWR VPWR RF.registers\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7395_ _3647_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6415_ _3098_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9134_ clknet_leaf_5_CLK _0294_ VGND VGND VPWR VPWR RF.registers\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6346_ _3050_ RF.registers\[22\]\[13\] _3044_ VGND VGND VPWR VPWR _3051_ sky130_fd_sc_hd__mux2_1
X_9065_ clknet_leaf_1_CLK _0225_ VGND VGND VPWR VPWR RF.registers\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8016_ _3976_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__clkbuf_1
X_6277_ _2621_ _2995_ _3001_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__o21bai_2
X_5228_ RF.registers\[28\]\[26\] RF.registers\[29\]\[26\] RF.registers\[30\]\[26\]
+ RF.registers\[31\]\[26\] _1881_ _1883_ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__mux4_1
X_5159_ _1913_ _1914_ _1889_ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8918_ clknet_leaf_47_CLK _0078_ VGND VGND VPWR VPWR RF.registers\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8849_ clknet_leaf_55_CLK _0009_ VGND VGND VPWR VPWR RF.registers\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4530_ _1282_ _1285_ _1071_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4461_ _1171_ _1188_ _1216_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6200_ _2621_ _2921_ _2928_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__o21bai_2
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7180_ _3532_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4392_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__clkbuf_4
X_6131_ _2586_ _2797_ VGND VGND VPWR VPWR _2863_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _2040_ _2796_ _2797_ _2421_ VGND VGND VPWR VPWR _2798_ sky130_fd_sc_hd__o31ai_1
X_5013_ RF.registers\[8\]\[21\] RF.registers\[9\]\[21\] RF.registers\[10\]\[21\] RF.registers\[11\]\[21\]
+ _1767_ _1768_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6964_ _3402_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6895_ RF.registers\[5\]\[23\] _3141_ _3362_ VGND VGND VPWR VPWR _3366_ sky130_fd_sc_hd__mux2_1
X_5915_ _1464_ _2536_ _2658_ VGND VGND VPWR VPWR _2659_ sky130_fd_sc_hd__or3_1
X_8703_ clknet_leaf_65_CLK _0887_ VGND VGND VPWR VPWR RF.registers\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8634_ clknet_leaf_29_CLK _0818_ VGND VGND VPWR VPWR RF.registers\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5846_ _1060_ _1083_ VGND VGND VPWR VPWR _2594_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8565_ _4266_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__clkbuf_1
X_5777_ _2524_ _2527_ _2501_ VGND VGND VPWR VPWR _2528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8496_ RF.registers\[11\]\[23\] net29 _4227_ VGND VGND VPWR VPWR _4231_ sky130_fd_sc_hd__mux2_1
X_7516_ _3043_ RF.registers\[27\]\[10\] _3711_ VGND VGND VPWR VPWR _3712_ sky130_fd_sc_hd__mux2_1
X_4728_ RF.registers\[20\]\[14\] RF.registers\[21\]\[14\] RF.registers\[22\]\[14\]
+ RF.registers\[23\]\[14\] _1324_ _1325_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7447_ _3663_ VGND VGND VPWR VPWR _3675_ sky130_fd_sc_hd__buf_4
X_4659_ _1025_ _1406_ _1410_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7378_ _3638_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9117_ clknet_leaf_22_CLK _0277_ VGND VGND VPWR VPWR RF.registers\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6329_ net44 VGND VGND VPWR VPWR _3039_ sky130_fd_sc_hd__clkbuf_2
X_9048_ clknet_leaf_38_CLK _0208_ VGND VGND VPWR VPWR RF.registers\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5700_ _2452_ _2453_ _2421_ VGND VGND VPWR VPWR _2454_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6680_ _3251_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5631_ _1167_ _2016_ VGND VGND VPWR VPWR _2386_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8350_ _4153_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__clkbuf_1
X_5562_ _1716_ _2317_ VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__nor2_1
X_4513_ RF.registers\[8\]\[21\] RF.registers\[9\]\[21\] RF.registers\[10\]\[21\] RF.registers\[11\]\[21\]
+ _1267_ _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8281_ _3130_ RF.registers\[13\]\[18\] _4108_ VGND VGND VPWR VPWR _4117_ sky130_fd_sc_hd__mux2_1
X_7301_ _3597_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5493_ _1669_ _2230_ _2248_ VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__o21ai_1
X_7232_ _3033_ RF.registers\[29\]\[5\] _3555_ VGND VGND VPWR VPWR _3561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4444_ _1027_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__buf_4
XFILLER_0_111_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7163_ _3523_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
X_4375_ _1129_ _1130_ _1035_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__mux2_1
X_6114_ _2800_ _2847_ _1877_ VGND VGND VPWR VPWR _2848_ sky130_fd_sc_hd__mux2_1
X_7094_ _3480_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
X_6045_ _1512_ _1602_ _1634_ _2658_ _2536_ VGND VGND VPWR VPWR _2782_ sky130_fd_sc_hd__a41o_1
XFILLER_0_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7996_ _3118_ RF.registers\[21\]\[12\] _3963_ VGND VGND VPWR VPWR _3966_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6947_ _3393_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6878_ RF.registers\[5\]\[15\] _3124_ _3351_ VGND VGND VPWR VPWR _3357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5829_ _2418_ VGND VGND VPWR VPWR _2577_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8617_ clknet_leaf_9_CLK _0801_ VGND VGND VPWR VPWR RF.registers\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8548_ RF.registers\[10\]\[16\] net21 _4255_ VGND VGND VPWR VPWR _4258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_680 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8479_ RF.registers\[11\]\[15\] net20 _4216_ VGND VGND VPWR VPWR _4222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7850_ _3888_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__clkbuf_1
X_6801_ _3316_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4993_ _1745_ _1746_ _1748_ _1697_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7781_ RF.registers\[9\]\[7\] _3470_ _3844_ VGND VGND VPWR VPWR _3852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9520_ clknet_leaf_12_CLK _0680_ VGND VGND VPWR VPWR RF.registers\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6732_ _3279_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__clkbuf_1
X_6663_ RF.registers\[8\]\[10\] _3113_ _3242_ VGND VGND VPWR VPWR _3243_ sky130_fd_sc_hd__mux2_1
X_9451_ clknet_leaf_86_CLK _0611_ VGND VGND VPWR VPWR RF.registers\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5614_ _1799_ _2306_ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__or2_1
X_8402_ _4181_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9382_ clknet_leaf_62_CLK _0542_ VGND VGND VPWR VPWR RF.registers\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6594_ _3194_ VGND VGND VPWR VPWR _3206_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5545_ RF.registers\[4\]\[4\] RF.registers\[5\]\[4\] RF.registers\[6\]\[4\] RF.registers\[7\]\[4\]
+ _1718_ _1679_ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__mux4_1
X_8333_ RF.registers\[16\]\[10\] _3476_ _4144_ VGND VGND VPWR VPWR _4145_ sky130_fd_sc_hd__mux2_1
X_5476_ RF.registers\[28\]\[9\] RF.registers\[29\]\[9\] RF.registers\[30\]\[9\] RF.registers\[31\]\[9\]
+ _1675_ _1692_ VGND VGND VPWR VPWR _2232_ sky130_fd_sc_hd__mux4_1
X_8264_ _4096_ VGND VGND VPWR VPWR _4108_ sky130_fd_sc_hd__buf_4
X_7215_ _3550_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_4427_ _1044_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__clkbuf_4
X_8195_ _4071_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7146_ RF.registers\[19\]\[30\] _3450_ _3455_ VGND VGND VPWR VPWR _3514_ sky130_fd_sc_hd__mux2_1
X_4358_ RF.registers\[16\]\[2\] RF.registers\[17\]\[2\] RF.registers\[18\]\[2\] RF.registers\[19\]\[2\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__mux4_1
X_4289_ RF.registers\[4\]\[4\] RF.registers\[5\]\[4\] RF.registers\[6\]\[4\] RF.registers\[7\]\[4\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__mux4_1
X_7077_ RF.registers\[19\]\[6\] _3468_ _3456_ VGND VGND VPWR VPWR _3469_ sky130_fd_sc_hd__mux2_1
X_6028_ _2755_ _2760_ _2766_ _2621_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__o22a_1
XFILLER_0_96_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7979_ _3101_ RF.registers\[21\]\[4\] _3952_ VGND VGND VPWR VPWR _3957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload12 clknet_leaf_94_CLK VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_4
Xclkload34 clknet_leaf_71_CLK VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__clkinv_4
Xclkload23 clknet_leaf_85_CLK VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__inv_6
Xclkload78 clknet_leaf_45_CLK VGND VGND VPWR VPWR clkload78/Y sky130_fd_sc_hd__clkinv_4
Xclkload67 clknet_leaf_23_CLK VGND VGND VPWR VPWR clkload67/X sky130_fd_sc_hd__clkbuf_4
Xclkload56 clknet_leaf_12_CLK VGND VGND VPWR VPWR clkload56/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5330_ RF.registers\[16\]\[1\] RF.registers\[17\]\[1\] RF.registers\[18\]\[1\] RF.registers\[19\]\[1\]
+ _1673_ _1690_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__mux4_1
Xclkload45 clknet_leaf_61_CLK VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload89 clknet_leaf_34_CLK VGND VGND VPWR VPWR clkload89/X sky130_fd_sc_hd__clkbuf_4
X_5261_ _1668_ _2016_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7000_ RF.registers\[3\]\[8\] _3109_ _3413_ VGND VGND VPWR VPWR _3422_ sky130_fd_sc_hd__mux2_1
X_5192_ RF.registers\[20\]\[28\] RF.registers\[21\]\[28\] RF.registers\[22\]\[28\]
+ RF.registers\[23\]\[28\] _1882_ _1884_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__mux4_1
X_8951_ clknet_leaf_49_CLK _0111_ VGND VGND VPWR VPWR RF.registers\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_7902_ _3915_ VGND VGND VPWR VPWR _3916_ sky130_fd_sc_hd__buf_6
XFILLER_0_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8882_ clknet_leaf_54_CLK _0042_ VGND VGND VPWR VPWR RF.registers\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7833_ _3021_ _3193_ VGND VGND VPWR VPWR _3879_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_19_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7764_ _3842_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4976_ _1639_ _1731_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__or2_1
X_6715_ _3270_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__clkbuf_1
X_9503_ clknet_leaf_65_CLK _0663_ VGND VGND VPWR VPWR RF.registers\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7695_ RF.registers\[2\]\[31\] _3452_ _3771_ VGND VGND VPWR VPWR _3806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload6 clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_4
X_9434_ clknet_leaf_35_CLK _0594_ VGND VGND VPWR VPWR RF.registers\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6646_ RF.registers\[8\]\[2\] _3097_ _3231_ VGND VGND VPWR VPWR _3234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9365_ clknet_leaf_29_CLK _0525_ VGND VGND VPWR VPWR RF.registers\[20\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6577_ _3197_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8316_ RF.registers\[16\]\[2\] _3460_ _4133_ VGND VGND VPWR VPWR _4136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5528_ _2282_ _2283_ _1738_ VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9296_ clknet_leaf_7_CLK _0456_ VGND VGND VPWR VPWR RF.registers\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8247_ _4099_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__clkbuf_1
X_5459_ RF.registers\[16\]\[8\] RF.registers\[17\]\[8\] RF.registers\[18\]\[8\] RF.registers\[19\]\[8\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2215_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8178_ RF.registers\[1\]\[1\] _3458_ _4061_ VGND VGND VPWR VPWR _4063_ sky130_fd_sc_hd__mux2_1
X_7129_ net29 VGND VGND VPWR VPWR _3504_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_38_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_70_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_70_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4830_ _1205_ _1585_ _1170_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4761_ RF.registers\[24\]\[8\] RF.registers\[25\]\[8\] RF.registers\[26\]\[8\] RF.registers\[27\]\[8\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7480_ _3692_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
X_4692_ _1416_ _1447_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__or2b_1
X_6500_ net10 net9 net46 VGND VGND VPWR VPWR _3154_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6431_ net44 VGND VGND VPWR VPWR _3109_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_113_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6362_ _3061_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__clkbuf_1
X_9150_ clknet_leaf_67_CLK _0310_ VGND VGND VPWR VPWR RF.registers\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8101_ _4021_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__clkbuf_1
X_5313_ RF.registers\[24\]\[2\] RF.registers\[25\]\[2\] RF.registers\[26\]\[2\] RF.registers\[27\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2069_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_61_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_61_CLK sky130_fd_sc_hd__clkbuf_8
X_9081_ clknet_leaf_27_CLK _0241_ VGND VGND VPWR VPWR RF.registers\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6293_ RF.registers\[10\]\[29\] _3013_ _3007_ VGND VGND VPWR VPWR _3014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5244_ RF.registers\[20\]\[25\] RF.registers\[21\]\[25\] RF.registers\[22\]\[25\]
+ RF.registers\[23\]\[25\] _1822_ _1823_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__mux4_1
X_8032_ _3984_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__clkbuf_1
X_5175_ RF.registers\[24\]\[29\] RF.registers\[25\]\[29\] RF.registers\[26\]\[29\]
+ RF.registers\[27\]\[29\] _1705_ _1708_ VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8934_ clknet_leaf_61_CLK _0094_ VGND VGND VPWR VPWR RF.registers\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8865_ clknet_leaf_72_CLK _0025_ VGND VGND VPWR VPWR RF.registers\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_7816_ _3870_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8796_ clknet_leaf_16_CLK _0980_ VGND VGND VPWR VPWR RF.registers\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7747_ _3071_ RF.registers\[30\]\[23\] _3830_ VGND VGND VPWR VPWR _3834_ sky130_fd_sc_hd__mux2_1
X_4959_ _1700_ _1714_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7678_ _3797_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6629_ _3224_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__clkbuf_1
X_9417_ clknet_leaf_86_CLK _0577_ VGND VGND VPWR VPWR RF.registers\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9348_ clknet_leaf_95_CLK _0508_ VGND VGND VPWR VPWR RF.registers\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9279_ clknet_leaf_72_CLK _0439_ VGND VGND VPWR VPWR RF.registers\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_528 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_43_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_43_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6980_ _3410_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5931_ _1800_ _2194_ _2176_ VGND VGND VPWR VPWR _2675_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5862_ _2353_ _2358_ VGND VGND VPWR VPWR _2609_ sky130_fd_sc_hd__and2_1
X_8650_ clknet_leaf_82_CLK _0834_ VGND VGND VPWR VPWR RF.registers\[0\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_7601_ _3756_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
X_5793_ _2511_ _2512_ _2518_ _2542_ VGND VGND VPWR VPWR _2543_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_8_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4813_ RF.registers\[0\]\[11\] RF.registers\[1\]\[11\] RF.registers\[2\]\[11\] RF.registers\[3\]\[11\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__mux4_1
X_8581_ clknet_leaf_59_CLK _0765_ VGND VGND VPWR VPWR RF.registers\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7532_ _3060_ RF.registers\[27\]\[18\] _3711_ VGND VGND VPWR VPWR _3720_ sky130_fd_sc_hd__mux2_1
X_4744_ RF.registers\[24\]\[15\] RF.registers\[25\]\[15\] RF.registers\[26\]\[15\]
+ RF.registers\[27\]\[15\] _1324_ _1325_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4675_ RF.registers\[20\]\[22\] RF.registers\[21\]\[22\] RF.registers\[22\]\[22\]
+ RF.registers\[23\]\[22\] _1182_ _1184_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__mux4_1
XFILLER_0_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9202_ clknet_leaf_42_CLK _0362_ VGND VGND VPWR VPWR RF.registers\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_7463_ _3683_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_34_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_34_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7394_ _3058_ RF.registers\[26\]\[17\] _3639_ VGND VGND VPWR VPWR _3647_ sky130_fd_sc_hd__mux2_1
X_6414_ RF.registers\[17\]\[2\] _3097_ _3093_ VGND VGND VPWR VPWR _3098_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6345_ net18 VGND VGND VPWR VPWR _3050_ sky130_fd_sc_hd__buf_2
X_9133_ clknet_leaf_2_CLK _0293_ VGND VGND VPWR VPWR RF.registers\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6276_ _2720_ _2737_ _2996_ _2472_ _3000_ VGND VGND VPWR VPWR _3001_ sky130_fd_sc_hd__a221o_1
X_9064_ clknet_leaf_1_CLK _0224_ VGND VGND VPWR VPWR RF.registers\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8015_ _3137_ RF.registers\[21\]\[21\] _3974_ VGND VGND VPWR VPWR _3976_ sky130_fd_sc_hd__mux2_1
X_5227_ _1981_ _1982_ _1901_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5158_ RF.registers\[12\]\[30\] RF.registers\[13\]\[30\] RF.registers\[14\]\[30\]
+ RF.registers\[15\]\[30\] _1881_ _1883_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5089_ _1843_ _1844_ _1686_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__mux2_1
X_8917_ clknet_leaf_28_CLK _0077_ VGND VGND VPWR VPWR RF.registers\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8848_ clknet_leaf_55_CLK _0008_ VGND VGND VPWR VPWR RF.registers\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8779_ clknet_leaf_82_CLK _0963_ VGND VGND VPWR VPWR RF.registers\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_25_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4460_ _1197_ _1206_ _1212_ _1214_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_16_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_16_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4391_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6130_ _2621_ _2856_ _2862_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_55_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _2737_ VGND VGND VPWR VPWR _2797_ sky130_fd_sc_hd__inv_2
X_5012_ _1707_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6963_ RF.registers\[4\]\[23\] _3141_ _3398_ VGND VGND VPWR VPWR _3402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6894_ _3365_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5914_ _2657_ VGND VGND VPWR VPWR _2658_ sky130_fd_sc_hd__buf_2
X_8702_ clknet_leaf_67_CLK _0886_ VGND VGND VPWR VPWR RF.registers\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8633_ clknet_leaf_30_CLK _0817_ VGND VGND VPWR VPWR RF.registers\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5845_ _1111_ _1125_ _1145_ _1166_ VGND VGND VPWR VPWR _2593_ sky130_fd_sc_hd__nand4_2
XFILLER_0_118_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8564_ RF.registers\[10\]\[24\] net30 _3006_ VGND VGND VPWR VPWR _4266_ sky130_fd_sc_hd__mux2_1
X_5776_ _2363_ _2456_ _2526_ VGND VGND VPWR VPWR _2527_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8495_ _4230_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__clkbuf_1
X_7515_ _3699_ VGND VGND VPWR VPWR _3711_ sky130_fd_sc_hd__buf_4
XFILLER_0_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ RF.registers\[16\]\[14\] RF.registers\[17\]\[14\] RF.registers\[18\]\[14\]
+ RF.registers\[19\]\[14\] _1324_ _1325_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__mux4_1
X_7446_ _3674_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4658_ _1078_ _1413_ _1057_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4589_ RF.registers\[0\]\[30\] RF.registers\[1\]\[30\] RF.registers\[2\]\[30\] RF.registers\[3\]\[30\]
+ _1262_ _1263_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__mux4_1
X_9116_ clknet_leaf_22_CLK _0276_ VGND VGND VPWR VPWR RF.registers\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_7377_ _3041_ RF.registers\[26\]\[9\] _3628_ VGND VGND VPWR VPWR _3638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6328_ _3038_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__clkbuf_1
X_9047_ clknet_leaf_31_CLK _0207_ VGND VGND VPWR VPWR RF.registers\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6259_ _1923_ _2983_ VGND VGND VPWR VPWR _2985_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_4_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_5_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5630_ _2383_ _2384_ VGND VGND VPWR VPWR _2385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5561_ _2315_ _2316_ _1711_ VGND VGND VPWR VPWR _2317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4512_ _1202_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8280_ _4116_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__clkbuf_1
X_5492_ _1668_ _2247_ VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__nand2_1
X_7300_ _3033_ RF.registers\[31\]\[5\] _3591_ VGND VGND VPWR VPWR _3597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7231_ _3560_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4443_ _1198_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7162_ RF.registers\[7\]\[5\] _3466_ _3517_ VGND VGND VPWR VPWR _3523_ sky130_fd_sc_hd__mux2_1
X_4374_ RF.registers\[16\]\[1\] RF.registers\[17\]\[1\] RF.registers\[18\]\[1\] RF.registers\[19\]\[1\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__mux4_1
X_6113_ _1781_ _1756_ VGND VGND VPWR VPWR _2847_ sky130_fd_sc_hd__and2_1
X_7093_ RF.registers\[19\]\[11\] _3479_ _3477_ VGND VGND VPWR VPWR _3480_ sky130_fd_sc_hd__mux2_1
X_6044_ _2408_ _2775_ _2776_ _2781_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_68_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7995_ _3965_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6946_ RF.registers\[4\]\[15\] _3124_ _3387_ VGND VGND VPWR VPWR _3393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6877_ _3356_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5828_ _2504_ _2564_ _2576_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__a21o_1
XFILLER_0_8_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8616_ clknet_leaf_96_CLK _0800_ VGND VGND VPWR VPWR RF.registers\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8547_ _4257_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__clkbuf_1
X_5759_ _2509_ _2510_ VGND VGND VPWR VPWR _2511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8478_ _4221_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7429_ _3025_ RF.registers\[25\]\[1\] _3664_ VGND VGND VPWR VPWR _3666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6800_ RF.registers\[6\]\[10\] _3113_ _3315_ VGND VGND VPWR VPWR _3316_ sky130_fd_sc_hd__mux2_1
X_4992_ _1712_ _1747_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7780_ _3851_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6731_ _3043_ RF.registers\[14\]\[10\] _3278_ VGND VGND VPWR VPWR _3279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6662_ _3230_ VGND VGND VPWR VPWR _3242_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9450_ clknet_leaf_86_CLK _0610_ VGND VGND VPWR VPWR RF.registers\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_5613_ _1167_ _2063_ VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8401_ RF.registers\[12\]\[10\] _3476_ _4180_ VGND VGND VPWR VPWR _4181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9381_ clknet_leaf_59_CLK _0541_ VGND VGND VPWR VPWR RF.registers\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8332_ _4132_ VGND VGND VPWR VPWR _4144_ sky130_fd_sc_hd__buf_4
X_6593_ _3205_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__clkbuf_1
X_5544_ _1716_ _2299_ VGND VGND VPWR VPWR _2300_ sky130_fd_sc_hd__nor2_1
X_5475_ RF.registers\[24\]\[9\] RF.registers\[25\]\[9\] RF.registers\[26\]\[9\] RF.registers\[27\]\[9\]
+ _1675_ _1692_ VGND VGND VPWR VPWR _2231_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8263_ _4107_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__clkbuf_1
X_7214_ RF.registers\[7\]\[30\] _3450_ _3516_ VGND VGND VPWR VPWR _3550_ sky130_fd_sc_hd__mux2_1
X_4426_ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8194_ RF.registers\[1\]\[9\] _3474_ _4061_ VGND VGND VPWR VPWR _4071_ sky130_fd_sc_hd__mux2_1
X_7145_ _3513_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4357_ RF.registers\[28\]\[2\] RF.registers\[29\]\[2\] RF.registers\[30\]\[2\] RF.registers\[31\]\[2\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__mux4_1
X_4288_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__buf_4
X_7076_ net42 VGND VGND VPWR VPWR _3468_ sky130_fd_sc_hd__buf_2
X_6027_ _2763_ _2765_ VGND VGND VPWR VPWR _2766_ sky130_fd_sc_hd__xnor2_1
X_7978_ _3956_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6929_ RF.registers\[4\]\[7\] _3107_ _3376_ VGND VGND VPWR VPWR _3384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9579_ clknet_leaf_89_CLK _0739_ VGND VGND VPWR VPWR RF.registers\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload13 clknet_leaf_95_CLK VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__bufinv_16
Xclkload35 clknet_leaf_72_CLK VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__clkinvlp_2
Xclkload24 clknet_leaf_86_CLK VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__clkinv_4
Xclkload68 clknet_leaf_24_CLK VGND VGND VPWR VPWR clkload68/Y sky130_fd_sc_hd__inv_6
Xclkload57 clknet_leaf_13_CLK VGND VGND VPWR VPWR clkload57/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload46 clknet_leaf_62_CLK VGND VGND VPWR VPWR clkload46/Y sky130_fd_sc_hd__inv_6
XFILLER_0_121_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload79 clknet_leaf_51_CLK VGND VGND VPWR VPWR clkload79/Y sky130_fd_sc_hd__inv_8
X_5260_ _1638_ _2015_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5191_ RF.registers\[16\]\[28\] RF.registers\[17\]\[28\] RF.registers\[18\]\[28\]
+ RF.registers\[19\]\[28\] _1882_ _1884_ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__mux4_1
X_8950_ clknet_leaf_48_CLK _0110_ VGND VGND VPWR VPWR RF.registers\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_7901_ _3005_ _3090_ VGND VGND VPWR VPWR _3915_ sky130_fd_sc_hd__nor2_2
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8881_ clknet_leaf_56_CLK _0041_ VGND VGND VPWR VPWR RF.registers\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_7832_ _3878_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4975_ _1672_ _1698_ _1715_ _1730_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__a2bb2o_2
X_7763_ _3087_ RF.registers\[30\]\[31\] _3807_ VGND VGND VPWR VPWR _3842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9502_ clknet_leaf_68_CLK _0662_ VGND VGND VPWR VPWR RF.registers\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6714_ _3027_ RF.registers\[14\]\[2\] _3267_ VGND VGND VPWR VPWR _3270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9433_ clknet_leaf_49_CLK _0593_ VGND VGND VPWR VPWR RF.registers\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_7694_ _3805_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload7 clknet_leaf_0_CLK VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinv_4
X_6645_ _3233_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9364_ clknet_leaf_37_CLK _0524_ VGND VGND VPWR VPWR RF.registers\[20\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6576_ _3025_ RF.registers\[15\]\[1\] _3195_ VGND VGND VPWR VPWR _3197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9295_ clknet_leaf_4_CLK _0455_ VGND VGND VPWR VPWR RF.registers\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8315_ _4135_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5527_ RF.registers\[0\]\[7\] RF.registers\[1\]\[7\] RF.registers\[2\]\[7\] RF.registers\[3\]\[7\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8246_ _3095_ RF.registers\[13\]\[1\] _4097_ VGND VGND VPWR VPWR _4099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5458_ RF.registers\[20\]\[8\] RF.registers\[21\]\[8\] RF.registers\[22\]\[8\] RF.registers\[23\]\[8\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2214_ sky130_fd_sc_hd__mux4_1
X_8177_ _4062_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__clkbuf_1
X_4409_ _1088_ _1164_ net8 VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a21oi_2
X_5389_ RF.registers\[20\]\[13\] RF.registers\[21\]\[13\] RF.registers\[22\]\[13\]
+ RF.registers\[23\]\[13\] _1673_ _1690_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__mux4_1
X_7128_ _3503_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7059_ RF.registers\[19\]\[0\] _3454_ _3456_ VGND VGND VPWR VPWR _3457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ RF.registers\[28\]\[8\] RF.registers\[29\]\[8\] RF.registers\[30\]\[8\] RF.registers\[31\]\[8\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4691_ _1430_ _1446_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6430_ _3108_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6361_ _3060_ RF.registers\[22\]\[18\] _3044_ VGND VGND VPWR VPWR _3061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8100_ RF.registers\[20\]\[29\] _3448_ _4011_ VGND VGND VPWR VPWR _4021_ sky130_fd_sc_hd__mux2_1
X_5312_ RF.registers\[28\]\[2\] RF.registers\[29\]\[2\] RF.registers\[30\]\[2\] RF.registers\[31\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6292_ net35 VGND VGND VPWR VPWR _3013_ sky130_fd_sc_hd__buf_2
X_9080_ clknet_leaf_38_CLK _0240_ VGND VGND VPWR VPWR RF.registers\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8031_ _3013_ RF.registers\[21\]\[29\] _3974_ VGND VGND VPWR VPWR _3984_ sky130_fd_sc_hd__mux2_1
X_5243_ _1980_ _1998_ VGND VGND VPWR VPWR _1999_ sky130_fd_sc_hd__or2_1
X_5174_ RF.registers\[28\]\[29\] RF.registers\[29\]\[29\] RF.registers\[30\]\[29\]
+ RF.registers\[31\]\[29\] _1705_ _1708_ VGND VGND VPWR VPWR _1930_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8933_ clknet_leaf_81_CLK _0093_ VGND VGND VPWR VPWR RF.registers\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8864_ clknet_leaf_69_CLK _0024_ VGND VGND VPWR VPWR RF.registers\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_7815_ RF.registers\[9\]\[23\] _3504_ _3866_ VGND VGND VPWR VPWR _3870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8795_ clknet_leaf_44_CLK _0979_ VGND VGND VPWR VPWR RF.registers\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4958_ _1709_ _1710_ _1713_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__mux2_1
X_7746_ _3833_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7677_ RF.registers\[2\]\[22\] _3502_ _3794_ VGND VGND VPWR VPWR _3797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4889_ net3 VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6628_ _3077_ RF.registers\[15\]\[26\] _3217_ VGND VGND VPWR VPWR _3224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9416_ clknet_leaf_78_CLK _0576_ VGND VGND VPWR VPWR RF.registers\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9347_ clknet_leaf_75_CLK _0507_ VGND VGND VPWR VPWR RF.registers\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6559_ _3186_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9278_ clknet_leaf_68_CLK _0438_ VGND VGND VPWR VPWR RF.registers\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8229_ _4089_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5930_ _2212_ _2429_ VGND VGND VPWR VPWR _2674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5861_ _2457_ _2525_ _1877_ VGND VGND VPWR VPWR _2608_ sky130_fd_sc_hd__mux2_1
X_7600_ _3060_ RF.registers\[28\]\[18\] _3747_ VGND VGND VPWR VPWR _3756_ sky130_fd_sc_hd__mux2_1
X_5792_ _2509_ _2541_ _2517_ VGND VGND VPWR VPWR _2542_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_1_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8580_ clknet_leaf_94_CLK _0764_ VGND VGND VPWR VPWR RF.registers\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4812_ RF.registers\[4\]\[11\] RF.registers\[5\]\[11\] RF.registers\[6\]\[11\] RF.registers\[7\]\[11\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7531_ _3719_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
X_4743_ RF.registers\[28\]\[15\] RF.registers\[29\]\[15\] RF.registers\[30\]\[15\]
+ RF.registers\[31\]\[15\] _1262_ _1263_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7462_ _3058_ RF.registers\[25\]\[17\] _3675_ VGND VGND VPWR VPWR _3683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4674_ _1239_ _1421_ _1425_ _1429_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9201_ clknet_leaf_6_CLK _0361_ VGND VGND VPWR VPWR RF.registers\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6413_ net36 VGND VGND VPWR VPWR _3097_ sky130_fd_sc_hd__buf_2
XFILLER_0_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7393_ _3646_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9132_ clknet_leaf_1_CLK _0292_ VGND VGND VPWR VPWR RF.registers\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6344_ _3049_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__clkbuf_1
X_6275_ _2530_ _2859_ _2999_ _1087_ VGND VGND VPWR VPWR _3000_ sky130_fd_sc_hd__o211a_1
X_9063_ clknet_leaf_58_CLK _0223_ VGND VGND VPWR VPWR RF.registers\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5226_ RF.registers\[16\]\[26\] RF.registers\[17\]\[26\] RF.registers\[18\]\[26\]
+ RF.registers\[19\]\[26\] _1881_ _1883_ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__mux4_1
X_8014_ _3975_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_47_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5157_ RF.registers\[8\]\[30\] RF.registers\[9\]\[30\] RF.registers\[10\]\[30\] RF.registers\[11\]\[30\]
+ _1881_ _1883_ VGND VGND VPWR VPWR _1913_ sky130_fd_sc_hd__mux4_1
X_5088_ RF.registers\[16\]\[17\] RF.registers\[17\]\[17\] RF.registers\[18\]\[17\]
+ RF.registers\[19\]\[17\] _1689_ _1693_ VGND VGND VPWR VPWR _1844_ sky130_fd_sc_hd__mux4_1
X_8916_ clknet_leaf_24_CLK _0076_ VGND VGND VPWR VPWR RF.registers\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8847_ clknet_leaf_57_CLK _0007_ VGND VGND VPWR VPWR RF.registers\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_56_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8778_ clknet_leaf_82_CLK _0962_ VGND VGND VPWR VPWR RF.registers\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7729_ _3824_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4390_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6060_ _2585_ _2578_ _2426_ VGND VGND VPWR VPWR _2796_ sky130_fd_sc_hd__mux2_1
X_5011_ _1704_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6962_ _3401_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
X_6893_ RF.registers\[5\]\[22\] _3139_ _3362_ VGND VGND VPWR VPWR _3365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8701_ clknet_leaf_17_CLK _0885_ VGND VGND VPWR VPWR RF.registers\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5913_ _1416_ _1573_ _2506_ _2535_ VGND VGND VPWR VPWR _2657_ sky130_fd_sc_hd__and4b_1
XFILLER_0_118_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8632_ clknet_leaf_38_CLK _0816_ VGND VGND VPWR VPWR RF.registers\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5844_ _2038_ _2590_ _2591_ _2253_ VGND VGND VPWR VPWR _2592_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_66_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8563_ _4265_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5775_ _2327_ _2525_ VGND VGND VPWR VPWR _2526_ sky130_fd_sc_hd__nand2_1
X_7514_ _3710_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
X_8494_ RF.registers\[11\]\[22\] net28 _4227_ VGND VGND VPWR VPWR _4230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4726_ RF.registers\[28\]\[14\] RF.registers\[29\]\[14\] RF.registers\[30\]\[14\]
+ RF.registers\[31\]\[14\] _1324_ _1325_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7445_ _3041_ RF.registers\[25\]\[9\] _3664_ VGND VGND VPWR VPWR _3674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4657_ _1411_ _1412_ _1040_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7376_ _3637_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
X_9115_ clknet_leaf_35_CLK _0275_ VGND VGND VPWR VPWR RF.registers\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4588_ RF.registers\[4\]\[30\] RF.registers\[5\]\[30\] RF.registers\[6\]\[30\] RF.registers\[7\]\[30\]
+ _1262_ _1263_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__mux4_1
X_6327_ _3037_ RF.registers\[22\]\[7\] _3023_ VGND VGND VPWR VPWR _3038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9046_ clknet_leaf_33_CLK _0206_ VGND VGND VPWR VPWR RF.registers\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6258_ _1923_ _2983_ VGND VGND VPWR VPWR _2984_ sky130_fd_sc_hd__nor2_1
X_5209_ _1963_ _1964_ _1745_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__mux2_1
X_6189_ _2916_ _2917_ VGND VGND VPWR VPWR _2918_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5560_ RF.registers\[12\]\[5\] RF.registers\[13\]\[5\] RF.registers\[14\]\[5\] RF.registers\[15\]\[5\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2316_ sky130_fd_sc_hd__mux4_1
X_4511_ _1200_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5491_ _1842_ _2246_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7230_ _3031_ RF.registers\[29\]\[4\] _3555_ VGND VGND VPWR VPWR _3560_ sky130_fd_sc_hd__mux2_1
X_4442_ _1040_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__buf_4
XFILLER_0_111_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7161_ _3522_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4373_ RF.registers\[20\]\[1\] RF.registers\[21\]\[1\] RF.registers\[22\]\[1\] RF.registers\[23\]\[1\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6112_ _2102_ _2554_ VGND VGND VPWR VPWR _2846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7092_ net16 VGND VGND VPWR VPWR _3479_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6043_ _2625_ _2731_ _2779_ _2496_ _2780_ VGND VGND VPWR VPWR _2781_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_68_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7994_ _3116_ RF.registers\[21\]\[11\] _3963_ VGND VGND VPWR VPWR _3965_ sky130_fd_sc_hd__mux2_1
X_6945_ _3392_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6876_ RF.registers\[5\]\[14\] _3122_ _3351_ VGND VGND VPWR VPWR _3356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5827_ _2496_ _2569_ _2572_ _2468_ _2575_ VGND VGND VPWR VPWR _2576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8615_ clknet_leaf_83_CLK _0799_ VGND VGND VPWR VPWR RF.registers\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5758_ _2305_ _2508_ VGND VGND VPWR VPWR _2510_ sky130_fd_sc_hd__and2_1
X_8546_ RF.registers\[10\]\[15\] net20 _4255_ VGND VGND VPWR VPWR _4257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4709_ RF.registers\[20\]\[13\] RF.registers\[21\]\[13\] RF.registers\[22\]\[13\]
+ RF.registers\[23\]\[13\] _1027_ _1029_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__mux4_1
X_8477_ RF.registers\[11\]\[14\] net19 _4216_ VGND VGND VPWR VPWR _4221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5689_ _1961_ _1999_ _2347_ VGND VGND VPWR VPWR _2443_ sky130_fd_sc_hd__mux2_1
X_7428_ _3665_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_79_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7359_ _3019_ RF.registers\[26\]\[0\] _3628_ VGND VGND VPWR VPWR _3629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9029_ clknet_leaf_59_CLK _0189_ VGND VGND VPWR VPWR RF.registers\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4991_ RF.registers\[8\]\[22\] RF.registers\[9\]\[22\] RF.registers\[10\]\[22\] RF.registers\[11\]\[22\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6730_ _3266_ VGND VGND VPWR VPWR _3278_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ _3241_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8400_ _4168_ VGND VGND VPWR VPWR _4180_ sky130_fd_sc_hd__buf_4
X_5612_ _1167_ _2081_ VGND VGND VPWR VPWR _2367_ sky130_fd_sc_hd__or2_1
X_9380_ clknet_leaf_95_CLK _0540_ VGND VGND VPWR VPWR RF.registers\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6592_ _3041_ RF.registers\[15\]\[9\] _3195_ VGND VGND VPWR VPWR _3205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5543_ _2297_ _2298_ _1738_ VGND VGND VPWR VPWR _2299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8331_ _4143_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5474_ _1639_ _2229_ VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8262_ _3111_ RF.registers\[13\]\[9\] _4097_ VGND VGND VPWR VPWR _4107_ sky130_fd_sc_hd__mux2_1
X_7213_ _3549_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
X_4425_ _1042_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__buf_4
X_8193_ _4070_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__clkbuf_1
X_7144_ RF.registers\[19\]\[29\] _3448_ _3498_ VGND VGND VPWR VPWR _3513_ sky130_fd_sc_hd__mux2_1
X_4356_ RF.registers\[24\]\[2\] RF.registers\[25\]\[2\] RF.registers\[26\]\[2\] RF.registers\[27\]\[2\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7075_ _3467_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
X_4287_ A2[1] VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__clkbuf_4
X_6026_ _2744_ _2749_ _2764_ VGND VGND VPWR VPWR _2765_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7977_ _3099_ RF.registers\[21\]\[3\] _3952_ VGND VGND VPWR VPWR _3956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6928_ _3383_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6859_ RF.registers\[5\]\[6\] _3105_ _3340_ VGND VGND VPWR VPWR _3347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9578_ clknet_leaf_87_CLK _0738_ VGND VGND VPWR VPWR RF.registers\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8529_ RF.registers\[10\]\[7\] net43 _4244_ VGND VGND VPWR VPWR _4248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload14 clknet_leaf_96_CLK VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinv_1
Xclkload25 clknet_leaf_87_CLK VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload69 clknet_leaf_26_CLK VGND VGND VPWR VPWR clkload69/Y sky130_fd_sc_hd__inv_8
Xclkload58 clknet_leaf_14_CLK VGND VGND VPWR VPWR clkload58/Y sky130_fd_sc_hd__inv_6
Xclkload36 clknet_leaf_74_CLK VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_3_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload47 clknet_leaf_63_CLK VGND VGND VPWR VPWR clkload47/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5190_ RF.registers\[28\]\[28\] RF.registers\[29\]\[28\] RF.registers\[30\]\[28\]
+ RF.registers\[31\]\[28\] _1882_ _1884_ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_10_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7900_ _3914_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8880_ clknet_leaf_56_CLK _0040_ VGND VGND VPWR VPWR RF.registers\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7831_ RF.registers\[9\]\[31\] _3452_ _3843_ VGND VGND VPWR VPWR _3878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4974_ _1717_ _1727_ _1729_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__a21oi_1
X_7762_ _3841_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7693_ RF.registers\[2\]\[30\] _3450_ _3771_ VGND VGND VPWR VPWR _3805_ sky130_fd_sc_hd__mux2_1
X_9501_ clknet_leaf_18_CLK _0661_ VGND VGND VPWR VPWR RF.registers\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6713_ _3269_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9432_ clknet_leaf_39_CLK _0592_ VGND VGND VPWR VPWR RF.registers\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6644_ RF.registers\[8\]\[1\] _3095_ _3231_ VGND VGND VPWR VPWR _3233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload8 clknet_leaf_89_CLK VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9363_ clknet_leaf_30_CLK _0523_ VGND VGND VPWR VPWR RF.registers\[20\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6575_ _3196_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9294_ clknet_leaf_21_CLK _0454_ VGND VGND VPWR VPWR RF.registers\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8314_ RF.registers\[16\]\[1\] _3458_ _4133_ VGND VGND VPWR VPWR _4135_ sky130_fd_sc_hd__mux2_1
X_5526_ RF.registers\[4\]\[7\] RF.registers\[5\]\[7\] RF.registers\[6\]\[7\] RF.registers\[7\]\[7\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2282_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_76_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5457_ _1169_ _2194_ _2212_ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__o21ba_1
X_8245_ _4098_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4408_ _1162_ _1163_ _1035_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5388_ _1638_ VGND VGND VPWR VPWR _2144_ sky130_fd_sc_hd__inv_2
X_8176_ RF.registers\[1\]\[0\] _3454_ _4061_ VGND VGND VPWR VPWR _4062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7127_ RF.registers\[19\]\[22\] _3502_ _3498_ VGND VGND VPWR VPWR _3503_ sky130_fd_sc_hd__mux2_1
X_4339_ RF.registers\[28\]\[3\] RF.registers\[29\]\[3\] RF.registers\[30\]\[3\] RF.registers\[31\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7058_ _3455_ VGND VGND VPWR VPWR _3456_ sky130_fd_sc_hd__buf_6
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6009_ _2668_ _2745_ _2748_ VGND VGND VPWR VPWR _2749_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_120_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4690_ _1239_ _1437_ _1445_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6360_ net23 VGND VGND VPWR VPWR _3060_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5311_ _2065_ _2066_ _1645_ VGND VGND VPWR VPWR _2067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6291_ _3012_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__clkbuf_1
X_8030_ _3983_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5242_ _1839_ _1997_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__nor2_1
X_5173_ _1927_ _1928_ _1745_ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 A1[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_8932_ clknet_leaf_77_CLK _0092_ VGND VGND VPWR VPWR RF.registers\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8863_ clknet_leaf_66_CLK _0023_ VGND VGND VPWR VPWR RF.registers\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_7814_ _3869_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8794_ clknet_leaf_46_CLK _0978_ VGND VGND VPWR VPWR RF.registers\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7745_ _3069_ RF.registers\[30\]\[22\] _3830_ VGND VGND VPWR VPWR _3833_ sky130_fd_sc_hd__mux2_1
X_4957_ _1712_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7676_ _3796_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4888_ RF.registers\[16\]\[0\] RF.registers\[17\]\[0\] RF.registers\[18\]\[0\] RF.registers\[19\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6627_ _3223_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9415_ clknet_leaf_59_CLK _0575_ VGND VGND VPWR VPWR RF.registers\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6558_ RF.registers\[0\]\[26\] _3002_ _3179_ VGND VGND VPWR VPWR _3186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9346_ clknet_leaf_91_CLK _0506_ VGND VGND VPWR VPWR RF.registers\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6489_ RF.registers\[17\]\[27\] _3009_ _3135_ VGND VGND VPWR VPWR _3148_ sky130_fd_sc_hd__mux2_1
X_9277_ clknet_leaf_18_CLK _0437_ VGND VGND VPWR VPWR RF.registers\[23\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5509_ _2263_ _2264_ _1712_ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__mux2_1
X_8228_ RF.registers\[1\]\[25\] _3508_ _4083_ VGND VGND VPWR VPWR _4089_ sky130_fd_sc_hd__mux2_1
X_8159_ _4052_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5860_ _2504_ _2604_ _2606_ VGND VGND VPWR VPWR _2607_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4811_ _1071_ _1566_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5791_ _2323_ _2515_ VGND VGND VPWR VPWR _2541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7530_ _3058_ RF.registers\[27\]\[17\] _3711_ VGND VGND VPWR VPWR _3719_ sky130_fd_sc_hd__mux2_1
X_4742_ _1496_ _1497_ _1259_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4673_ _1254_ _1428_ _1170_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7461_ _3682_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9200_ clknet_leaf_6_CLK _0360_ VGND VGND VPWR VPWR RF.registers\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6412_ _3096_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7392_ _3056_ RF.registers\[26\]\[16\] _3639_ VGND VGND VPWR VPWR _3646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9131_ clknet_leaf_0_CLK _0291_ VGND VGND VPWR VPWR RF.registers\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6343_ _3048_ RF.registers\[22\]\[12\] _3044_ VGND VGND VPWR VPWR _3049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6274_ _2254_ _2925_ _2998_ _2337_ VGND VGND VPWR VPWR _2999_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9062_ clknet_leaf_63_CLK _0222_ VGND VGND VPWR VPWR RF.registers\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_102_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5225_ RF.registers\[20\]\[26\] RF.registers\[21\]\[26\] RF.registers\[22\]\[26\]
+ RF.registers\[23\]\[26\] _1881_ _1883_ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__mux4_1
X_8013_ _3134_ RF.registers\[21\]\[20\] _3974_ VGND VGND VPWR VPWR _3975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5156_ _1908_ _1911_ _1700_ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5087_ RF.registers\[20\]\[17\] RF.registers\[21\]\[17\] RF.registers\[22\]\[17\]
+ RF.registers\[23\]\[17\] _1689_ _1693_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__mux4_1
X_8915_ clknet_leaf_27_CLK _0075_ VGND VGND VPWR VPWR RF.registers\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8846_ clknet_leaf_56_CLK _0006_ VGND VGND VPWR VPWR RF.registers\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_111_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5989_ _2716_ _2722_ _2729_ _2621_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__o22a_1
X_8777_ clknet_leaf_82_CLK _0961_ VGND VGND VPWR VPWR RF.registers\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7728_ _3052_ RF.registers\[30\]\[14\] _3819_ VGND VGND VPWR VPWR _3824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7659_ _3787_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_115_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9329_ clknet_leaf_19_CLK _0489_ VGND VGND VPWR VPWR RF.registers\[21\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _1700_ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6961_ RF.registers\[4\]\[22\] _3139_ _3398_ VGND VGND VPWR VPWR _3401_ sky130_fd_sc_hd__mux2_1
X_8700_ clknet_leaf_17_CLK _0884_ VGND VGND VPWR VPWR RF.registers\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6892_ _3364_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__clkbuf_1
X_5912_ _2504_ _2647_ _2653_ _2656_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__o2bb2a_1
X_8631_ clknet_leaf_32_CLK _0815_ VGND VGND VPWR VPWR RF.registers\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5843_ _2039_ _2102_ VGND VGND VPWR VPWR _2591_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_66_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8562_ RF.registers\[10\]\[23\] net29 _4255_ VGND VGND VPWR VPWR _4265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5774_ _2369_ _2360_ VGND VGND VPWR VPWR _2525_ sky130_fd_sc_hd__nand2_1
X_7513_ _3041_ RF.registers\[27\]\[9\] _3700_ VGND VGND VPWR VPWR _3710_ sky130_fd_sc_hd__mux2_1
X_8493_ _4229_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4725_ RF.registers\[24\]\[14\] RF.registers\[25\]\[14\] RF.registers\[26\]\[14\]
+ RF.registers\[27\]\[14\] _1324_ _1325_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7444_ _3673_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__clkbuf_1
X_4656_ RF.registers\[0\]\[7\] RF.registers\[1\]\[7\] RF.registers\[2\]\[7\] RF.registers\[3\]\[7\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4587_ _1211_ _1342_ _1078_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7375_ _3039_ RF.registers\[26\]\[8\] _3628_ VGND VGND VPWR VPWR _3637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9114_ clknet_leaf_25_CLK _0274_ VGND VGND VPWR VPWR RF.registers\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6326_ net43 VGND VGND VPWR VPWR _3037_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9045_ clknet_leaf_25_CLK _0205_ VGND VGND VPWR VPWR RF.registers\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6257_ _1348_ _2982_ VGND VGND VPWR VPWR _2983_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5208_ RF.registers\[16\]\[27\] RF.registers\[17\]\[27\] RF.registers\[18\]\[27\]
+ RF.registers\[19\]\[27\] _1767_ _1768_ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__mux4_1
X_6188_ _1978_ _2915_ VGND VGND VPWR VPWR _2917_ sky130_fd_sc_hd__nand2_1
X_5139_ _1689_ VGND VGND VPWR VPWR _1895_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8829_ clknet_leaf_14_CLK _1013_ VGND VGND VPWR VPWR RF.registers\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ _1260_ _1265_ _1187_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__mux2_1
X_5490_ _1671_ _2237_ _2245_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4441_ _1190_ _1196_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7160_ RF.registers\[7\]\[4\] _3464_ _3517_ VGND VGND VPWR VPWR _3522_ sky130_fd_sc_hd__mux2_1
X_6111_ _2840_ _2844_ VGND VGND VPWR VPWR _2845_ sky130_fd_sc_hd__xor2_1
X_4372_ _1087_ _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7091_ _3478_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6042_ _2420_ _2738_ _2333_ VGND VGND VPWR VPWR _2780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7993_ _3964_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6944_ RF.registers\[4\]\[14\] _3122_ _3387_ VGND VGND VPWR VPWR _3392_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6875_ _3355_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8614_ clknet_leaf_61_CLK _0798_ VGND VGND VPWR VPWR RF.registers\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5826_ _2105_ _2573_ _2574_ _2373_ VGND VGND VPWR VPWR _2575_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5757_ _2305_ _2508_ VGND VGND VPWR VPWR _2509_ sky130_fd_sc_hd__nor2_1
X_8545_ _4256_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4708_ _1215_ _1455_ _1463_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__o21ai_4
X_8476_ _4220_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5688_ _1926_ _2178_ VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__or2b_1
X_7427_ _3019_ RF.registers\[25\]\[0\] _3664_ VGND VGND VPWR VPWR _3665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4639_ RF.registers\[4\]\[6\] RF.registers\[5\]\[6\] RF.registers\[6\]\[6\] RF.registers\[7\]\[6\]
+ _1072_ _1073_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7358_ _3627_ VGND VGND VPWR VPWR _3628_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_9_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7289_ _3590_ VGND VGND VPWR VPWR _3591_ sky130_fd_sc_hd__buf_8
X_6309_ _3025_ RF.registers\[22\]\[1\] _3023_ VGND VGND VPWR VPWR _3026_ sky130_fd_sc_hd__mux2_1
X_9028_ clknet_leaf_96_CLK _0188_ VGND VGND VPWR VPWR RF.registers\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4990_ RF.registers\[12\]\[22\] RF.registers\[13\]\[22\] RF.registers\[14\]\[22\]
+ RF.registers\[15\]\[22\] _1720_ _1723_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6660_ RF.registers\[8\]\[9\] _3111_ _3231_ VGND VGND VPWR VPWR _3241_ sky130_fd_sc_hd__mux2_1
X_5611_ _2365_ VGND VGND VPWR VPWR _2366_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6591_ _3204_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5542_ RF.registers\[8\]\[4\] RF.registers\[9\]\[4\] RF.registers\[10\]\[4\] RF.registers\[11\]\[4\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2298_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8330_ RF.registers\[16\]\[9\] _3474_ _4133_ VGND VGND VPWR VPWR _4143_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_91_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_91_CLK sky130_fd_sc_hd__clkbuf_8
X_5473_ _1671_ _2220_ _2224_ _2228_ VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_14_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8261_ _4106_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__clkbuf_1
X_4424_ RF.registers\[28\]\[29\] RF.registers\[29\]\[29\] RF.registers\[30\]\[29\]
+ RF.registers\[31\]\[29\] _1173_ _1175_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7212_ RF.registers\[7\]\[29\] _3448_ _3539_ VGND VGND VPWR VPWR _3549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8192_ RF.registers\[1\]\[8\] _3472_ _4061_ VGND VGND VPWR VPWR _4070_ sky130_fd_sc_hd__mux2_1
X_7143_ _3512_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_4355_ _1110_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__clkbuf_4
X_7074_ RF.registers\[19\]\[5\] _3466_ _3456_ VGND VGND VPWR VPWR _3467_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_3_0__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_4286_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__clkbuf_8
X_6025_ _1874_ _2743_ VGND VGND VPWR VPWR _2764_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7976_ _3955_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6927_ RF.registers\[4\]\[6\] _3105_ _3376_ VGND VGND VPWR VPWR _3383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6858_ _3346_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5809_ _1415_ _2557_ VGND VGND VPWR VPWR _2558_ sky130_fd_sc_hd__xor2_1
X_9577_ clknet_leaf_88_CLK _0737_ VGND VGND VPWR VPWR RF.registers\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6789_ RF.registers\[6\]\[5\] _3103_ _3304_ VGND VGND VPWR VPWR _3310_ sky130_fd_sc_hd__mux2_1
X_8528_ _4247_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_82_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_82_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8459_ _4211_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload15 clknet_leaf_97_CLK VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__inv_6
Xclkbuf_leaf_73_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_73_CLK sky130_fd_sc_hd__clkbuf_8
Xclkload26 clknet_leaf_98_CLK VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinv_4
Xclkload59 clknet_leaf_15_CLK VGND VGND VPWR VPWR clkload59/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload37 clknet_leaf_75_CLK VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload48 clknet_leaf_80_CLK VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__inv_8
XFILLER_0_121_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7830_ _3877_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7761_ _3085_ RF.registers\[30\]\[30\] _3807_ VGND VGND VPWR VPWR _3841_ sky130_fd_sc_hd__mux2_1
X_4973_ _1728_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_19_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7692_ _3804_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__clkbuf_1
X_9500_ clknet_leaf_17_CLK _0660_ VGND VGND VPWR VPWR RF.registers\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6712_ _3025_ RF.registers\[14\]\[1\] _3267_ VGND VGND VPWR VPWR _3269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9431_ clknet_leaf_49_CLK _0591_ VGND VGND VPWR VPWR RF.registers\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6643_ _3232_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_90_CLK VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__bufinv_16
X_9362_ clknet_leaf_41_CLK _0522_ VGND VGND VPWR VPWR RF.registers\[20\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6574_ _3019_ RF.registers\[15\]\[0\] _3195_ VGND VGND VPWR VPWR _3196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_64_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_64_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9293_ clknet_leaf_4_CLK _0453_ VGND VGND VPWR VPWR RF.registers\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8313_ _4134_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__clkbuf_1
X_5525_ _1699_ _2280_ VGND VGND VPWR VPWR _2281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5456_ _1168_ _2211_ VGND VGND VPWR VPWR _2212_ sky130_fd_sc_hd__and2_1
X_8244_ _3089_ RF.registers\[13\]\[0\] _4097_ VGND VGND VPWR VPWR _4098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4407_ RF.registers\[0\]\[0\] RF.registers\[1\]\[0\] RF.registers\[2\]\[0\] RF.registers\[3\]\[0\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5387_ _1169_ _2124_ _2142_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8175_ _4060_ VGND VGND VPWR VPWR _4061_ sky130_fd_sc_hd__clkbuf_8
X_7126_ net28 VGND VGND VPWR VPWR _3502_ sky130_fd_sc_hd__clkbuf_4
X_4338_ _1088_ _1093_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__nand2_1
X_7057_ _3090_ _3411_ VGND VGND VPWR VPWR _3455_ sky130_fd_sc_hd__nor2_2
X_4269_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__clkbuf_8
X_6008_ _2123_ _2724_ _2746_ _2747_ VGND VGND VPWR VPWR _2748_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ RF.registers\[18\]\[27\] _3444_ _3938_ VGND VGND VPWR VPWR _3946_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_55_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_55_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_46_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_46_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6290_ RF.registers\[10\]\[28\] _3011_ _3007_ VGND VGND VPWR VPWR _3012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5310_ RF.registers\[16\]\[2\] RF.registers\[17\]\[2\] RF.registers\[18\]\[2\] RF.registers\[19\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2066_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5241_ _1842_ _1996_ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5172_ RF.registers\[16\]\[29\] RF.registers\[17\]\[29\] RF.registers\[18\]\[29\]
+ RF.registers\[19\]\[29\] _1705_ _1708_ VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 A1[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
X_8931_ clknet_leaf_75_CLK _0091_ VGND VGND VPWR VPWR RF.registers\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_8862_ clknet_leaf_67_CLK _0022_ VGND VGND VPWR VPWR RF.registers\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8793_ clknet_leaf_50_CLK _0977_ VGND VGND VPWR VPWR RF.registers\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_7813_ RF.registers\[9\]\[22\] _3502_ _3866_ VGND VGND VPWR VPWR _3869_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7744_ _3832_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4956_ _1711_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7675_ RF.registers\[2\]\[21\] _3500_ _3794_ VGND VGND VPWR VPWR _3796_ sky130_fd_sc_hd__mux2_1
X_4887_ RF.registers\[20\]\[0\] RF.registers\[21\]\[0\] RF.registers\[22\]\[0\] RF.registers\[23\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__mux4_1
X_6626_ _3075_ RF.registers\[15\]\[25\] _3217_ VGND VGND VPWR VPWR _3223_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_37_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_37_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9414_ clknet_leaf_61_CLK _0574_ VGND VGND VPWR VPWR RF.registers\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6557_ _3185_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9345_ clknet_leaf_93_CLK _0505_ VGND VGND VPWR VPWR RF.registers\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5508_ RF.registers\[12\]\[6\] RF.registers\[13\]\[6\] RF.registers\[14\]\[6\] RF.registers\[15\]\[6\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__mux4_1
X_6488_ _3147_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__clkbuf_1
X_9276_ clknet_leaf_18_CLK _0436_ VGND VGND VPWR VPWR RF.registers\[23\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_8227_ _4088_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__clkbuf_1
X_5439_ RF.registers\[24\]\[10\] RF.registers\[25\]\[10\] RF.registers\[26\]\[10\]
+ RF.registers\[27\]\[10\] _1674_ _1691_ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__mux4_1
X_8158_ RF.registers\[24\]\[24\] _3506_ _4047_ VGND VGND VPWR VPWR _4052_ sky130_fd_sc_hd__mux2_1
X_7109_ _3490_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_8089_ _4015_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_89_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_28_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4810_ _1564_ _1565_ _1048_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5790_ _2271_ _2538_ VGND VGND VPWR VPWR _2540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4741_ RF.registers\[16\]\[15\] RF.registers\[17\]\[15\] RF.registers\[18\]\[15\]
+ RF.registers\[19\]\[15\] _1262_ _1263_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4672_ _1426_ _1427_ _1211_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_19_CLK sky130_fd_sc_hd__clkbuf_8
X_7460_ _3056_ RF.registers\[25\]\[16\] _3675_ VGND VGND VPWR VPWR _3682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6411_ RF.registers\[17\]\[1\] _3095_ _3093_ VGND VGND VPWR VPWR _3096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7391_ _3645_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9130_ clknet_leaf_8_CLK _0290_ VGND VGND VPWR VPWR RF.registers\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6342_ net17 VGND VGND VPWR VPWR _3048_ sky130_fd_sc_hd__clkbuf_2
X_6273_ _2958_ _2997_ _2363_ VGND VGND VPWR VPWR _2998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9061_ clknet_leaf_59_CLK _0221_ VGND VGND VPWR VPWR RF.registers\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8012_ _3951_ VGND VGND VPWR VPWR _3974_ sky130_fd_sc_hd__buf_4
X_5224_ _1800_ _1979_ VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__nor2_1
X_5155_ _1909_ _1910_ _1745_ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5086_ _1638_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__clkbuf_4
X_8914_ clknet_leaf_42_CLK _0074_ VGND VGND VPWR VPWR RF.registers\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8845_ clknet_leaf_57_CLK _0005_ VGND VGND VPWR VPWR RF.registers\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5988_ _2725_ _2728_ VGND VGND VPWR VPWR _2729_ sky130_fd_sc_hd__xnor2_1
X_8776_ clknet_leaf_78_CLK _0960_ VGND VGND VPWR VPWR RF.registers\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4939_ _1688_ _1694_ _1686_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7727_ _3823_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__clkbuf_1
X_7658_ RF.registers\[2\]\[13\] _3483_ _3783_ VGND VGND VPWR VPWR _3787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6609_ _3058_ RF.registers\[15\]\[17\] _3206_ VGND VGND VPWR VPWR _3214_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7589_ _3750_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9328_ clknet_leaf_15_CLK _0488_ VGND VGND VPWR VPWR RF.registers\[21\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_9259_ clknet_leaf_2_CLK _0419_ VGND VGND VPWR VPWR RF.registers\[23\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_8_CLK sky130_fd_sc_hd__clkbuf_8
X_6960_ _3400_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5911_ _2654_ _2655_ VGND VGND VPWR VPWR _2656_ sky130_fd_sc_hd__or2_1
X_6891_ RF.registers\[5\]\[21\] _3137_ _3362_ VGND VGND VPWR VPWR _3364_ sky130_fd_sc_hd__mux2_1
X_8630_ clknet_leaf_47_CLK _0814_ VGND VGND VPWR VPWR RF.registers\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5842_ _1666_ _2040_ VGND VGND VPWR VPWR _2590_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_66_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8561_ _4264_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5773_ _2338_ _2365_ VGND VGND VPWR VPWR _2524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4724_ _1215_ _1471_ _1475_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__a2bb2o_1
X_7512_ _3709_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8492_ RF.registers\[11\]\[21\] net27 _4227_ VGND VGND VPWR VPWR _4229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7443_ _3039_ RF.registers\[25\]\[8\] _3664_ VGND VGND VPWR VPWR _3673_ sky130_fd_sc_hd__mux2_1
X_4655_ RF.registers\[4\]\[7\] RF.registers\[5\]\[7\] RF.registers\[6\]\[7\] RF.registers\[7\]\[7\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4586_ RF.registers\[8\]\[30\] RF.registers\[9\]\[30\] RF.registers\[10\]\[30\] RF.registers\[11\]\[30\]
+ _1182_ _1184_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__mux4_1
X_7374_ _3636_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
X_9113_ clknet_leaf_27_CLK _0273_ VGND VGND VPWR VPWR RF.registers\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6325_ _3036_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__clkbuf_1
X_9044_ clknet_leaf_23_CLK _0204_ VGND VGND VPWR VPWR RF.registers\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6256_ _2741_ _2981_ VGND VGND VPWR VPWR _2982_ sky130_fd_sc_hd__nor2_1
X_5207_ RF.registers\[20\]\[27\] RF.registers\[21\]\[27\] RF.registers\[22\]\[27\]
+ RF.registers\[23\]\[27\] _1767_ _1768_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__mux4_1
X_6187_ _1978_ _2915_ VGND VGND VPWR VPWR _2916_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5138_ _1773_ _1893_ VGND VGND VPWR VPWR _1894_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5069_ RF.registers\[28\]\[19\] RF.registers\[29\]\[19\] RF.registers\[30\]\[19\]
+ RF.registers\[31\]\[19\] _1676_ _1681_ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8828_ clknet_leaf_16_CLK _1012_ VGND VGND VPWR VPWR RF.registers\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8759_ clknet_leaf_47_CLK _0943_ VGND VGND VPWR VPWR RF.registers\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_130_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4440_ RF.registers\[12\]\[29\] RF.registers\[13\]\[29\] RF.registers\[14\]\[29\]
+ RF.registers\[15\]\[29\] _1192_ _1195_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_414 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4371_ _1111_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__and2_2
X_6110_ _2827_ _2831_ _2843_ VGND VGND VPWR VPWR _2844_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7090_ RF.registers\[19\]\[10\] _3476_ _3477_ VGND VGND VPWR VPWR _3478_ sky130_fd_sc_hd__mux2_1
X_6041_ _2704_ _2778_ _1879_ VGND VGND VPWR VPWR _2779_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7992_ _3113_ RF.registers\[21\]\[10\] _3963_ VGND VGND VPWR VPWR _3964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6943_ _3391_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6874_ RF.registers\[5\]\[13\] _3120_ _3351_ VGND VGND VPWR VPWR _3355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5825_ _2255_ _2461_ _2463_ _2337_ VGND VGND VPWR VPWR _2574_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8613_ clknet_leaf_63_CLK _0797_ VGND VGND VPWR VPWR RF.registers\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5756_ _1060_ _2507_ VGND VGND VPWR VPWR _2508_ sky130_fd_sc_hd__xnor2_1
X_8544_ RF.registers\[10\]\[14\] net19 _4255_ VGND VGND VPWR VPWR _4256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5687_ _2252_ _2437_ _2440_ VGND VGND VPWR VPWR _2441_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8475_ RF.registers\[11\]\[13\] net18 _4216_ VGND VGND VPWR VPWR _4220_ sky130_fd_sc_hd__mux2_1
X_4707_ _1457_ _1459_ _1462_ _1071_ _1057_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7426_ _3663_ VGND VGND VPWR VPWR _3664_ sky130_fd_sc_hd__buf_6
X_4638_ _1036_ _1393_ _1037_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7357_ _3020_ _3626_ VGND VGND VPWR VPWR _3627_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_9_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4569_ _1029_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_92_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7288_ _3193_ _3553_ VGND VGND VPWR VPWR _3590_ sky130_fd_sc_hd__nand2_4
X_6308_ net25 VGND VGND VPWR VPWR _3025_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6239_ _2965_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
X_9027_ clknet_leaf_75_CLK _0187_ VGND VGND VPWR VPWR RF.registers\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5610_ _1169_ _2098_ _1803_ VGND VGND VPWR VPWR _2365_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6590_ _3039_ RF.registers\[15\]\[8\] _3195_ VGND VGND VPWR VPWR _3204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5541_ RF.registers\[12\]\[4\] RF.registers\[13\]\[4\] RF.registers\[14\]\[4\] RF.registers\[15\]\[4\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8260_ _3109_ RF.registers\[13\]\[8\] _4097_ VGND VGND VPWR VPWR _4106_ sky130_fd_sc_hd__mux2_1
X_7211_ _3548_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5472_ _1717_ _2227_ _1729_ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4423_ _1176_ _1177_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__mux2_1
X_8191_ _4069_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__clkbuf_1
X_7142_ RF.registers\[19\]\[28\] _3446_ _3498_ VGND VGND VPWR VPWR _3512_ sky130_fd_sc_hd__mux2_1
X_4354_ _1057_ _1094_ _1098_ _1102_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a32o_2
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7073_ net41 VGND VGND VPWR VPWR _3466_ sky130_fd_sc_hd__buf_2
X_6024_ _1858_ _2762_ VGND VGND VPWR VPWR _2763_ sky130_fd_sc_hd__xor2_1
X_4285_ A2[0] VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7975_ _3097_ RF.registers\[21\]\[2\] _3952_ VGND VGND VPWR VPWR _3955_ sky130_fd_sc_hd__mux2_1
X_6926_ _3382_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6857_ RF.registers\[5\]\[5\] _3103_ _3340_ VGND VGND VPWR VPWR _3346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5808_ _1399_ _2506_ _2535_ _2411_ VGND VGND VPWR VPWR _2557_ sky130_fd_sc_hd__a31o_1
X_6788_ _3309_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__clkbuf_1
X_9576_ clknet_leaf_88_CLK _0736_ VGND VGND VPWR VPWR RF.registers\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5739_ _2490_ _2179_ _2426_ VGND VGND VPWR VPWR _2491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8527_ RF.registers\[10\]\[6\] net42 _4244_ VGND VGND VPWR VPWR _4247_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8458_ RF.registers\[11\]\[5\] net41 _4205_ VGND VGND VPWR VPWR _4211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7409_ _3073_ RF.registers\[26\]\[24\] _3650_ VGND VGND VPWR VPWR _3655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8389_ _4174_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload16 clknet_leaf_2_CLK VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload38 clknet_leaf_76_CLK VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__clkinv_1
Xclkload27 clknet_leaf_64_CLK VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__bufinv_16
Xclkload49 clknet_leaf_81_CLK VGND VGND VPWR VPWR clkload49/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7760_ _3840_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4972_ net5 VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7691_ RF.registers\[2\]\[29\] _3448_ _3794_ VGND VGND VPWR VPWR _3804_ sky130_fd_sc_hd__mux2_1
X_6711_ _3268_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__clkbuf_1
X_9430_ clknet_leaf_48_CLK _0590_ VGND VGND VPWR VPWR RF.registers\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6642_ RF.registers\[8\]\[0\] _3089_ _3231_ VGND VGND VPWR VPWR _3232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9361_ clknet_leaf_18_CLK _0521_ VGND VGND VPWR VPWR RF.registers\[20\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8312_ RF.registers\[16\]\[0\] _3454_ _4133_ VGND VGND VPWR VPWR _4134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6573_ _3194_ VGND VGND VPWR VPWR _3195_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5524_ _2278_ _2279_ _1685_ VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__mux2_1
X_9292_ clknet_leaf_3_CLK _0452_ VGND VGND VPWR VPWR RF.registers\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5455_ _1639_ _2210_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__or2_1
X_8243_ _4096_ VGND VGND VPWR VPWR _4097_ sky130_fd_sc_hd__clkbuf_8
X_8174_ _3091_ _3153_ VGND VGND VPWR VPWR _4060_ sky130_fd_sc_hd__nor2_4
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4406_ RF.registers\[4\]\[0\] RF.registers\[5\]\[0\] RF.registers\[6\]\[0\] RF.registers\[7\]\[0\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__mux4_1
X_7125_ _3501_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5386_ _1669_ _2141_ VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__nor2_1
X_4337_ _1091_ _1092_ _1040_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7056_ net14 VGND VGND VPWR VPWR _3454_ sky130_fd_sc_hd__buf_2
X_4268_ net8 VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__inv_2
X_6007_ _2123_ _2724_ _2726_ VGND VGND VPWR VPWR _2747_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_120_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7958_ _3945_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7889_ _3002_ RF.registers\[23\]\[26\] _3902_ VGND VGND VPWR VPWR _3909_ sky130_fd_sc_hd__mux2_1
X_6909_ RF.registers\[5\]\[30\] _3015_ _3339_ VGND VGND VPWR VPWR _3373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9559_ clknet_leaf_47_CLK _0719_ VGND VGND VPWR VPWR RF.registers\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5240_ _1777_ _1987_ _1995_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_58_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5171_ RF.registers\[20\]\[29\] RF.registers\[21\]\[29\] RF.registers\[22\]\[29\]
+ RF.registers\[23\]\[29\] _1705_ _1708_ VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8930_ clknet_leaf_91_CLK _0090_ VGND VGND VPWR VPWR RF.registers\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xinput3 A1[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
X_8861_ clknet_leaf_14_CLK _0021_ VGND VGND VPWR VPWR RF.registers\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_7812_ _3868_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__clkbuf_1
X_8792_ clknet_leaf_40_CLK _0976_ VGND VGND VPWR VPWR RF.registers\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7743_ _3067_ RF.registers\[30\]\[21\] _3830_ VGND VGND VPWR VPWR _3832_ sky130_fd_sc_hd__mux2_1
X_4955_ net3 VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7674_ _3795_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4886_ net2 VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__clkbuf_4
X_6625_ _3222_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9413_ clknet_leaf_81_CLK _0573_ VGND VGND VPWR VPWR RF.registers\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6556_ RF.registers\[0\]\[25\] _3145_ _3179_ VGND VGND VPWR VPWR _3185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9344_ clknet_leaf_70_CLK _0504_ VGND VGND VPWR VPWR RF.registers\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9275_ clknet_leaf_46_CLK _0435_ VGND VGND VPWR VPWR RF.registers\[23\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5507_ RF.registers\[8\]\[6\] RF.registers\[9\]\[6\] RF.registers\[10\]\[6\] RF.registers\[11\]\[6\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2263_ sky130_fd_sc_hd__mux4_1
X_8226_ RF.registers\[1\]\[24\] _3506_ _4083_ VGND VGND VPWR VPWR _4088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6487_ RF.registers\[17\]\[26\] _3002_ _3135_ VGND VGND VPWR VPWR _3147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5438_ _2144_ _2193_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8157_ _4051_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5369_ RF.registers\[20\]\[14\] RF.registers\[21\]\[14\] RF.registers\[22\]\[14\]
+ RF.registers\[23\]\[14\] _1733_ _1679_ VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__mux4_1
X_8088_ RF.registers\[20\]\[23\] _3504_ _4011_ VGND VGND VPWR VPWR _4015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7108_ RF.registers\[19\]\[16\] _3489_ _3477_ VGND VGND VPWR VPWR _3490_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7039_ RF.registers\[3\]\[26\] _3442_ _3435_ VGND VGND VPWR VPWR _3443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4740_ RF.registers\[20\]\[15\] RF.registers\[21\]\[15\] RF.registers\[22\]\[15\]
+ RF.registers\[23\]\[15\] _1262_ _1263_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4671_ RF.registers\[0\]\[23\] RF.registers\[1\]\[23\] RF.registers\[2\]\[23\] RF.registers\[3\]\[23\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7390_ _3054_ RF.registers\[26\]\[15\] _3639_ VGND VGND VPWR VPWR _3645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6410_ net25 VGND VGND VPWR VPWR _3095_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6341_ _3047_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6272_ _2379_ _2377_ VGND VGND VPWR VPWR _2997_ sky130_fd_sc_hd__or2_1
X_9060_ clknet_leaf_96_CLK _0220_ VGND VGND VPWR VPWR RF.registers\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_5223_ _1842_ _1978_ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__nor2_1
X_8011_ _3973_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5154_ RF.registers\[24\]\[30\] RF.registers\[25\]\[30\] RF.registers\[26\]\[30\]
+ RF.registers\[27\]\[30\] _1895_ _1897_ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__mux4_1
XFILLER_0_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5085_ _1669_ _1821_ _1840_ VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_16_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8913_ clknet_leaf_19_CLK _0073_ VGND VGND VPWR VPWR RF.registers\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8844_ clknet_leaf_83_CLK _0004_ VGND VGND VPWR VPWR RF.registers\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5987_ _2726_ _2727_ VGND VGND VPWR VPWR _2728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8775_ clknet_leaf_60_CLK _0959_ VGND VGND VPWR VPWR RF.registers\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_4938_ RF.registers\[24\]\[23\] RF.registers\[25\]\[23\] RF.registers\[26\]\[23\]
+ RF.registers\[27\]\[23\] _1689_ _1693_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__mux4_1
X_7726_ _3050_ RF.registers\[30\]\[13\] _3819_ VGND VGND VPWR VPWR _3823_ sky130_fd_sc_hd__mux2_1
X_4869_ _1621_ _1624_ _1213_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_25_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7657_ _3786_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6608_ _3213_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7588_ _3048_ RF.registers\[28\]\[12\] _3747_ VGND VGND VPWR VPWR _3750_ sky130_fd_sc_hd__mux2_1
X_6539_ RF.registers\[0\]\[17\] _3128_ _3168_ VGND VGND VPWR VPWR _3176_ sky130_fd_sc_hd__mux2_1
X_9327_ clknet_leaf_5_CLK _0487_ VGND VGND VPWR VPWR RF.registers\[21\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9258_ clknet_leaf_9_CLK _0418_ VGND VGND VPWR VPWR RF.registers\[23\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8209_ RF.registers\[1\]\[16\] _3489_ _4072_ VGND VGND VPWR VPWR _4079_ sky130_fd_sc_hd__mux2_1
X_9189_ clknet_leaf_80_CLK _0349_ VGND VGND VPWR VPWR RF.registers\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_43_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5910_ _2471_ _2605_ _2591_ _2462_ VGND VGND VPWR VPWR _2655_ sky130_fd_sc_hd__a22o_1
X_6890_ _3363_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5841_ _1880_ _2588_ _2421_ VGND VGND VPWR VPWR _2589_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8560_ RF.registers\[10\]\[22\] net28 _4255_ VGND VGND VPWR VPWR _4264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5772_ _1111_ _2522_ _2487_ _2382_ VGND VGND VPWR VPWR _2523_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8491_ _4228_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__clkbuf_1
X_4723_ _1205_ _1478_ _1170_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7511_ _3039_ RF.registers\[27\]\[8\] _3700_ VGND VGND VPWR VPWR _3709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7442_ _3672_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4654_ _1071_ _1409_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4585_ _1189_ _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7373_ _3037_ RF.registers\[26\]\[7\] _3628_ VGND VGND VPWR VPWR _3636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9112_ clknet_leaf_38_CLK _0272_ VGND VGND VPWR VPWR RF.registers\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6324_ _3035_ RF.registers\[22\]\[6\] _3023_ VGND VGND VPWR VPWR _3036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9043_ clknet_leaf_25_CLK _0203_ VGND VGND VPWR VPWR RF.registers\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6255_ _1238_ _2929_ VGND VGND VPWR VPWR _2981_ sky130_fd_sc_hd__nor2_1
X_5206_ _1926_ _1961_ _1877_ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__mux2_2
X_6186_ _1315_ _2914_ VGND VGND VPWR VPWR _2915_ sky130_fd_sc_hd__xor2_1
X_5137_ _1891_ _1892_ _1889_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5068_ RF.registers\[24\]\[19\] RF.registers\[25\]\[19\] RF.registers\[26\]\[19\]
+ RF.registers\[27\]\[19\] _1822_ _1823_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__mux4_1
X_8827_ clknet_leaf_44_CLK _1011_ VGND VGND VPWR VPWR RF.registers\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8758_ clknet_leaf_33_CLK _0942_ VGND VGND VPWR VPWR RF.registers\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7709_ _3033_ RF.registers\[30\]\[5\] _3808_ VGND VGND VPWR VPWR _3814_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8689_ clknet_leaf_12_CLK _0873_ VGND VGND VPWR VPWR RF.registers\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4370_ _1125_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6040_ _2734_ _2777_ _1877_ VGND VGND VPWR VPWR _2778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7991_ _3951_ VGND VGND VPWR VPWR _3963_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6942_ RF.registers\[4\]\[13\] _3120_ _3387_ VGND VGND VPWR VPWR _3391_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6873_ _3354_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__clkbuf_1
X_5824_ _2470_ _2460_ _2252_ VGND VGND VPWR VPWR _2573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8612_ clknet_leaf_95_CLK _0796_ VGND VGND VPWR VPWR RF.registers\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5755_ _2411_ _2506_ VGND VGND VPWR VPWR _2507_ sky130_fd_sc_hd__nor2_1
X_8543_ _3006_ VGND VGND VPWR VPWR _4255_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_20_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5686_ _2252_ _2439_ VGND VGND VPWR VPWR _2440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8474_ _4219_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__clkbuf_1
X_4706_ _1460_ _1461_ _1048_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7425_ _3552_ _3626_ VGND VGND VPWR VPWR _3663_ sky130_fd_sc_hd__nand2_4
XFILLER_0_72_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4637_ RF.registers\[12\]\[6\] RF.registers\[13\]\[6\] RF.registers\[14\]\[6\] RF.registers\[15\]\[6\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7356_ net11 net12 net13 VGND VGND VPWR VPWR _3626_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_9_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4568_ _1027_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_92_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4499_ _1248_ _1250_ _1253_ _1254_ _1170_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__a221o_1
X_7287_ _3589_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
X_6307_ _3024_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__clkbuf_1
X_6238_ _2957_ _2963_ _2964_ VGND VGND VPWR VPWR _2965_ sky130_fd_sc_hd__or3_1
X_9026_ clknet_leaf_92_CLK _0186_ VGND VGND VPWR VPWR RF.registers\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6169_ _2613_ _2737_ _2898_ _2899_ VGND VGND VPWR VPWR _2900_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5540_ _2292_ _2295_ _1696_ VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5471_ _2225_ _2226_ _1739_ VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7210_ RF.registers\[7\]\[28\] _3446_ _3539_ VGND VGND VPWR VPWR _3548_ sky130_fd_sc_hd__mux2_1
X_4422_ _1036_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8190_ RF.registers\[1\]\[7\] _3470_ _4061_ VGND VGND VPWR VPWR _4069_ sky130_fd_sc_hd__mux2_1
X_7141_ _3511_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
X_4353_ _1088_ _1108_ net8 VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7072_ _3465_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
X_4284_ _1034_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__buf_4
X_6023_ _1601_ _2761_ VGND VGND VPWR VPWR _2762_ sky130_fd_sc_hd__xor2_1
X_7974_ _3954_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6925_ RF.registers\[4\]\[5\] _3103_ _3376_ VGND VGND VPWR VPWR _3382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6856_ _3345_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5807_ _2504_ _2544_ _2545_ _2556_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__a31o_1
X_6787_ RF.registers\[6\]\[4\] _3101_ _3304_ VGND VGND VPWR VPWR _3309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9575_ clknet_leaf_81_CLK _0735_ VGND VGND VPWR VPWR RF.registers\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_5738_ _1878_ VGND VGND VPWR VPWR _2490_ sky130_fd_sc_hd__inv_2
X_8526_ _4246_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5669_ _1876_ VGND VGND VPWR VPWR _2423_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8457_ _4210_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7408_ _3654_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__clkbuf_1
X_8388_ RF.registers\[12\]\[4\] _3464_ _4169_ VGND VGND VPWR VPWR _4174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7339_ _3617_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_8_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9009_ clknet_leaf_19_CLK _0169_ VGND VGND VPWR VPWR RF.registers\[31\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload17 clknet_leaf_3_CLK VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_11_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload39 clknet_leaf_77_CLK VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload28 clknet_leaf_65_CLK VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_50_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _1724_ _1725_ _1726_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7690_ _3803_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__clkbuf_1
X_6710_ _3019_ RF.registers\[14\]\[0\] _3267_ VGND VGND VPWR VPWR _3268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6641_ _3230_ VGND VGND VPWR VPWR _3231_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9360_ clknet_leaf_11_CLK _0520_ VGND VGND VPWR VPWR RF.registers\[20\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6572_ _3192_ _3193_ VGND VGND VPWR VPWR _3194_ sky130_fd_sc_hd__nand2_4
X_8311_ _4132_ VGND VGND VPWR VPWR _4133_ sky130_fd_sc_hd__buf_6
XFILLER_0_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9291_ clknet_leaf_98_CLK _0451_ VGND VGND VPWR VPWR RF.registers\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5523_ RF.registers\[8\]\[7\] RF.registers\[9\]\[7\] RF.registers\[10\]\[7\] RF.registers\[11\]\[7\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_76_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8242_ _3552_ _3192_ VGND VGND VPWR VPWR _4096_ sky130_fd_sc_hd__nand2_2
X_5454_ _1670_ _2201_ _2205_ _2209_ VGND VGND VPWR VPWR _2210_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_42_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8173_ _4059_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__clkbuf_1
X_5385_ _1639_ _2140_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__nor2_1
X_4405_ _1038_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nand2_1
X_7124_ RF.registers\[19\]\[21\] _3500_ _3498_ VGND VGND VPWR VPWR _3501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4336_ RF.registers\[16\]\[3\] RF.registers\[17\]\[3\] RF.registers\[18\]\[3\] RF.registers\[19\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7055_ _3453_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
X_6006_ _2712_ _2713_ _2725_ VGND VGND VPWR VPWR _2746_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_120_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7957_ RF.registers\[18\]\[26\] _3442_ _3938_ VGND VGND VPWR VPWR _3945_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7888_ _3908_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__clkbuf_1
X_6908_ _3372_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6839_ RF.registers\[6\]\[29\] _3013_ _3326_ VGND VGND VPWR VPWR _3336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9558_ clknet_leaf_34_CLK _0718_ VGND VGND VPWR VPWR RF.registers\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8509_ _4237_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__clkbuf_1
X_9489_ clknet_leaf_18_CLK _0649_ VGND VGND VPWR VPWR RF.registers\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5170_ _1169_ _1905_ _1925_ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_71_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 A1[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8860_ clknet_leaf_38_CLK _0020_ VGND VGND VPWR VPWR RF.registers\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8791_ clknet_leaf_49_CLK _0975_ VGND VGND VPWR VPWR RF.registers\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_7811_ RF.registers\[9\]\[21\] _3500_ _3866_ VGND VGND VPWR VPWR _3868_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4954_ RF.registers\[12\]\[23\] RF.registers\[13\]\[23\] RF.registers\[14\]\[23\]
+ RF.registers\[15\]\[23\] _1705_ _1708_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__mux4_1
X_7742_ _3831_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7673_ RF.registers\[2\]\[20\] _3497_ _3794_ VGND VGND VPWR VPWR _3795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4885_ net1 VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__buf_4
X_9412_ clknet_leaf_77_CLK _0572_ VGND VGND VPWR VPWR RF.registers\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6624_ _3073_ RF.registers\[15\]\[24\] _3217_ VGND VGND VPWR VPWR _3222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6555_ _3184_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9343_ clknet_leaf_65_CLK _0503_ VGND VGND VPWR VPWR RF.registers\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9274_ clknet_leaf_37_CLK _0434_ VGND VGND VPWR VPWR RF.registers\[23\]\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_89_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5506_ _2258_ _2261_ _1696_ VGND VGND VPWR VPWR _2262_ sky130_fd_sc_hd__mux2_1
X_6486_ _3146_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__clkbuf_1
X_8225_ _4087_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__clkbuf_1
X_5437_ _1670_ _2184_ _2188_ _2192_ VGND VGND VPWR VPWR _2193_ sky130_fd_sc_hd__o22a_2
X_8156_ RF.registers\[24\]\[23\] _3504_ _4047_ VGND VGND VPWR VPWR _4051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5368_ _1639_ _2123_ VGND VGND VPWR VPWR _2124_ sky130_fd_sc_hd__nor2_1
X_8087_ _4014_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__clkbuf_1
X_7107_ net21 VGND VGND VPWR VPWR _3489_ sky130_fd_sc_hd__clkbuf_4
X_5299_ RF.registers\[12\]\[3\] RF.registers\[13\]\[3\] RF.registers\[14\]\[3\] RF.registers\[15\]\[3\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__mux4_1
X_4319_ RF.registers\[12\]\[5\] RF.registers\[13\]\[5\] RF.registers\[14\]\[5\] RF.registers\[15\]\[5\]
+ _1072_ _1073_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_89_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7038_ net32 VGND VGND VPWR VPWR _3442_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_98_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8989_ clknet_leaf_22_CLK _0149_ VGND VGND VPWR VPWR RF.registers\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4670_ RF.registers\[4\]\[23\] RF.registers\[5\]\[23\] RF.registers\[6\]\[23\] RF.registers\[7\]\[23\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6340_ _3046_ RF.registers\[22\]\[11\] _3044_ VGND VGND VPWR VPWR _3047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6271_ _2942_ VGND VGND VPWR VPWR _2996_ sky130_fd_sc_hd__inv_2
X_5222_ _1777_ _1969_ _1973_ _1977_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__o2bb2a_2
X_8010_ _3132_ RF.registers\[21\]\[19\] _3963_ VGND VGND VPWR VPWR _3973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5153_ RF.registers\[28\]\[30\] RF.registers\[29\]\[30\] RF.registers\[30\]\[30\]
+ RF.registers\[31\]\[30\] _1895_ _1897_ VGND VGND VPWR VPWR _1909_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5084_ _1758_ _1838_ _1839_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8912_ clknet_leaf_7_CLK _0072_ VGND VGND VPWR VPWR RF.registers\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8843_ clknet_leaf_78_CLK _0003_ VGND VGND VPWR VPWR RF.registers\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_84_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5986_ _2712_ _2714_ VGND VGND VPWR VPWR _2727_ sky130_fd_sc_hd__or2b_1
X_8774_ clknet_leaf_61_CLK _0958_ VGND VGND VPWR VPWR RF.registers\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_4937_ _1692_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__buf_4
X_7725_ _3822_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 _1416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _1622_ _1623_ _1259_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__mux2_1
X_7656_ RF.registers\[2\]\[12\] _3481_ _3783_ VGND VGND VPWR VPWR _3786_ sky130_fd_sc_hd__mux2_1
X_6607_ _3056_ RF.registers\[15\]\[16\] _3206_ VGND VGND VPWR VPWR _3213_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_3_6__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_9326_ clknet_leaf_21_CLK _0486_ VGND VGND VPWR VPWR RF.registers\[21\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4799_ RF.registers\[0\]\[10\] RF.registers\[1\]\[10\] RF.registers\[2\]\[10\] RF.registers\[3\]\[10\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__mux4_1
X_7587_ _3749_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6538_ _3175_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6469_ _3092_ VGND VGND VPWR VPWR _3135_ sky130_fd_sc_hd__buf_4
X_9257_ clknet_leaf_9_CLK _0417_ VGND VGND VPWR VPWR RF.registers\[23\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8208_ _4078_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__clkbuf_1
X_9188_ clknet_leaf_96_CLK _0348_ VGND VGND VPWR VPWR RF.registers\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8139_ RF.registers\[24\]\[15\] _3487_ _4036_ VGND VGND VPWR VPWR _4042_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5840_ _2040_ _2372_ VGND VGND VPWR VPWR _2588_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5771_ _2388_ _2397_ _1126_ VGND VGND VPWR VPWR _2522_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8490_ RF.registers\[11\]\[20\] net26 _4227_ VGND VGND VPWR VPWR _4228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4722_ _1476_ _1477_ _1198_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__mux2_1
X_7510_ _3708_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7441_ _3037_ RF.registers\[25\]\[7\] _3664_ VGND VGND VPWR VPWR _3672_ sky130_fd_sc_hd__mux2_1
Xinput40 WD3[4] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
X_4653_ _1407_ _1408_ _1040_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__mux2_1
X_4584_ RF.registers\[12\]\[30\] RF.registers\[13\]\[30\] RF.registers\[14\]\[30\]
+ RF.registers\[15\]\[30\] _1220_ _1222_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__mux4_1
X_7372_ _3635_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
X_9111_ clknet_leaf_31_CLK _0271_ VGND VGND VPWR VPWR RF.registers\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6323_ net42 VGND VGND VPWR VPWR _3035_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9042_ clknet_leaf_41_CLK _0202_ VGND VGND VPWR VPWR RF.registers\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6254_ _2974_ _2797_ _2979_ _2421_ VGND VGND VPWR VPWR _2980_ sky130_fd_sc_hd__o211a_1
X_5205_ _1944_ _1960_ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6185_ _1447_ _1299_ _2901_ _2871_ _2741_ VGND VGND VPWR VPWR _2914_ sky130_fd_sc_hd__a41o_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5136_ RF.registers\[12\]\[31\] RF.registers\[13\]\[31\] RF.registers\[14\]\[31\]
+ RF.registers\[15\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__mux4_1
X_5067_ _1735_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_4_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8826_ clknet_leaf_42_CLK _1010_ VGND VGND VPWR VPWR RF.registers\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8757_ clknet_leaf_29_CLK _0941_ VGND VGND VPWR VPWR RF.registers\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5969_ _1494_ _2710_ VGND VGND VPWR VPWR _2711_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7708_ _3813_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8688_ clknet_leaf_12_CLK _0872_ VGND VGND VPWR VPWR RF.registers\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_7639_ RF.registers\[2\]\[4\] _3464_ _3772_ VGND VGND VPWR VPWR _3777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9309_ clknet_leaf_18_CLK _0469_ VGND VGND VPWR VPWR RF.registers\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7990_ _3962_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_1
X_6941_ _3390_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6872_ RF.registers\[5\]\[12\] _3118_ _3351_ VGND VGND VPWR VPWR _3354_ sky130_fd_sc_hd__mux2_1
X_9591_ clknet_leaf_47_CLK _0751_ VGND VGND VPWR VPWR RF.registers\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5823_ _2472_ _2570_ _2571_ _1111_ VGND VGND VPWR VPWR _2572_ sky130_fd_sc_hd__a22o_1
X_8611_ clknet_leaf_75_CLK _0795_ VGND VGND VPWR VPWR RF.registers\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8542_ _4254_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__clkbuf_1
X_5754_ _1110_ _1125_ _1144_ _1166_ VGND VGND VPWR VPWR _2506_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_94_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_94_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5685_ _2178_ _1802_ _2438_ VGND VGND VPWR VPWR _2439_ sky130_fd_sc_hd__o21ai_1
X_8473_ RF.registers\[11\]\[12\] net17 _4216_ VGND VGND VPWR VPWR _4219_ sky130_fd_sc_hd__mux2_1
X_4705_ RF.registers\[12\]\[12\] RF.registers\[13\]\[12\] RF.registers\[14\]\[12\]
+ RF.registers\[15\]\[12\] _1181_ _1183_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7424_ _3662_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4636_ _1048_ _1391_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7355_ _3625_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4567_ _1319_ _1322_ _1213_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6306_ _3019_ RF.registers\[22\]\[0\] _3023_ VGND VGND VPWR VPWR _3024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7286_ _3087_ RF.registers\[29\]\[31\] _3554_ VGND VGND VPWR VPWR _3589_ sky130_fd_sc_hd__mux2_1
X_4498_ _1205_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6237_ _2701_ _2797_ VGND VGND VPWR VPWR _2964_ sky130_fd_sc_hd__nor2_1
X_9025_ clknet_leaf_97_CLK _0185_ VGND VGND VPWR VPWR RF.registers\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6168_ _2390_ _2864_ _2333_ VGND VGND VPWR VPWR _2899_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5119_ _1758_ _1874_ _1800_ VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__o21ai_1
X_6099_ _2806_ _2827_ _2831_ _2833_ VGND VGND VPWR VPWR _2834_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_28_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8809_ clknet_leaf_82_CLK _0993_ VGND VGND VPWR VPWR RF.registers\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_85_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_76_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_76_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5470_ RF.registers\[0\]\[8\] RF.registers\[1\]\[8\] RF.registers\[2\]\[8\] RF.registers\[3\]\[8\]
+ _1734_ _1735_ VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__mux4_1
X_4421_ RF.registers\[16\]\[29\] RF.registers\[17\]\[29\] RF.registers\[18\]\[29\]
+ RF.registers\[19\]\[29\] _1173_ _1175_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7140_ RF.registers\[19\]\[27\] _3444_ _3498_ VGND VGND VPWR VPWR _3511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4352_ _1103_ _1106_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__mux2_1
X_4283_ _1030_ _1031_ _1032_ _1033_ _1036_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__mux4_1
X_7071_ RF.registers\[19\]\[4\] _3464_ _3456_ VGND VGND VPWR VPWR _3465_ sky130_fd_sc_hd__mux2_1
X_6022_ _1512_ _1587_ _2658_ _2741_ VGND VGND VPWR VPWR _2761_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7973_ _3095_ RF.registers\[21\]\[1\] _3952_ VGND VGND VPWR VPWR _3954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6924_ _3381_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ RF.registers\[5\]\[4\] _3101_ _3340_ VGND VGND VPWR VPWR _3345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5806_ _2496_ _2549_ _2552_ _2555_ VGND VGND VPWR VPWR _2556_ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9574_ clknet_leaf_60_CLK _0734_ VGND VGND VPWR VPWR RF.registers\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_67_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_67_CLK sky130_fd_sc_hd__clkbuf_8
X_6786_ _3308_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5737_ _1666_ _2488_ VGND VGND VPWR VPWR _2489_ sky130_fd_sc_hd__nor2_1
X_8525_ RF.registers\[10\]\[5\] net41 _4244_ VGND VGND VPWR VPWR _4246_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8456_ RF.registers\[11\]\[4\] net40 _4205_ VGND VGND VPWR VPWR _4210_ sky130_fd_sc_hd__mux2_1
X_7407_ _3071_ RF.registers\[26\]\[23\] _3650_ VGND VGND VPWR VPWR _3654_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5668_ _1128_ _2420_ _2421_ VGND VGND VPWR VPWR _2422_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4619_ _1371_ _1372_ _1373_ _1374_ _1190_ _1254_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5599_ _2352_ _2353_ VGND VGND VPWR VPWR _2354_ sky130_fd_sc_hd__and2_1
X_8387_ _4173_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__clkbuf_1
X_7338_ _3071_ RF.registers\[31\]\[23\] _3613_ VGND VGND VPWR VPWR _3617_ sky130_fd_sc_hd__mux2_1
X_7269_ _3580_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
X_9008_ clknet_leaf_6_CLK _0168_ VGND VGND VPWR VPWR RF.registers\[31\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_58_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_58_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_136_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload18 clknet_leaf_4_CLK VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_11_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload29 clknet_leaf_66_CLK VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_6
XFILLER_0_35_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4970_ _1685_ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_49_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_49_CLK sky130_fd_sc_hd__clkbuf_8
X_6640_ _3003_ _3155_ VGND VGND VPWR VPWR _3230_ sky130_fd_sc_hd__nor2_2
XFILLER_0_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6571_ net10 net9 net46 VGND VGND VPWR VPWR _3193_ sky130_fd_sc_hd__and3_2
XFILLER_0_6_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8310_ _3090_ _3155_ VGND VGND VPWR VPWR _4132_ sky130_fd_sc_hd__nor2_2
XFILLER_0_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5522_ RF.registers\[12\]\[7\] RF.registers\[13\]\[7\] RF.registers\[14\]\[7\] RF.registers\[15\]\[7\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2278_ sky130_fd_sc_hd__mux4_1
X_9290_ clknet_leaf_7_CLK _0450_ VGND VGND VPWR VPWR RF.registers\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8241_ _4095_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5453_ _1828_ _2208_ _1728_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_136_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8172_ RF.registers\[24\]\[31\] _3452_ _4024_ VGND VGND VPWR VPWR _4059_ sky130_fd_sc_hd__mux2_1
X_5384_ _1670_ _2131_ _2135_ _2139_ VGND VGND VPWR VPWR _2140_ sky130_fd_sc_hd__a2bb2o_2
X_4404_ _1158_ _1159_ _1047_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__mux2_1
X_7123_ net27 VGND VGND VPWR VPWR _3500_ sky130_fd_sc_hd__clkbuf_4
X_4335_ RF.registers\[20\]\[3\] RF.registers\[21\]\[3\] RF.registers\[22\]\[3\] RF.registers\[23\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__mux4_1
X_7054_ RF.registers\[3\]\[31\] _3452_ _3412_ VGND VGND VPWR VPWR _3453_ sky130_fd_sc_hd__mux2_1
X_6005_ _2663_ _2689_ _2712_ _2725_ VGND VGND VPWR VPWR _2745_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7956_ _3944_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_120_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7887_ _3145_ RF.registers\[23\]\[25\] _3902_ VGND VGND VPWR VPWR _3908_ sky130_fd_sc_hd__mux2_1
X_6907_ RF.registers\[5\]\[29\] _3013_ _3362_ VGND VGND VPWR VPWR _3372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6838_ _3335_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9557_ clknet_leaf_35_CLK _0717_ VGND VGND VPWR VPWR RF.registers\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8508_ RF.registers\[11\]\[29\] net35 _4227_ VGND VGND VPWR VPWR _4237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6769_ _3298_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9488_ clknet_leaf_10_CLK _0648_ VGND VGND VPWR VPWR RF.registers\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8439_ _4200_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 A1[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_0_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7810_ _3867_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__clkbuf_1
X_8790_ clknet_leaf_47_CLK _0974_ VGND VGND VPWR VPWR RF.registers\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_4953_ RF.registers\[8\]\[23\] RF.registers\[9\]\[23\] RF.registers\[10\]\[23\] RF.registers\[11\]\[23\]
+ _1705_ _1708_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__mux4_1
X_7741_ _3064_ RF.registers\[30\]\[20\] _3830_ VGND VGND VPWR VPWR _3831_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7672_ _3771_ VGND VGND VPWR VPWR _3794_ sky130_fd_sc_hd__buf_4
XFILLER_0_117_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6623_ _3221_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9411_ clknet_leaf_74_CLK _0571_ VGND VGND VPWR VPWR RF.registers\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_4884_ net5 VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6554_ RF.registers\[0\]\[24\] _3143_ _3179_ VGND VGND VPWR VPWR _3184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9342_ clknet_leaf_67_CLK _0502_ VGND VGND VPWR VPWR RF.registers\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9273_ clknet_leaf_31_CLK _0433_ VGND VGND VPWR VPWR RF.registers\[23\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_6485_ RF.registers\[17\]\[25\] _3145_ _3135_ VGND VGND VPWR VPWR _3146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5505_ _2259_ _2260_ _2044_ VGND VGND VPWR VPWR _2261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8224_ RF.registers\[1\]\[23\] _3504_ _4083_ VGND VGND VPWR VPWR _4087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5436_ _1828_ _2191_ _1728_ VGND VGND VPWR VPWR _2192_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8155_ _4050_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__clkbuf_1
X_5367_ _1671_ _2110_ _2122_ VGND VGND VPWR VPWR _2123_ sky130_fd_sc_hd__o21ai_4
X_8086_ RF.registers\[20\]\[22\] _3502_ _4011_ VGND VGND VPWR VPWR _4014_ sky130_fd_sc_hd__mux2_1
X_7106_ _3488_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_5298_ RF.registers\[8\]\[3\] RF.registers\[9\]\[3\] RF.registers\[10\]\[3\] RF.registers\[11\]\[3\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2054_ sky130_fd_sc_hd__mux4_1
X_4318_ RF.registers\[8\]\[5\] RF.registers\[9\]\[5\] RF.registers\[10\]\[5\] RF.registers\[11\]\[5\]
+ _1072_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__mux4_1
X_7037_ _3441_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8988_ clknet_leaf_23_CLK _0148_ VGND VGND VPWR VPWR RF.registers\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_7939_ _3935_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6270_ _2991_ _2994_ VGND VGND VPWR VPWR _2995_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5221_ _1766_ _1976_ _1672_ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5152_ _1906_ _1907_ _1745_ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__mux2_1
X_5083_ _1667_ VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__clkbuf_4
X_8911_ clknet_leaf_4_CLK _0071_ VGND VGND VPWR VPWR RF.registers\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8842_ clknet_leaf_83_CLK _0002_ VGND VGND VPWR VPWR RF.registers\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8773_ clknet_leaf_82_CLK _0957_ VGND VGND VPWR VPWR RF.registers\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5985_ _2140_ _2711_ VGND VGND VPWR VPWR _2726_ sky130_fd_sc_hd__or2_1
X_7724_ _3048_ RF.registers\[30\]\[12\] _3819_ VGND VGND VPWR VPWR _3822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4936_ _1691_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_10 _3075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4867_ RF.registers\[24\]\[18\] RF.registers\[25\]\[18\] RF.registers\[26\]\[18\]
+ RF.registers\[27\]\[18\] _1200_ _1202_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__mux4_1
XANTENNA_21 _1712_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7655_ _3785_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6606_ _3212_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7586_ _3046_ RF.registers\[28\]\[11\] _3747_ VGND VGND VPWR VPWR _3749_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6537_ RF.registers\[0\]\[16\] _3126_ _3168_ VGND VGND VPWR VPWR _3175_ sky130_fd_sc_hd__mux2_1
X_9325_ clknet_leaf_8_CLK _0485_ VGND VGND VPWR VPWR RF.registers\[21\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_4798_ RF.registers\[4\]\[10\] RF.registers\[5\]\[10\] RF.registers\[6\]\[10\] RF.registers\[7\]\[10\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6468_ net26 VGND VGND VPWR VPWR _3134_ sky130_fd_sc_hd__buf_2
X_9256_ clknet_leaf_88_CLK _0416_ VGND VGND VPWR VPWR RF.registers\[23\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6399_ _3086_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__clkbuf_1
X_8207_ RF.registers\[1\]\[15\] _3487_ _4072_ VGND VGND VPWR VPWR _4078_ sky130_fd_sc_hd__mux2_1
X_5419_ _1670_ _2166_ _2170_ _2174_ VGND VGND VPWR VPWR _2175_ sky130_fd_sc_hd__a2bb2o_2
X_9187_ clknet_leaf_74_CLK _0347_ VGND VGND VPWR VPWR RF.registers\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8138_ _4041_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__clkbuf_1
X_8069_ RF.registers\[20\]\[14\] _3485_ _4000_ VGND VGND VPWR VPWR _4005_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5770_ _2503_ _2520_ VGND VGND VPWR VPWR _2521_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4721_ RF.registers\[0\]\[13\] RF.registers\[1\]\[13\] RF.registers\[2\]\[13\] RF.registers\[3\]\[13\]
+ _1172_ _1279_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7440_ _3671_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_1
X_4652_ RF.registers\[8\]\[7\] RF.registers\[9\]\[7\] RF.registers\[10\]\[7\] RF.registers\[11\]\[7\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput30 WD3[24] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XFILLER_0_127_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9110_ clknet_leaf_33_CLK _0270_ VGND VGND VPWR VPWR RF.registers\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_4583_ _1335_ _1336_ _1337_ _1338_ _1189_ _1205_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput41 WD3[5] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
X_7371_ _3035_ RF.registers\[26\]\[6\] _3628_ VGND VGND VPWR VPWR _3635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6322_ _3034_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6253_ _2255_ _2910_ _2978_ VGND VGND VPWR VPWR _2979_ sky130_fd_sc_hd__o21ai_1
X_9041_ clknet_leaf_19_CLK _0201_ VGND VGND VPWR VPWR RF.registers\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5204_ _1839_ _1959_ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__nor2_1
X_6184_ _2408_ _2906_ _2907_ _2913_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__o22a_1
X_5135_ RF.registers\[8\]\[31\] RF.registers\[9\]\[31\] RF.registers\[10\]\[31\] RF.registers\[11\]\[31\]
+ _1882_ _1884_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5066_ _1782_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__clkbuf_8
X_8825_ clknet_leaf_50_CLK _1009_ VGND VGND VPWR VPWR RF.registers\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8756_ clknet_leaf_43_CLK _0940_ VGND VGND VPWR VPWR RF.registers\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5968_ _1464_ _1480_ _2657_ _2411_ VGND VGND VPWR VPWR _2710_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7707_ _3031_ RF.registers\[30\]\[4\] _3808_ VGND VGND VPWR VPWR _3813_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4919_ _1674_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5899_ _2642_ _2643_ VGND VGND VPWR VPWR _2644_ sky130_fd_sc_hd__nand2_1
X_8687_ clknet_leaf_11_CLK _0871_ VGND VGND VPWR VPWR RF.registers\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7638_ _3776_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7569_ _3029_ RF.registers\[28\]\[3\] _3736_ VGND VGND VPWR VPWR _3740_ sky130_fd_sc_hd__mux2_1
X_9308_ clknet_leaf_23_CLK _0468_ VGND VGND VPWR VPWR RF.registers\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_9239_ clknet_leaf_50_CLK _0399_ VGND VGND VPWR VPWR RF.registers\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6940_ RF.registers\[4\]\[12\] _3118_ _3387_ VGND VGND VPWR VPWR _3390_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6871_ _3353_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__clkbuf_1
X_9590_ clknet_leaf_34_CLK _0750_ VGND VGND VPWR VPWR RF.registers\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_5822_ _2474_ _2469_ _1126_ VGND VGND VPWR VPWR _2571_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8610_ clknet_leaf_76_CLK _0794_ VGND VGND VPWR VPWR RF.registers\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_5753_ _2496_ _2502_ _2504_ VGND VGND VPWR VPWR _2505_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8541_ RF.registers\[10\]\[13\] net18 _4244_ VGND VGND VPWR VPWR _4254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4704_ RF.registers\[8\]\[12\] RF.registers\[9\]\[12\] RF.registers\[10\]\[12\] RF.registers\[11\]\[12\]
+ _1181_ _1183_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5684_ _1841_ _2347_ VGND VGND VPWR VPWR _2438_ sky130_fd_sc_hd__or2b_1
X_8472_ _4218_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__clkbuf_1
X_7423_ _3087_ RF.registers\[26\]\[31\] _3627_ VGND VGND VPWR VPWR _3662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4635_ RF.registers\[8\]\[6\] RF.registers\[9\]\[6\] RF.registers\[10\]\[6\] RF.registers\[11\]\[6\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7354_ _3087_ RF.registers\[31\]\[31\] _3590_ VGND VGND VPWR VPWR _3625_ sky130_fd_sc_hd__mux2_1
X_4566_ _1320_ _1321_ _1198_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6305_ _3022_ VGND VGND VPWR VPWR _3023_ sky130_fd_sc_hd__buf_6
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7285_ _3588_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_4497_ _1251_ _1252_ _1211_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__mux2_1
X_9024_ clknet_leaf_74_CLK _0184_ VGND VGND VPWR VPWR RF.registers\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6236_ _1087_ _2960_ _2961_ _2962_ _1127_ VGND VGND VPWR VPWR _2963_ sky130_fd_sc_hd__a32o_1
X_6167_ _2105_ _2754_ _2897_ _1087_ VGND VGND VPWR VPWR _2898_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5118_ _1777_ _1865_ _1869_ _1873_ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__o2bb2a_2
X_6098_ _2830_ _2832_ _2503_ VGND VGND VPWR VPWR _2833_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_123_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5049_ RF.registers\[20\]\[18\] RF.registers\[21\]\[18\] RF.registers\[22\]\[18\]
+ RF.registers\[23\]\[18\] _1719_ _1722_ VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_28_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8808_ clknet_leaf_81_CLK _0992_ VGND VGND VPWR VPWR RF.registers\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8739_ clknet_leaf_76_CLK _0923_ VGND VGND VPWR VPWR RF.registers\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4420_ RF.registers\[20\]\[29\] RF.registers\[21\]\[29\] RF.registers\[22\]\[29\]
+ RF.registers\[23\]\[29\] _1173_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4351_ _1034_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4282_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__buf_4
X_7070_ net40 VGND VGND VPWR VPWR _3464_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _2757_ _2731_ _2758_ _2759_ VGND VGND VPWR VPWR _2760_ sky130_fd_sc_hd__a211o_1
X_7972_ _3953_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__clkbuf_1
X_6923_ RF.registers\[4\]\[4\] _3101_ _3376_ VGND VGND VPWR VPWR _3381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6854_ _3344_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5805_ _1666_ _2554_ VGND VGND VPWR VPWR _2555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6785_ RF.registers\[6\]\[3\] _3099_ _3304_ VGND VGND VPWR VPWR _3308_ sky130_fd_sc_hd__mux2_1
X_9573_ clknet_leaf_80_CLK _0733_ VGND VGND VPWR VPWR RF.registers\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5736_ _2040_ _2486_ _2487_ _1962_ VGND VGND VPWR VPWR _2488_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8524_ _4245_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_33_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5667_ _2333_ VGND VGND VPWR VPWR _2421_ sky130_fd_sc_hd__buf_2
XFILLER_0_60_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8455_ _4209_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4618_ RF.registers\[20\]\[24\] RF.registers\[21\]\[24\] RF.registers\[22\]\[24\]
+ RF.registers\[23\]\[24\] _1360_ _1361_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__mux4_1
X_7406_ _3653_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5598_ _1668_ _2247_ VGND VGND VPWR VPWR _2353_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8386_ RF.registers\[12\]\[3\] _3462_ _4169_ VGND VGND VPWR VPWR _4173_ sky130_fd_sc_hd__mux2_1
X_4549_ _1303_ _1304_ _1259_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__mux2_1
X_7337_ _3616_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7268_ _3069_ RF.registers\[29\]\[22\] _3577_ VGND VGND VPWR VPWR _3580_ sky130_fd_sc_hd__mux2_1
X_6219_ _2105_ _2802_ _2946_ _1085_ VGND VGND VPWR VPWR _2947_ sky130_fd_sc_hd__o211a_1
X_9007_ clknet_leaf_5_CLK _0167_ VGND VGND VPWR VPWR RF.registers\[31\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_7199_ _3542_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload19 clknet_leaf_8_CLK VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_11_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6570_ net13 net12 net11 VGND VGND VPWR VPWR _3192_ sky130_fd_sc_hd__and3b_2
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5521_ _2273_ _2274_ _2275_ _2276_ _1711_ _1716_ VGND VGND VPWR VPWR _2277_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8240_ RF.registers\[1\]\[31\] _3452_ _4060_ VGND VGND VPWR VPWR _4095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5452_ _2206_ _2207_ _1738_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__mux2_1
X_8171_ _4058_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__clkbuf_1
X_5383_ _1828_ _2138_ _1728_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4403_ RF.registers\[12\]\[0\] RF.registers\[13\]\[0\] RF.registers\[14\]\[0\] RF.registers\[15\]\[0\]
+ _1149_ _1028_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7122_ _3499_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_4334_ _1043_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__buf_4
X_7053_ net38 VGND VGND VPWR VPWR _3452_ sky130_fd_sc_hd__buf_2
X_6004_ _1874_ _2743_ VGND VGND VPWR VPWR _2744_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7955_ RF.registers\[18\]\[25\] _3508_ _3938_ VGND VGND VPWR VPWR _3944_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7886_ _3907_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6906_ _3371_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6837_ RF.registers\[6\]\[28\] _3011_ _3326_ VGND VGND VPWR VPWR _3335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9556_ clknet_leaf_42_CLK _0716_ VGND VGND VPWR VPWR RF.registers\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8507_ _4236_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__clkbuf_1
X_6768_ _3081_ RF.registers\[14\]\[28\] _3289_ VGND VGND VPWR VPWR _3298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6699_ _3261_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5719_ _2347_ _1169_ _1905_ VGND VGND VPWR VPWR _2472_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9487_ clknet_leaf_6_CLK _0647_ VGND VGND VPWR VPWR RF.registers\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8438_ RF.registers\[12\]\[28\] net34 _4191_ VGND VGND VPWR VPWR _4200_ sky130_fd_sc_hd__mux2_1
X_8369_ _4163_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_131_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 A2[2] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7740_ _3807_ VGND VGND VPWR VPWR _3830_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4952_ _1707_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4883_ _1638_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__buf_2
X_7671_ _3793_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6622_ _3071_ RF.registers\[15\]\[23\] _3217_ VGND VGND VPWR VPWR _3221_ sky130_fd_sc_hd__mux2_1
X_9410_ clknet_leaf_76_CLK _0570_ VGND VGND VPWR VPWR RF.registers\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6553_ _3183_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9341_ clknet_leaf_18_CLK _0501_ VGND VGND VPWR VPWR RF.registers\[21\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6484_ net31 VGND VGND VPWR VPWR _3145_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9272_ clknet_leaf_39_CLK _0432_ VGND VGND VPWR VPWR RF.registers\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5504_ RF.registers\[24\]\[6\] RF.registers\[25\]\[6\] RF.registers\[26\]\[6\] RF.registers\[27\]\[6\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2260_ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8223_ _4086_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5435_ _2189_ _2190_ _1738_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8154_ RF.registers\[24\]\[22\] _3502_ _4047_ VGND VGND VPWR VPWR _4050_ sky130_fd_sc_hd__mux2_1
X_5366_ _2112_ _2116_ _2121_ _1828_ _1728_ VGND VGND VPWR VPWR _2122_ sky130_fd_sc_hd__a221o_1
X_8085_ _4013_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__clkbuf_1
X_7105_ RF.registers\[19\]\[15\] _3487_ _3477_ VGND VGND VPWR VPWR _3488_ sky130_fd_sc_hd__mux2_1
X_4317_ _1043_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__buf_4
X_5297_ _2052_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__buf_4
X_7036_ RF.registers\[3\]\[25\] _3145_ _3435_ VGND VGND VPWR VPWR _3441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8987_ clknet_leaf_46_CLK _0147_ VGND VGND VPWR VPWR RF.registers\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7938_ RF.registers\[18\]\[17\] _3491_ _3927_ VGND VGND VPWR VPWR _3935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7869_ _3898_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9539_ clknet_leaf_76_CLK _0699_ VGND VGND VPWR VPWR RF.registers\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5220_ _1974_ _1975_ _1745_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5151_ RF.registers\[16\]\[30\] RF.registers\[17\]\[30\] RF.registers\[18\]\[30\]
+ RF.registers\[19\]\[30\] _1895_ _1897_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__mux4_1
X_5082_ _1671_ _1829_ _1833_ _1837_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__a2bb2o_2
X_8910_ clknet_leaf_21_CLK _0070_ VGND VGND VPWR VPWR RF.registers\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8841_ clknet_leaf_82_CLK _0001_ VGND VGND VPWR VPWR RF.registers\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8772_ clknet_leaf_78_CLK _0956_ VGND VGND VPWR VPWR RF.registers\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_5984_ _2123_ _2724_ VGND VGND VPWR VPWR _2725_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7723_ _3821_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4935_ _1690_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_11 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4866_ RF.registers\[28\]\[18\] RF.registers\[29\]\[18\] RF.registers\[30\]\[18\]
+ RF.registers\[31\]\[18\] _1200_ _1202_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__mux4_1
X_7654_ RF.registers\[2\]\[11\] _3479_ _3783_ VGND VGND VPWR VPWR _3785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6605_ _3054_ RF.registers\[15\]\[15\] _3206_ VGND VGND VPWR VPWR _3212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7585_ _3748_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4797_ _1038_ _1552_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6536_ _3174_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9324_ clknet_leaf_2_CLK _0484_ VGND VGND VPWR VPWR RF.registers\[21\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6467_ _3133_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__clkbuf_1
X_9255_ clknet_leaf_58_CLK _0415_ VGND VGND VPWR VPWR RF.registers\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_6398_ _3085_ RF.registers\[22\]\[30\] _3022_ VGND VGND VPWR VPWR _3086_ sky130_fd_sc_hd__mux2_1
X_8206_ _4077_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__clkbuf_1
X_9186_ clknet_leaf_93_CLK _0346_ VGND VGND VPWR VPWR RF.registers\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_5418_ _1828_ _2173_ _1728_ VGND VGND VPWR VPWR _2174_ sky130_fd_sc_hd__a21oi_1
X_5349_ _2104_ VGND VGND VPWR VPWR _2105_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8137_ RF.registers\[24\]\[14\] _3485_ _4036_ VGND VGND VPWR VPWR _4041_ sky130_fd_sc_hd__mux2_1
X_8068_ _4004_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__clkbuf_1
X_7019_ RF.registers\[3\]\[17\] _3128_ _3424_ VGND VGND VPWR VPWR _3432_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4720_ RF.registers\[4\]\[13\] RF.registers\[5\]\[13\] RF.registers\[6\]\[13\] RF.registers\[7\]\[13\]
+ _1172_ _1279_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4651_ RF.registers\[12\]\[7\] RF.registers\[13\]\[7\] RF.registers\[14\]\[7\] RF.registers\[15\]\[7\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__mux4_1
Xinput31 WD3[25] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
Xinput20 WD3[15] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4582_ RF.registers\[20\]\[30\] RF.registers\[21\]\[30\] RF.registers\[22\]\[30\]
+ RF.registers\[23\]\[30\] _1267_ _1268_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7370_ _3634_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
Xinput42 WD3[6] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6321_ _3033_ RF.registers\[22\]\[5\] _3023_ VGND VGND VPWR VPWR _3034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6252_ _2104_ _2849_ _2977_ _1086_ VGND VGND VPWR VPWR _2978_ sky130_fd_sc_hd__o211a_1
X_9040_ clknet_leaf_6_CLK _0200_ VGND VGND VPWR VPWR RF.registers\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5203_ _1842_ _1958_ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__nor2_1
X_6183_ _2504_ _2908_ _2912_ VGND VGND VPWR VPWR _2913_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5134_ _1885_ _1886_ _1887_ _1888_ _1889_ _1773_ VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__mux4_1
X_5065_ _1758_ _1820_ VGND VGND VPWR VPWR _1821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8824_ clknet_leaf_40_CLK _1008_ VGND VGND VPWR VPWR RF.registers\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8755_ clknet_leaf_30_CLK _0939_ VGND VGND VPWR VPWR RF.registers\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5967_ _2550_ _2591_ _2708_ VGND VGND VPWR VPWR _2709_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8686_ clknet_leaf_15_CLK _0870_ VGND VGND VPWR VPWR RF.registers\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7706_ _3812_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__clkbuf_1
X_4918_ _1673_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_23_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5898_ _2193_ _2640_ _2641_ VGND VGND VPWR VPWR _2643_ sky130_fd_sc_hd__nand3_1
X_7637_ RF.registers\[2\]\[3\] _3462_ _3772_ VGND VGND VPWR VPWR _3776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4849_ _1603_ _1604_ _1178_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7568_ _3739_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
X_9307_ clknet_leaf_46_CLK _0467_ VGND VGND VPWR VPWR RF.registers\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_7499_ _3027_ RF.registers\[27\]\[2\] _3700_ VGND VGND VPWR VPWR _3703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6519_ _3165_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__clkbuf_1
X_9238_ clknet_leaf_34_CLK _0398_ VGND VGND VPWR VPWR RF.registers\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9169_ clknet_leaf_40_CLK _0329_ VGND VGND VPWR VPWR RF.registers\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6870_ RF.registers\[5\]\[11\] _3116_ _3351_ VGND VGND VPWR VPWR _3353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5821_ _2039_ _2251_ VGND VGND VPWR VPWR _2570_ sky130_fd_sc_hd__and2_1
X_5752_ _2503_ VGND VGND VPWR VPWR _2504_ sky130_fd_sc_hd__buf_2
X_8540_ _4253_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4703_ _1287_ _1458_ _1088_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__o21a_1
X_5683_ _2036_ _1757_ _2347_ VGND VGND VPWR VPWR _2437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8471_ RF.registers\[11\]\[11\] net16 _4216_ VGND VGND VPWR VPWR _4218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7422_ _3661_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4634_ _1386_ _1387_ _1388_ _1389_ _1048_ _1088_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_96_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7353_ _3624_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
X_4565_ RF.registers\[24\]\[31\] RF.registers\[25\]\[31\] RF.registers\[26\]\[31\]
+ RF.registers\[27\]\[31\] _1200_ _1202_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6304_ _3020_ _3021_ VGND VGND VPWR VPWR _3022_ sky130_fd_sc_hd__nand2_2
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7284_ _3085_ RF.registers\[29\]\[30\] _3554_ VGND VGND VPWR VPWR _3588_ sky130_fd_sc_hd__mux2_1
X_4496_ RF.registers\[0\]\[20\] RF.registers\[1\]\[20\] RF.registers\[2\]\[20\] RF.registers\[3\]\[20\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9023_ clknet_leaf_73_CLK _0183_ VGND VGND VPWR VPWR RF.registers\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_6235_ _2102_ _2692_ VGND VGND VPWR VPWR _2962_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6166_ _2255_ _2821_ _2896_ _2337_ VGND VGND VPWR VPWR _2897_ sky130_fd_sc_hd__o22a_1
X_6097_ _2806_ _2827_ VGND VGND VPWR VPWR _2832_ sky130_fd_sc_hd__nor2_1
X_5117_ _1700_ _1872_ _1671_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__o21ai_1
X_5048_ _1757_ _1802_ _1803_ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8807_ clknet_leaf_60_CLK _0991_ VGND VGND VPWR VPWR RF.registers\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8738_ clknet_leaf_91_CLK _0922_ VGND VGND VPWR VPWR RF.registers\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6999_ _3421_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8669_ clknet_leaf_39_CLK _0853_ VGND VGND VPWR VPWR RF.registers\[0\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4350_ RF.registers\[0\]\[3\] RF.registers\[1\]\[3\] RF.registers\[2\]\[3\] RF.registers\[3\]\[3\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4281_ net7 VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _2102_ _2406_ VGND VGND VPWR VPWR _2759_ sky130_fd_sc_hd__nor2_1
X_7971_ _3089_ RF.registers\[21\]\[0\] _3952_ VGND VGND VPWR VPWR _3953_ sky130_fd_sc_hd__mux2_1
X_6922_ _3380_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6853_ RF.registers\[5\]\[3\] _3099_ _3340_ VGND VGND VPWR VPWR _3344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5804_ _2442_ _2487_ _2553_ _2040_ VGND VGND VPWR VPWR _2554_ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6784_ _3307_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9572_ clknet_leaf_88_CLK _0732_ VGND VGND VPWR VPWR RF.registers\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5735_ _2039_ _2251_ VGND VGND VPWR VPWR _2487_ sky130_fd_sc_hd__nand2_1
X_8523_ RF.registers\[10\]\[4\] net40 _4244_ VGND VGND VPWR VPWR _4245_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5666_ _2363_ _2417_ _2419_ VGND VGND VPWR VPWR _2420_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8454_ RF.registers\[11\]\[3\] net39 _4205_ VGND VGND VPWR VPWR _4209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4617_ RF.registers\[16\]\[24\] RF.registers\[17\]\[24\] RF.registers\[18\]\[24\]
+ RF.registers\[19\]\[24\] _1360_ _1361_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__mux4_1
X_7405_ _3069_ RF.registers\[26\]\[22\] _3650_ VGND VGND VPWR VPWR _3653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5597_ _1839_ _2211_ VGND VGND VPWR VPWR _2352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8385_ _4172_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4548_ RF.registers\[24\]\[27\] RF.registers\[25\]\[27\] RF.registers\[26\]\[27\]
+ RF.registers\[27\]\[27\] _1262_ _1263_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__mux4_1
X_7336_ _3069_ RF.registers\[31\]\[22\] _3613_ VGND VGND VPWR VPWR _3616_ sky130_fd_sc_hd__mux2_1
X_7267_ _3579_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
X_4479_ _1233_ _1234_ _1189_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__mux2_1
X_6218_ _2255_ _2867_ _2945_ _2337_ VGND VGND VPWR VPWR _2946_ sky130_fd_sc_hd__o22a_1
X_9006_ clknet_leaf_20_CLK _0166_ VGND VGND VPWR VPWR RF.registers\[31\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7198_ RF.registers\[7\]\[22\] _3502_ _3539_ VGND VGND VPWR VPWR _3542_ sky130_fd_sc_hd__mux2_1
X_6149_ _1731_ _2853_ VGND VGND VPWR VPWR _2881_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_107_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5520_ RF.registers\[20\]\[7\] RF.registers\[21\]\[7\] RF.registers\[22\]\[7\] RF.registers\[23\]\[7\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5451_ RF.registers\[0\]\[10\] RF.registers\[1\]\[10\] RF.registers\[2\]\[10\] RF.registers\[3\]\[10\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__mux4_1
X_8170_ RF.registers\[24\]\[30\] _3450_ _4024_ VGND VGND VPWR VPWR _4058_ sky130_fd_sc_hd__mux2_1
X_5382_ _2136_ _2137_ _1738_ VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4402_ RF.registers\[8\]\[0\] RF.registers\[9\]\[0\] RF.registers\[10\]\[0\] RF.registers\[11\]\[0\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__mux4_1
X_7121_ RF.registers\[19\]\[20\] _3497_ _3498_ VGND VGND VPWR VPWR _3499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4333_ _1041_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__clkbuf_8
X_7052_ _3451_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
X_6003_ _1587_ _2742_ VGND VGND VPWR VPWR _2743_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7954_ _3943_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_120_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ RF.registers\[5\]\[28\] _3011_ _3362_ VGND VGND VPWR VPWR _3371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7885_ _3143_ RF.registers\[23\]\[24\] _3902_ VGND VGND VPWR VPWR _3907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6836_ _3334_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6767_ _3297_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__clkbuf_1
X_9555_ clknet_leaf_29_CLK _0715_ VGND VGND VPWR VPWR RF.registers\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8506_ RF.registers\[11\]\[28\] net34 _4227_ VGND VGND VPWR VPWR _4236_ sky130_fd_sc_hd__mux2_1
X_5718_ _2469_ _2470_ _2251_ VGND VGND VPWR VPWR _2471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6698_ RF.registers\[8\]\[27\] _3009_ _3253_ VGND VGND VPWR VPWR _3261_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9486_ clknet_leaf_20_CLK _0646_ VGND VGND VPWR VPWR RF.registers\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8437_ _4199_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__clkbuf_1
X_5649_ _2397_ _2403_ _1125_ VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8368_ RF.registers\[16\]\[27\] _3444_ _4155_ VGND VGND VPWR VPWR _4163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7319_ _3052_ RF.registers\[31\]\[14\] _3602_ VGND VGND VPWR VPWR _3607_ sky130_fd_sc_hd__mux2_1
X_8299_ _4126_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput7 A2[3] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4951_ _1706_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__buf_4
X_4882_ _1637_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__clkbuf_4
X_7670_ RF.registers\[2\]\[19\] _3495_ _3783_ VGND VGND VPWR VPWR _3793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6621_ _3220_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9340_ clknet_leaf_18_CLK _0500_ VGND VGND VPWR VPWR RF.registers\[21\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6552_ RF.registers\[0\]\[23\] _3141_ _3179_ VGND VGND VPWR VPWR _3183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9271_ clknet_leaf_32_CLK _0431_ VGND VGND VPWR VPWR RF.registers\[23\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6483_ _3144_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5503_ RF.registers\[28\]\[6\] RF.registers\[29\]\[6\] RF.registers\[30\]\[6\] RF.registers\[31\]\[6\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8222_ RF.registers\[1\]\[22\] _3502_ _4083_ VGND VGND VPWR VPWR _4086_ sky130_fd_sc_hd__mux2_1
X_5434_ RF.registers\[0\]\[11\] RF.registers\[1\]\[11\] RF.registers\[2\]\[11\] RF.registers\[3\]\[11\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__mux4_1
X_8153_ _4049_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7104_ net20 VGND VGND VPWR VPWR _3487_ sky130_fd_sc_hd__buf_2
XFILLER_0_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5365_ _2119_ _2120_ _1738_ VGND VGND VPWR VPWR _2121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8084_ RF.registers\[20\]\[21\] _3500_ _4011_ VGND VGND VPWR VPWR _4013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5296_ _1690_ VGND VGND VPWR VPWR _2052_ sky130_fd_sc_hd__clkbuf_4
X_4316_ _1041_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__buf_4
X_7035_ _3440_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8986_ clknet_leaf_25_CLK _0146_ VGND VGND VPWR VPWR RF.registers\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_7937_ _3934_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_67_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7868_ _3126_ RF.registers\[23\]\[16\] _3891_ VGND VGND VPWR VPWR _3898_ sky130_fd_sc_hd__mux2_1
X_6819_ _3325_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7799_ _3861_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9538_ clknet_leaf_91_CLK _0698_ VGND VGND VPWR VPWR RF.registers\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9469_ clknet_leaf_15_CLK _0629_ VGND VGND VPWR VPWR RF.registers\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_94_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5150_ RF.registers\[20\]\[30\] RF.registers\[21\]\[30\] RF.registers\[22\]\[30\]
+ RF.registers\[23\]\[30\] _1895_ _1897_ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__mux4_1
X_5081_ _1717_ _1836_ _1729_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_88_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8840_ clknet_leaf_79_CLK _0000_ VGND VGND VPWR VPWR RF.registers\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5983_ _1511_ _2723_ VGND VGND VPWR VPWR _2724_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8771_ clknet_leaf_79_CLK _0955_ VGND VGND VPWR VPWR RF.registers\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_4934_ _1642_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__buf_4
X_7722_ _3046_ RF.registers\[30\]\[11\] _3819_ VGND VGND VPWR VPWR _3821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_12 _3132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4865_ _1619_ _1620_ _1259_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__mux2_1
X_7653_ _3784_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7584_ _3043_ RF.registers\[28\]\[10\] _3747_ VGND VGND VPWR VPWR _3748_ sky130_fd_sc_hd__mux2_1
X_4796_ _1550_ _1551_ _1047_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__mux2_1
X_6604_ _3211_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6535_ RF.registers\[0\]\[15\] _3124_ _3168_ VGND VGND VPWR VPWR _3174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9323_ clknet_leaf_1_CLK _0483_ VGND VGND VPWR VPWR RF.registers\[21\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9254_ clknet_leaf_62_CLK _0414_ VGND VGND VPWR VPWR RF.registers\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6466_ RF.registers\[17\]\[19\] _3132_ _3114_ VGND VGND VPWR VPWR _3133_ sky130_fd_sc_hd__mux2_1
X_8205_ RF.registers\[1\]\[14\] _3485_ _4072_ VGND VGND VPWR VPWR _4077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6397_ net37 VGND VGND VPWR VPWR _3085_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9185_ clknet_leaf_97_CLK _0345_ VGND VGND VPWR VPWR RF.registers\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5417_ _2171_ _2172_ _1738_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5348_ _1111_ VGND VGND VPWR VPWR _2104_ sky130_fd_sc_hd__clkbuf_4
X_8136_ _4040_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8067_ RF.registers\[20\]\[13\] _3483_ _4000_ VGND VGND VPWR VPWR _4004_ sky130_fd_sc_hd__mux2_1
X_5279_ _1799_ _2034_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__and2_1
X_7018_ _3431_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
X_8969_ clknet_leaf_1_CLK _0129_ VGND VGND VPWR VPWR RF.registers\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4650_ _1402_ _1405_ _1038_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput21 WD3[16] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput10 A3[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput32 WD3[26] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
X_4581_ RF.registers\[16\]\[30\] RF.registers\[17\]\[30\] RF.registers\[18\]\[30\]
+ RF.registers\[19\]\[30\] _1267_ _1268_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput43 WD3[7] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
X_6320_ net41 VGND VGND VPWR VPWR _3033_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6251_ _1944_ _2975_ _2976_ VGND VGND VPWR VPWR _2977_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_30_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_30_CLK sky130_fd_sc_hd__clkbuf_8
X_5202_ _1777_ _1949_ _1957_ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__a21oi_4
X_6182_ _2530_ _2779_ _2911_ _1087_ VGND VGND VPWR VPWR _2912_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5133_ _1713_ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5064_ _1671_ _1811_ _1815_ _1819_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__a2bb2o_2
X_8823_ clknet_leaf_49_CLK _1007_ VGND VGND VPWR VPWR RF.registers\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8754_ clknet_leaf_43_CLK _0938_ VGND VGND VPWR VPWR RF.registers\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5966_ _2553_ _2588_ _2679_ _2442_ _2333_ VGND VGND VPWR VPWR _2708_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_97_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_97_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5897_ _2640_ _2641_ _2193_ VGND VGND VPWR VPWR _2642_ sky130_fd_sc_hd__a21o_1
X_8685_ clknet_leaf_10_CLK _0869_ VGND VGND VPWR VPWR RF.registers\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_7705_ _3029_ RF.registers\[30\]\[3\] _3808_ VGND VGND VPWR VPWR _3812_ sky130_fd_sc_hd__mux2_1
X_4917_ _1641_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_23_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4848_ RF.registers\[16\]\[19\] RF.registers\[17\]\[19\] RF.registers\[18\]\[19\]
+ RF.registers\[19\]\[19\] _1220_ _1222_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__mux4_1
X_7636_ _3775_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9306_ clknet_leaf_24_CLK _0466_ VGND VGND VPWR VPWR RF.registers\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_7567_ _3027_ RF.registers\[28\]\[2\] _3736_ VGND VGND VPWR VPWR _3739_ sky130_fd_sc_hd__mux2_1
X_4779_ _1047_ _1534_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7498_ _3702_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
X_6518_ RF.registers\[0\]\[7\] _3107_ _3157_ VGND VGND VPWR VPWR _3165_ sky130_fd_sc_hd__mux2_1
X_9237_ clknet_leaf_34_CLK _0397_ VGND VGND VPWR VPWR RF.registers\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6449_ _3121_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_21_CLK sky130_fd_sc_hd__clkbuf_8
X_9168_ clknet_leaf_57_CLK _0328_ VGND VGND VPWR VPWR RF.registers\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8119_ _4031_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9099_ clknet_leaf_98_CLK _0259_ VGND VGND VPWR VPWR RF.registers\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_88_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_88_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_12_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5820_ _2568_ VGND VGND VPWR VPWR _2569_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_79_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_79_CLK sky130_fd_sc_hd__clkbuf_8
X_5751_ net48 VGND VGND VPWR VPWR _2503_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8470_ _4217_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__clkbuf_1
X_4702_ RF.registers\[0\]\[12\] RF.registers\[1\]\[12\] RF.registers\[2\]\[12\] RF.registers\[3\]\[12\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7421_ _3085_ RF.registers\[26\]\[30\] _3627_ VGND VGND VPWR VPWR _3661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5682_ _2105_ _2427_ _2435_ VGND VGND VPWR VPWR _2436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4633_ RF.registers\[20\]\[6\] RF.registers\[21\]\[6\] RF.registers\[22\]\[6\] RF.registers\[23\]\[6\]
+ _1219_ _1221_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7352_ _3085_ RF.registers\[31\]\[30\] _3590_ VGND VGND VPWR VPWR _3624_ sky130_fd_sc_hd__mux2_1
X_4564_ RF.registers\[28\]\[31\] RF.registers\[29\]\[31\] RF.registers\[30\]\[31\]
+ RF.registers\[31\]\[31\] _1200_ _1202_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__mux4_1
X_7283_ _3587_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
X_6303_ net12 net11 net13 VGND VGND VPWR VPWR _3021_ sky130_fd_sc_hd__and3b_2
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4495_ RF.registers\[4\]\[20\] RF.registers\[5\]\[20\] RF.registers\[6\]\[20\] RF.registers\[7\]\[20\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__mux4_1
X_6234_ _1111_ _2822_ _2896_ _2254_ VGND VGND VPWR VPWR _2961_ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9022_ clknet_leaf_69_CLK _0182_ VGND VGND VPWR VPWR RF.registers\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6165_ _2857_ _2895_ _2327_ VGND VGND VPWR VPWR _2896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6096_ _2830_ VGND VGND VPWR VPWR _2831_ sky130_fd_sc_hd__inv_2
X_5116_ _1870_ _1871_ _1726_ VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__mux2_1
X_5047_ _1145_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_123_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8806_ clknet_leaf_61_CLK _0990_ VGND VGND VPWR VPWR RF.registers\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_40_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6998_ RF.registers\[3\]\[7\] _3107_ _3413_ VGND VGND VPWR VPWR _3421_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5949_ _2378_ _2381_ _2178_ VGND VGND VPWR VPWR _2692_ sky130_fd_sc_hd__mux2_1
X_8737_ clknet_leaf_93_CLK _0921_ VGND VGND VPWR VPWR RF.registers\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8668_ clknet_leaf_38_CLK _0852_ VGND VGND VPWR VPWR RF.registers\[0\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8599_ clknet_leaf_32_CLK _0783_ VGND VGND VPWR VPWR RF.registers\[22\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_7619_ _3079_ RF.registers\[28\]\[27\] _3758_ VGND VGND VPWR VPWR _3766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_1_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_1_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4280_ _1035_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7970_ _3951_ VGND VGND VPWR VPWR _3952_ sky130_fd_sc_hd__buf_6
X_6921_ RF.registers\[4\]\[3\] _3099_ _3376_ VGND VGND VPWR VPWR _3380_ sky130_fd_sc_hd__mux2_1
X_6852_ _3343_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5803_ _2443_ _2437_ _1879_ VGND VGND VPWR VPWR _2553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9571_ clknet_leaf_77_CLK _0731_ VGND VGND VPWR VPWR RF.registers\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8522_ _3006_ VGND VGND VPWR VPWR _4244_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6783_ RF.registers\[6\]\[2\] _3097_ _3304_ VGND VGND VPWR VPWR _3307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5734_ _2037_ _1804_ _2251_ VGND VGND VPWR VPWR _2486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5665_ _1147_ _2418_ VGND VGND VPWR VPWR _2419_ sky130_fd_sc_hd__nand2_1
X_8453_ _4208_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4616_ RF.registers\[28\]\[24\] RF.registers\[29\]\[24\] RF.registers\[30\]\[24\]
+ RF.registers\[31\]\[24\] _1360_ _1361_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__mux4_1
X_7404_ _3652_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8384_ RF.registers\[12\]\[2\] _3460_ _4169_ VGND VGND VPWR VPWR _4172_ sky130_fd_sc_hd__mux2_1
X_7335_ _3615_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5596_ _2349_ _2350_ VGND VGND VPWR VPWR _2351_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4547_ RF.registers\[28\]\[27\] RF.registers\[29\]\[27\] RF.registers\[30\]\[27\]
+ RF.registers\[31\]\[27\] _1262_ _1263_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__mux4_1
X_7266_ _3067_ RF.registers\[29\]\[21\] _3577_ VGND VGND VPWR VPWR _3579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4478_ RF.registers\[12\]\[28\] RF.registers\[13\]\[28\] RF.registers\[14\]\[28\]
+ RF.registers\[15\]\[28\] _1182_ _1184_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__mux4_1
X_7197_ _3541_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6217_ _2909_ _2944_ _2178_ VGND VGND VPWR VPWR _2945_ sky130_fd_sc_hd__mux2_1
X_9005_ clknet_leaf_3_CLK _0165_ VGND VGND VPWR VPWR RF.registers\[31\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6148_ _1731_ _2853_ _2838_ VGND VGND VPWR VPWR _2880_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _2667_ _2745_ VGND VGND VPWR VPWR _2815_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5450_ RF.registers\[4\]\[10\] RF.registers\[5\]\[10\] RF.registers\[6\]\[10\] RF.registers\[7\]\[10\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4401_ _1038_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5381_ RF.registers\[0\]\[14\] RF.registers\[1\]\[14\] RF.registers\[2\]\[14\] RF.registers\[3\]\[14\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2137_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7120_ _3455_ VGND VGND VPWR VPWR _3498_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4332_ _1050_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__buf_4
X_7051_ RF.registers\[3\]\[30\] _3450_ _3412_ VGND VGND VPWR VPWR _3451_ sky130_fd_sc_hd__mux2_1
X_6002_ _1512_ _2658_ _2741_ VGND VGND VPWR VPWR _2742_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7953_ RF.registers\[18\]\[24\] _3506_ _3938_ VGND VGND VPWR VPWR _3943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6904_ _3370_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7884_ _3906_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6835_ RF.registers\[6\]\[27\] _3009_ _3326_ VGND VGND VPWR VPWR _3334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6766_ _3079_ RF.registers\[14\]\[27\] _3289_ VGND VGND VPWR VPWR _3297_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_114_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9554_ clknet_leaf_41_CLK _0714_ VGND VGND VPWR VPWR RF.registers\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8505_ _4235_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__clkbuf_1
X_5717_ _2396_ _2400_ _1877_ VGND VGND VPWR VPWR _2470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6697_ _3260_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__clkbuf_1
X_9485_ clknet_leaf_4_CLK _0645_ VGND VGND VPWR VPWR RF.registers\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8436_ RF.registers\[12\]\[27\] net33 _4191_ VGND VGND VPWR VPWR _4199_ sky130_fd_sc_hd__mux2_1
X_5648_ _2400_ _2402_ _1145_ VGND VGND VPWR VPWR _2403_ sky130_fd_sc_hd__mux2_1
X_8367_ _4162_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__clkbuf_1
X_5579_ _1128_ _1663_ _2330_ _2334_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__o211ai_2
XFILLER_0_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8298_ _3002_ RF.registers\[13\]\[26\] _4119_ VGND VGND VPWR VPWR _4126_ sky130_fd_sc_hd__mux2_1
X_7318_ _3606_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
X_7249_ _3050_ RF.registers\[29\]\[13\] _3566_ VGND VGND VPWR VPWR _3570_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_123_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 A2[4] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_4
XFILLER_0_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4950_ _1678_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _1350_ _1385_ _1448_ _1636_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_86_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6620_ _3069_ RF.registers\[15\]\[22\] _3217_ VGND VGND VPWR VPWR _3220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6551_ _3182_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__clkbuf_1
X_5502_ _2256_ _2257_ _2044_ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9270_ clknet_leaf_48_CLK _0430_ VGND VGND VPWR VPWR RF.registers\[23\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6482_ RF.registers\[17\]\[24\] _3143_ _3135_ VGND VGND VPWR VPWR _3144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8221_ _4085_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5433_ RF.registers\[4\]\[11\] RF.registers\[5\]\[11\] RF.registers\[6\]\[11\] RF.registers\[7\]\[11\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2189_ sky130_fd_sc_hd__mux4_1
X_8152_ RF.registers\[24\]\[21\] _3500_ _4047_ VGND VGND VPWR VPWR _4049_ sky130_fd_sc_hd__mux2_1
X_5364_ RF.registers\[0\]\[15\] RF.registers\[1\]\[15\] RF.registers\[2\]\[15\] RF.registers\[3\]\[15\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4315_ _1037_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__clkbuf_8
X_7103_ _3486_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_8083_ _4012_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__clkbuf_1
X_5295_ _2050_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__buf_4
X_7034_ RF.registers\[3\]\[24\] _3143_ _3435_ VGND VGND VPWR VPWR _3440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8985_ clknet_leaf_26_CLK _0145_ VGND VGND VPWR VPWR RF.registers\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7936_ RF.registers\[18\]\[16\] _3489_ _3927_ VGND VGND VPWR VPWR _3934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7867_ _3897_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__clkbuf_1
X_6818_ RF.registers\[6\]\[19\] _3132_ _3315_ VGND VGND VPWR VPWR _3325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7798_ RF.registers\[9\]\[15\] _3487_ _3855_ VGND VGND VPWR VPWR _3861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6749_ _3062_ RF.registers\[14\]\[19\] _3278_ VGND VGND VPWR VPWR _3288_ sky130_fd_sc_hd__mux2_1
X_9537_ clknet_leaf_95_CLK _0697_ VGND VGND VPWR VPWR RF.registers\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9468_ clknet_leaf_16_CLK _0628_ VGND VGND VPWR VPWR RF.registers\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8419_ RF.registers\[12\]\[19\] _3495_ _4180_ VGND VGND VPWR VPWR _4190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9399_ clknet_leaf_31_CLK _0559_ VGND VGND VPWR VPWR RF.registers\[24\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_3_1__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_70_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5080_ _1834_ _1835_ _1686_ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5982_ _1495_ _2657_ _2536_ VGND VGND VPWR VPWR _2723_ sky130_fd_sc_hd__a21oi_1
X_8770_ clknet_leaf_91_CLK _0954_ VGND VGND VPWR VPWR RF.registers\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_4933_ _1675_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7721_ _3820_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 _3141_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4864_ RF.registers\[16\]\[18\] RF.registers\[17\]\[18\] RF.registers\[18\]\[18\]
+ RF.registers\[19\]\[18\] _1200_ _1202_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7652_ RF.registers\[2\]\[10\] _3476_ _3783_ VGND VGND VPWR VPWR _3784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7583_ _3735_ VGND VGND VPWR VPWR _3747_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4795_ RF.registers\[12\]\[10\] RF.registers\[13\]\[10\] RF.registers\[14\]\[10\]
+ RF.registers\[15\]\[10\] _1052_ _1090_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__mux4_1
X_6603_ _3052_ RF.registers\[15\]\[14\] _3206_ VGND VGND VPWR VPWR _3211_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6534_ _3173_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9322_ clknet_leaf_9_CLK _0482_ VGND VGND VPWR VPWR RF.registers\[21\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6465_ net24 VGND VGND VPWR VPWR _3132_ sky130_fd_sc_hd__buf_2
X_9253_ clknet_leaf_59_CLK _0413_ VGND VGND VPWR VPWR RF.registers\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8204_ _4076_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__clkbuf_1
X_5416_ RF.registers\[0\]\[12\] RF.registers\[1\]\[12\] RF.registers\[2\]\[12\] RF.registers\[3\]\[12\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6396_ _3084_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9184_ clknet_leaf_70_CLK _0344_ VGND VGND VPWR VPWR RF.registers\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_5347_ _1127_ _1663_ _2100_ _2102_ VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__a31o_1
X_8135_ RF.registers\[24\]\[13\] _3483_ _4036_ VGND VGND VPWR VPWR _4040_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5278_ _1639_ _2033_ VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8066_ _4003_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__clkbuf_1
X_7017_ RF.registers\[3\]\[16\] _3126_ _3424_ VGND VGND VPWR VPWR _3431_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8968_ clknet_leaf_96_CLK _0128_ VGND VGND VPWR VPWR RF.registers\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7919_ RF.registers\[18\]\[8\] _3472_ _3916_ VGND VGND VPWR VPWR _3925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8899_ clknet_leaf_76_CLK _0059_ VGND VGND VPWR VPWR RF.registers\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4580_ RF.registers\[28\]\[30\] RF.registers\[29\]\[30\] RF.registers\[30\]\[30\]
+ RF.registers\[31\]\[30\] _1201_ _1203_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__mux4_1
Xinput11 A3[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 WD3[17] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
Xinput33 WD3[27] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput44 WD3[8] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6250_ _2178_ _1980_ _1960_ _1127_ VGND VGND VPWR VPWR _2976_ sky130_fd_sc_hd__o31a_1
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5201_ _1951_ _1953_ _1956_ _1773_ _1672_ VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__o221a_1
X_6181_ _2254_ _2848_ _2910_ _2336_ VGND VGND VPWR VPWR _2911_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5132_ RF.registers\[20\]\[31\] RF.registers\[21\]\[31\] RF.registers\[22\]\[31\]
+ RF.registers\[23\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__mux4_1
X_5063_ _1717_ _1818_ _1729_ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8822_ clknet_leaf_47_CLK _1006_ VGND VGND VPWR VPWR RF.registers\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_125_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8753_ clknet_leaf_13_CLK _0937_ VGND VGND VPWR VPWR RF.registers\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5965_ _1087_ _2706_ VGND VGND VPWR VPWR _2707_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4916_ _1671_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__clkbuf_4
X_5896_ _2595_ _2639_ _1572_ VGND VGND VPWR VPWR _2641_ sky130_fd_sc_hd__a21o_1
X_7704_ _3811_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8684_ clknet_leaf_9_CLK _0868_ VGND VGND VPWR VPWR RF.registers\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4847_ RF.registers\[20\]\[19\] RF.registers\[21\]\[19\] RF.registers\[22\]\[19\]
+ RF.registers\[23\]\[19\] _1182_ _1184_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7635_ RF.registers\[2\]\[2\] _3460_ _3772_ VGND VGND VPWR VPWR _3775_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9305_ clknet_leaf_27_CLK _0465_ VGND VGND VPWR VPWR RF.registers\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7566_ _3738_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
X_4778_ RF.registers\[8\]\[9\] RF.registers\[9\]\[9\] RF.registers\[10\]\[9\] RF.registers\[11\]\[9\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__mux4_1
X_7497_ _3025_ RF.registers\[27\]\[1\] _3700_ VGND VGND VPWR VPWR _3702_ sky130_fd_sc_hd__mux2_1
X_6517_ _3164_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__clkbuf_1
X_9236_ clknet_leaf_43_CLK _0396_ VGND VGND VPWR VPWR RF.registers\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_6448_ RF.registers\[17\]\[13\] _3120_ _3114_ VGND VGND VPWR VPWR _3121_ sky130_fd_sc_hd__mux2_1
X_6379_ net30 VGND VGND VPWR VPWR _3073_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9167_ clknet_leaf_13_CLK _0327_ VGND VGND VPWR VPWR RF.registers\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8118_ RF.registers\[24\]\[5\] _3466_ _4025_ VGND VGND VPWR VPWR _4031_ sky130_fd_sc_hd__mux2_1
X_9098_ clknet_leaf_8_CLK _0258_ VGND VGND VPWR VPWR RF.registers\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_8049_ _3994_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5750_ _2497_ _2500_ _2501_ VGND VGND VPWR VPWR _2502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5681_ _2255_ _2431_ _2434_ _2373_ VGND VGND VPWR VPWR _2435_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4701_ _1198_ _1456_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__or2_1
X_7420_ _3660_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4632_ RF.registers\[16\]\[6\] RF.registers\[17\]\[6\] RF.registers\[18\]\[6\] RF.registers\[19\]\[6\]
+ _1219_ _1221_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7351_ _3623_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4563_ _1317_ _1318_ _1198_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7282_ _3083_ RF.registers\[29\]\[29\] _3577_ VGND VGND VPWR VPWR _3587_ sky130_fd_sc_hd__mux2_1
X_4494_ _1199_ _1249_ _1213_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__o21a_1
X_6302_ net9 _3004_ VGND VGND VPWR VPWR _3020_ sky130_fd_sc_hd__nor2_4
XFILLER_0_40_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6233_ _1148_ _2958_ _2959_ _2337_ VGND VGND VPWR VPWR _2960_ sky130_fd_sc_hd__a211o_1
X_9021_ clknet_leaf_22_CLK _0181_ VGND VGND VPWR VPWR RF.registers\[31\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6164_ _2386_ _2391_ VGND VGND VPWR VPWR _2895_ sky130_fd_sc_hd__nor2_1
X_6095_ _1779_ _2829_ VGND VGND VPWR VPWR _2830_ sky130_fd_sc_hd__xor2_1
X_5115_ RF.registers\[0\]\[16\] RF.registers\[1\]\[16\] RF.registers\[2\]\[16\] RF.registers\[3\]\[16\]
+ _1822_ _1823_ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5046_ _1781_ _1801_ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6997_ _3420_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
X_8805_ clknet_leaf_82_CLK _0989_ VGND VGND VPWR VPWR RF.registers\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5948_ _2661_ _2669_ _2689_ VGND VGND VPWR VPWR _2691_ sky130_fd_sc_hd__a21boi_1
X_8736_ clknet_leaf_73_CLK _0920_ VGND VGND VPWR VPWR RF.registers\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8667_ clknet_leaf_44_CLK _0851_ VGND VGND VPWR VPWR RF.registers\[0\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5879_ _2548_ _2624_ _2426_ VGND VGND VPWR VPWR _2625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8598_ clknet_leaf_48_CLK _0782_ VGND VGND VPWR VPWR RF.registers\[22\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7618_ _3765_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7549_ _3077_ RF.registers\[27\]\[26\] _3722_ VGND VGND VPWR VPWR _3729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9219_ clknet_leaf_77_CLK _0379_ VGND VGND VPWR VPWR RF.registers\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6920_ _3379_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6851_ RF.registers\[5\]\[2\] _3097_ _3340_ VGND VGND VPWR VPWR _3343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5802_ _2530_ _2550_ _2551_ _2373_ VGND VGND VPWR VPWR _2552_ sky130_fd_sc_hd__o211a_1
X_9570_ clknet_leaf_91_CLK _0730_ VGND VGND VPWR VPWR RF.registers\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8521_ _4243_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__clkbuf_1
X_6782_ _3306_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__clkbuf_1
X_5733_ _2459_ _2467_ _2477_ _2485_ _2408_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_33_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5664_ _2082_ _2099_ VGND VGND VPWR VPWR _2418_ sky130_fd_sc_hd__nand2_1
X_8452_ RF.registers\[11\]\[2\] net36 _4205_ VGND VGND VPWR VPWR _4208_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4615_ RF.registers\[24\]\[24\] RF.registers\[25\]\[24\] RF.registers\[26\]\[24\]
+ RF.registers\[27\]\[24\] _1360_ _1361_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__mux4_1
X_7403_ _3067_ RF.registers\[26\]\[21\] _3650_ VGND VGND VPWR VPWR _3652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5595_ _1668_ _2194_ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8383_ _4171_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__clkbuf_1
X_4546_ _1300_ _1301_ _1259_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__mux2_1
X_7334_ _3067_ RF.registers\[31\]\[21\] _3613_ VGND VGND VPWR VPWR _3615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4477_ RF.registers\[8\]\[28\] RF.registers\[9\]\[28\] RF.registers\[10\]\[28\] RF.registers\[11\]\[28\]
+ _1182_ _1184_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__mux4_1
X_7265_ _3578_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
X_7196_ RF.registers\[7\]\[21\] _3500_ _3539_ VGND VGND VPWR VPWR _3541_ sky130_fd_sc_hd__mux2_1
X_6216_ _1980_ _1960_ VGND VGND VPWR VPWR _2944_ sky130_fd_sc_hd__nor2_1
X_9004_ clknet_leaf_2_CLK _0164_ VGND VGND VPWR VPWR RF.registers\[31\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6147_ _2814_ _2815_ _2748_ _2816_ _2878_ VGND VGND VPWR VPWR _2879_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_107_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _2813_ _2665_ _2745_ _2600_ VGND VGND VPWR VPWR _2814_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_107_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5029_ _1783_ _1784_ _1739_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8719_ clknet_leaf_12_CLK _0903_ VGND VGND VPWR VPWR RF.registers\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4400_ _1154_ _1155_ _1107_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5380_ RF.registers\[4\]\[14\] RF.registers\[5\]\[14\] RF.registers\[6\]\[14\] RF.registers\[7\]\[14\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4331_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__buf_2
X_7050_ net37 VGND VGND VPWR VPWR _3450_ sky130_fd_sc_hd__buf_2
X_6001_ _2536_ VGND VGND VPWR VPWR _2741_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7952_ _3942_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__clkbuf_1
X_6903_ RF.registers\[5\]\[27\] _3009_ _3362_ VGND VGND VPWR VPWR _3370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7883_ _3141_ RF.registers\[23\]\[23\] _3902_ VGND VGND VPWR VPWR _3906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6834_ _3333_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6765_ _3296_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__clkbuf_1
X_9553_ clknet_leaf_13_CLK _0713_ VGND VGND VPWR VPWR RF.registers\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8504_ RF.registers\[11\]\[27\] net33 _4227_ VGND VGND VPWR VPWR _4235_ sky130_fd_sc_hd__mux2_1
X_5716_ _2387_ _2393_ _1146_ VGND VGND VPWR VPWR _2469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9484_ clknet_leaf_2_CLK _0644_ VGND VGND VPWR VPWR RF.registers\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8435_ _4198_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__clkbuf_1
X_6696_ RF.registers\[8\]\[26\] _3002_ _3253_ VGND VGND VPWR VPWR _3260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _1168_ _1821_ _2401_ VGND VGND VPWR VPWR _2402_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8366_ RF.registers\[16\]\[26\] _3442_ _4155_ VGND VGND VPWR VPWR _4162_ sky130_fd_sc_hd__mux2_1
X_5578_ _2331_ _2332_ _2333_ VGND VGND VPWR VPWR _2334_ sky130_fd_sc_hd__a21o_1
X_8297_ _4125_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__clkbuf_1
X_4529_ _1283_ _1284_ _1198_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__mux2_1
X_7317_ _3050_ RF.registers\[31\]\[13\] _3602_ VGND VGND VPWR VPWR _3606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7248_ _3569_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7179_ RF.registers\[7\]\[13\] _3483_ _3528_ VGND VGND VPWR VPWR _3532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 A3[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ _1512_ _1573_ _1635_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6550_ RF.registers\[0\]\[22\] _3139_ _3179_ VGND VGND VPWR VPWR _3182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5501_ RF.registers\[16\]\[6\] RF.registers\[17\]\[6\] RF.registers\[18\]\[6\] RF.registers\[19\]\[6\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6481_ net30 VGND VGND VPWR VPWR _3143_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_117_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8220_ RF.registers\[1\]\[21\] _3500_ _4083_ VGND VGND VPWR VPWR _4085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5432_ _1686_ _2185_ _2187_ _1699_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__o211a_1
X_8151_ _4048_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__clkbuf_1
X_5363_ RF.registers\[4\]\[15\] RF.registers\[5\]\[15\] RF.registers\[6\]\[15\] RF.registers\[7\]\[15\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4314_ _1064_ _1069_ _1037_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__mux2_1
X_7102_ RF.registers\[19\]\[14\] _3485_ _3477_ VGND VGND VPWR VPWR _3486_ sky130_fd_sc_hd__mux2_1
X_8082_ RF.registers\[20\]\[20\] _3497_ _4011_ VGND VGND VPWR VPWR _4012_ sky130_fd_sc_hd__mux2_1
X_5294_ _1673_ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__buf_4
X_7033_ _3439_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8984_ clknet_leaf_38_CLK _0144_ VGND VGND VPWR VPWR RF.registers\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7935_ _3933_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7866_ _3124_ RF.registers\[23\]\[15\] _3891_ VGND VGND VPWR VPWR _3897_ sky130_fd_sc_hd__mux2_1
X_6817_ _3324_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__clkbuf_1
X_7797_ _3860_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__clkbuf_1
X_9536_ clknet_leaf_72_CLK _0696_ VGND VGND VPWR VPWR RF.registers\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6748_ _3287_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9467_ clknet_leaf_45_CLK _0627_ VGND VGND VPWR VPWR RF.registers\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6679_ RF.registers\[8\]\[18\] _3130_ _3242_ VGND VGND VPWR VPWR _3251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9398_ clknet_leaf_48_CLK _0558_ VGND VGND VPWR VPWR RF.registers\[24\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8418_ _4189_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8349_ RF.registers\[16\]\[18\] _3493_ _4144_ VGND VGND VPWR VPWR _4153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5981_ _2571_ _2605_ _2720_ _1087_ _2721_ VGND VGND VPWR VPWR _2722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4932_ RF.registers\[28\]\[23\] RF.registers\[29\]\[23\] RF.registers\[30\]\[23\]
+ RF.registers\[31\]\[23\] _1676_ _1681_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__mux4_1
X_7720_ _3043_ RF.registers\[30\]\[10\] _3819_ VGND VGND VPWR VPWR _3820_ sky130_fd_sc_hd__mux2_1
X_7651_ _3771_ VGND VGND VPWR VPWR _3783_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_14 _3491_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4863_ RF.registers\[20\]\[18\] RF.registers\[21\]\[18\] RF.registers\[22\]\[18\]
+ RF.registers\[23\]\[18\] _1200_ _1202_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6602_ _3210_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7582_ _3746_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4794_ RF.registers\[8\]\[10\] RF.registers\[9\]\[10\] RF.registers\[10\]\[10\] RF.registers\[11\]\[10\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_115_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6533_ RF.registers\[0\]\[14\] _3122_ _3168_ VGND VGND VPWR VPWR _3173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9321_ clknet_leaf_88_CLK _0481_ VGND VGND VPWR VPWR RF.registers\[21\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_99_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6464_ _3131_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9252_ clknet_leaf_94_CLK _0412_ VGND VGND VPWR VPWR RF.registers\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8203_ RF.registers\[1\]\[13\] _3483_ _4072_ VGND VGND VPWR VPWR _4076_ sky130_fd_sc_hd__mux2_1
X_5415_ RF.registers\[4\]\[12\] RF.registers\[5\]\[12\] RF.registers\[6\]\[12\] RF.registers\[7\]\[12\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2171_ sky130_fd_sc_hd__mux4_1
X_6395_ _3083_ RF.registers\[22\]\[29\] _3065_ VGND VGND VPWR VPWR _3084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9183_ clknet_leaf_72_CLK _0343_ VGND VGND VPWR VPWR RF.registers\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5346_ _1060_ _2101_ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__nand2_4
X_8134_ _4039_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5277_ _1777_ _2024_ _2032_ VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8065_ RF.registers\[20\]\[12\] _3481_ _4000_ VGND VGND VPWR VPWR _4003_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7016_ _3430_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8967_ clknet_leaf_58_CLK _0127_ VGND VGND VPWR VPWR RF.registers\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7918_ _3924_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8898_ clknet_leaf_92_CLK _0058_ VGND VGND VPWR VPWR RF.registers\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7849_ _3107_ RF.registers\[23\]\[7\] _3880_ VGND VGND VPWR VPWR _3888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9519_ clknet_leaf_11_CLK _0679_ VGND VGND VPWR VPWR RF.registers\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 A3[3] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput34 WD3[28] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_126_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput23 WD3[18] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput45 WD3[9] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5200_ _1954_ _1955_ _1889_ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__mux2_1
X_6180_ _2866_ _2909_ _2327_ VGND VGND VPWR VPWR _2910_ sky130_fd_sc_hd__mux2_1
X_5131_ RF.registers\[16\]\[31\] RF.registers\[17\]\[31\] RF.registers\[18\]\[31\]
+ RF.registers\[19\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5062_ _1816_ _1817_ _1686_ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8821_ clknet_leaf_53_CLK _1005_ VGND VGND VPWR VPWR RF.registers\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8752_ clknet_leaf_12_CLK _0936_ VGND VGND VPWR VPWR RF.registers\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5964_ _2549_ _2705_ _2104_ VGND VGND VPWR VPWR _2706_ sky130_fd_sc_hd__mux2_1
X_7703_ _3027_ RF.registers\[30\]\[2\] _3808_ VGND VGND VPWR VPWR _3811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5895_ _1572_ _2595_ _2639_ VGND VGND VPWR VPWR _2640_ sky130_fd_sc_hd__nand3_1
X_4915_ _1670_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_23_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8683_ clknet_leaf_86_CLK _0867_ VGND VGND VPWR VPWR RF.registers\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4846_ _1587_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7634_ _3774_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
X_7565_ _3025_ RF.registers\[28\]\[1\] _3736_ VGND VGND VPWR VPWR _3738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9304_ clknet_leaf_38_CLK _0464_ VGND VGND VPWR VPWR RF.registers\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4777_ _1529_ _1530_ _1531_ _1532_ _1040_ _1038_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__mux4_1
X_6516_ RF.registers\[0\]\[6\] _3105_ _3157_ VGND VGND VPWR VPWR _3164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7496_ _3701_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
X_9235_ clknet_leaf_36_CLK _0395_ VGND VGND VPWR VPWR RF.registers\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6447_ net18 VGND VGND VPWR VPWR _3120_ sky130_fd_sc_hd__buf_2
XFILLER_0_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6378_ _3072_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__clkbuf_1
X_9166_ clknet_leaf_39_CLK _0326_ VGND VGND VPWR VPWR RF.registers\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8117_ _4030_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__clkbuf_1
X_5329_ RF.registers\[28\]\[1\] RF.registers\[29\]\[1\] RF.registers\[30\]\[1\] RF.registers\[31\]\[1\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__mux4_1
X_9097_ clknet_leaf_1_CLK _0257_ VGND VGND VPWR VPWR RF.registers\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_8048_ RF.registers\[20\]\[4\] _3464_ _3989_ VGND VGND VPWR VPWR _3994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5680_ _1148_ _2432_ _2433_ _2337_ VGND VGND VPWR VPWR _2434_ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4700_ RF.registers\[4\]\[12\] RF.registers\[5\]\[12\] RF.registers\[6\]\[12\] RF.registers\[7\]\[12\]
+ _1172_ _1279_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4631_ RF.registers\[28\]\[6\] RF.registers\[29\]\[6\] RF.registers\[30\]\[6\] RF.registers\[31\]\[6\]
+ _1219_ _1221_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7350_ _3083_ RF.registers\[31\]\[29\] _3613_ VGND VGND VPWR VPWR _3623_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4562_ RF.registers\[16\]\[31\] RF.registers\[17\]\[31\] RF.registers\[18\]\[31\]
+ RF.registers\[19\]\[31\] _1200_ _1202_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__mux4_1
X_7281_ _3586_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
X_4493_ RF.registers\[12\]\[20\] RF.registers\[13\]\[20\] RF.registers\[14\]\[20\]
+ RF.registers\[15\]\[20\] _1201_ _1203_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6301_ net14 VGND VGND VPWR VPWR _3019_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9020_ clknet_leaf_23_CLK _0180_ VGND VGND VPWR VPWR RF.registers\[31\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6232_ _2923_ _2384_ _1148_ VGND VGND VPWR VPWR _2959_ sky130_fd_sc_hd__a21oi_1
X_6163_ _2887_ _2893_ VGND VGND VPWR VPWR _2894_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_127_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _1277_ _2828_ VGND VGND VPWR VPWR _2829_ sky130_fd_sc_hd__xnor2_1
X_5114_ RF.registers\[4\]\[16\] RF.registers\[5\]\[16\] RF.registers\[6\]\[16\] RF.registers\[7\]\[16\]
+ _1822_ _1823_ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5045_ _1758_ _1798_ _1800_ VGND VGND VPWR VPWR _1801_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8804_ clknet_leaf_78_CLK _0988_ VGND VGND VPWR VPWR RF.registers\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6996_ RF.registers\[3\]\[6\] _3105_ _3413_ VGND VGND VPWR VPWR _3420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5947_ _2689_ _2669_ _2661_ VGND VGND VPWR VPWR _2690_ sky130_fd_sc_hd__and3b_1
X_8735_ clknet_leaf_64_CLK _0919_ VGND VGND VPWR VPWR RF.registers\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8666_ clknet_leaf_46_CLK _0850_ VGND VGND VPWR VPWR RF.registers\[0\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7617_ _3077_ RF.registers\[28\]\[26\] _3758_ VGND VGND VPWR VPWR _3765_ sky130_fd_sc_hd__mux2_1
X_5878_ _2623_ VGND VGND VPWR VPWR _2624_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8597_ clknet_leaf_28_CLK _0781_ VGND VGND VPWR VPWR RF.registers\[22\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4829_ _1583_ _1584_ _1036_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7548_ _3728_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7479_ _3075_ RF.registers\[25\]\[25\] _3686_ VGND VGND VPWR VPWR _3692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9218_ clknet_leaf_91_CLK _0378_ VGND VGND VPWR VPWR RF.registers\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9149_ clknet_leaf_23_CLK _0309_ VGND VGND VPWR VPWR RF.registers\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6850_ _3342_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5801_ _2254_ _2425_ _2431_ _2337_ VGND VGND VPWR VPWR _2551_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6781_ RF.registers\[6\]\[1\] _3095_ _3304_ VGND VGND VPWR VPWR _3306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5732_ _2482_ _2484_ VGND VGND VPWR VPWR _2485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8520_ RF.registers\[10\]\[3\] net39 _3007_ VGND VGND VPWR VPWR _4243_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5663_ _1662_ VGND VGND VPWR VPWR _2417_ sky130_fd_sc_hd__inv_2
X_8451_ _4207_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4614_ _1171_ _1359_ _1365_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_115_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7402_ _3651_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
X_5594_ _1758_ _2175_ _1839_ VGND VGND VPWR VPWR _2349_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8382_ RF.registers\[12\]\[1\] _3458_ _4169_ VGND VGND VPWR VPWR _4171_ sky130_fd_sc_hd__mux2_1
X_4545_ RF.registers\[16\]\[27\] RF.registers\[17\]\[27\] RF.registers\[18\]\[27\]
+ RF.registers\[19\]\[27\] _1262_ _1263_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__mux4_1
X_7333_ _3614_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4476_ _1199_ _1231_ _1213_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__a21o_1
X_7264_ _3064_ RF.registers\[29\]\[20\] _3577_ VGND VGND VPWR VPWR _3578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9003_ clknet_leaf_0_CLK _0163_ VGND VGND VPWR VPWR RF.registers\[31\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7195_ _3540_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
X_6215_ _1962_ _2942_ _2421_ VGND VGND VPWR VPWR _2943_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6146_ _2808_ _2830_ _2840_ _2854_ VGND VGND VPWR VPWR _2878_ sky130_fd_sc_hd__or4_1
XFILLER_0_99_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _2601_ VGND VGND VPWR VPWR _2813_ sky130_fd_sc_hd__inv_2
X_5028_ RF.registers\[16\]\[20\] RF.registers\[17\]\[20\] RF.registers\[18\]\[20\]
+ RF.registers\[19\]\[20\] _1782_ _1680_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6979_ RF.registers\[4\]\[31\] _3017_ _3375_ VGND VGND VPWR VPWR _3410_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8718_ clknet_leaf_14_CLK _0902_ VGND VGND VPWR VPWR RF.registers\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8649_ clknet_leaf_86_CLK _0833_ VGND VGND VPWR VPWR RF.registers\[0\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4330_ _1060_ _1085_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6000_ _2584_ _2731_ _2736_ _2496_ _2739_ VGND VGND VPWR VPWR _2740_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7951_ RF.registers\[18\]\[23\] _3504_ _3938_ VGND VGND VPWR VPWR _3942_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7882_ _3905_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__clkbuf_1
X_6902_ _3369_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6833_ RF.registers\[6\]\[26\] _3002_ _3326_ VGND VGND VPWR VPWR _3333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6764_ _3077_ RF.registers\[14\]\[26\] _3289_ VGND VGND VPWR VPWR _3296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9552_ clknet_leaf_12_CLK _0712_ VGND VGND VPWR VPWR RF.registers\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6695_ _3259_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8503_ _4234_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__clkbuf_1
X_5715_ _1666_ VGND VGND VPWR VPWR _2468_ sky130_fd_sc_hd__inv_2
X_9483_ clknet_leaf_98_CLK _0643_ VGND VGND VPWR VPWR RF.registers\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8434_ RF.registers\[12\]\[26\] net32 _4191_ VGND VGND VPWR VPWR _4198_ sky130_fd_sc_hd__mux2_1
X_5646_ _1667_ _1859_ VGND VGND VPWR VPWR _2401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8365_ _4161_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__clkbuf_1
X_5577_ net48 VGND VGND VPWR VPWR _2333_ sky130_fd_sc_hd__buf_2
XFILLER_0_25_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8296_ _3145_ RF.registers\[13\]\[25\] _4119_ VGND VGND VPWR VPWR _4125_ sky130_fd_sc_hd__mux2_1
X_4528_ RF.registers\[24\]\[26\] RF.registers\[25\]\[26\] RF.registers\[26\]\[26\]
+ RF.registers\[27\]\[26\] _1181_ _1183_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__mux4_1
X_7316_ _3605_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
X_4459_ _1025_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7247_ _3048_ RF.registers\[29\]\[12\] _3566_ VGND VGND VPWR VPWR _3569_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7178_ _3531_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6129_ _2496_ _2859_ _2861_ _2504_ VGND VGND VPWR VPWR _2862_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_37_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_46_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5500_ RF.registers\[20\]\[6\] RF.registers\[21\]\[6\] RF.registers\[22\]\[6\] RF.registers\[23\]\[6\]
+ _1733_ _1679_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_117_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6480_ _3142_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5431_ _1711_ _2186_ VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8150_ RF.registers\[24\]\[20\] _3497_ _4047_ VGND VGND VPWR VPWR _4048_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_60_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_60_CLK sky130_fd_sc_hd__clkbuf_8
X_5362_ _1678_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_130_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8081_ _3988_ VGND VGND VPWR VPWR _4011_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4313_ _1067_ _1068_ _1035_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__mux2_1
X_7101_ net19 VGND VGND VPWR VPWR _3485_ sky130_fd_sc_hd__clkbuf_4
X_7032_ RF.registers\[3\]\[23\] _3141_ _3435_ VGND VGND VPWR VPWR _3439_ sky130_fd_sc_hd__mux2_1
X_5293_ _2045_ _2048_ _1696_ VGND VGND VPWR VPWR _2049_ sky130_fd_sc_hd__mux2_1
X_8983_ clknet_leaf_31_CLK _0143_ VGND VGND VPWR VPWR RF.registers\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7934_ RF.registers\[18\]\[15\] _3487_ _3927_ VGND VGND VPWR VPWR _3933_ sky130_fd_sc_hd__mux2_1
X_7865_ _3896_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__clkbuf_1
X_6816_ RF.registers\[6\]\[18\] _3130_ _3315_ VGND VGND VPWR VPWR _3324_ sky130_fd_sc_hd__mux2_1
X_7796_ RF.registers\[9\]\[14\] _3485_ _3855_ VGND VGND VPWR VPWR _3860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6747_ _3060_ RF.registers\[14\]\[18\] _3278_ VGND VGND VPWR VPWR _3287_ sky130_fd_sc_hd__mux2_1
X_9535_ clknet_leaf_64_CLK _0695_ VGND VGND VPWR VPWR RF.registers\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9466_ clknet_leaf_37_CLK _0626_ VGND VGND VPWR VPWR RF.registers\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6678_ _3250_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__clkbuf_1
X_9397_ clknet_leaf_28_CLK _0557_ VGND VGND VPWR VPWR RF.registers\[24\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5629_ _1799_ _1979_ VGND VGND VPWR VPWR _2384_ sky130_fd_sc_hd__nand2_1
X_8417_ RF.registers\[12\]\[18\] _3493_ _4180_ VGND VGND VPWR VPWR _4189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_51_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8348_ _4152_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8279_ _3128_ RF.registers\[13\]\[17\] _4108_ VGND VGND VPWR VPWR _4116_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_42_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5980_ _2468_ _2530_ _2426_ _2472_ _2503_ VGND VGND VPWR VPWR _2721_ sky130_fd_sc_hd__a41o_1
X_4931_ _1682_ _1683_ _1686_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4862_ _1239_ _1609_ _1617_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__o21ai_1
X_7650_ _3782_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6601_ _3050_ RF.registers\[15\]\[13\] _3206_ VGND VGND VPWR VPWR _3210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_15 _3650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7581_ _3041_ RF.registers\[28\]\[9\] _3736_ VGND VGND VPWR VPWR _3746_ sky130_fd_sc_hd__mux2_1
X_4793_ _1545_ _1548_ _1037_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__mux2_1
X_9320_ clknet_leaf_88_CLK _0480_ VGND VGND VPWR VPWR RF.registers\[21\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6532_ _3172_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6463_ RF.registers\[17\]\[18\] _3130_ _3114_ VGND VGND VPWR VPWR _3131_ sky130_fd_sc_hd__mux2_1
X_9251_ clknet_leaf_76_CLK _0411_ VGND VGND VPWR VPWR RF.registers\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9182_ clknet_leaf_69_CLK _0342_ VGND VGND VPWR VPWR RF.registers\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8202_ _4075_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__clkbuf_1
X_5414_ _1699_ _2169_ VGND VGND VPWR VPWR _2170_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_33_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_33_CLK sky130_fd_sc_hd__clkbuf_8
X_6394_ net35 VGND VGND VPWR VPWR _3083_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8133_ RF.registers\[24\]\[12\] _3481_ _4036_ VGND VGND VPWR VPWR _4039_ sky130_fd_sc_hd__mux2_1
X_5345_ _1664_ _1084_ VGND VGND VPWR VPWR _2101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5276_ _2026_ _2028_ _2031_ _1766_ _1672_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__o221a_1
X_8064_ _4002_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7015_ RF.registers\[3\]\[15\] _3124_ _3424_ VGND VGND VPWR VPWR _3430_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8966_ clknet_leaf_62_CLK _0126_ VGND VGND VPWR VPWR RF.registers\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7917_ RF.registers\[18\]\[7\] _3470_ _3916_ VGND VGND VPWR VPWR _3924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8897_ clknet_leaf_94_CLK _0057_ VGND VGND VPWR VPWR RF.registers\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7848_ _3887_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7779_ RF.registers\[9\]\[6\] _3468_ _3844_ VGND VGND VPWR VPWR _3851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9518_ clknet_leaf_11_CLK _0678_ VGND VGND VPWR VPWR RF.registers\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9449_ clknet_leaf_86_CLK _0609_ VGND VGND VPWR VPWR RF.registers\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_24_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 A3[4] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
Xinput35 WD3[29] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 WD3[19] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput46 WE3 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_15_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5130_ RF.registers\[28\]\[31\] RF.registers\[29\]\[31\] RF.registers\[30\]\[31\]
+ RF.registers\[31\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__mux4_1
X_5061_ RF.registers\[0\]\[18\] RF.registers\[1\]\[18\] RF.registers\[2\]\[18\] RF.registers\[3\]\[18\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8820_ clknet_leaf_53_CLK _1004_ VGND VGND VPWR VPWR RF.registers\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5963_ _2624_ _2704_ _2501_ VGND VGND VPWR VPWR _2705_ sky130_fd_sc_hd__mux2_1
X_8751_ clknet_leaf_11_CLK _0935_ VGND VGND VPWR VPWR RF.registers\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_7702_ _3810_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__clkbuf_1
X_4914_ _1640_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5894_ _2638_ _1416_ _2593_ _2594_ VGND VGND VPWR VPWR _2639_ sky130_fd_sc_hd__or4_1
X_8682_ clknet_leaf_87_CLK _0866_ VGND VGND VPWR VPWR RF.registers\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4845_ _1215_ _1592_ _1596_ _1600_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7633_ RF.registers\[2\]\[1\] _3458_ _3772_ VGND VGND VPWR VPWR _3774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4776_ RF.registers\[24\]\[9\] RF.registers\[25\]\[9\] RF.registers\[26\]\[9\] RF.registers\[27\]\[9\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__mux4_1
X_7564_ _3737_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9303_ clknet_leaf_32_CLK _0463_ VGND VGND VPWR VPWR RF.registers\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6515_ _3163_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__clkbuf_1
X_7495_ _3019_ RF.registers\[27\]\[0\] _3700_ VGND VGND VPWR VPWR _3701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9234_ clknet_leaf_41_CLK _0394_ VGND VGND VPWR VPWR RF.registers\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6446_ _3119_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6377_ _3071_ RF.registers\[22\]\[23\] _3065_ VGND VGND VPWR VPWR _3072_ sky130_fd_sc_hd__mux2_1
X_9165_ clknet_leaf_83_CLK _0325_ VGND VGND VPWR VPWR RF.registers\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8116_ RF.registers\[24\]\[4\] _3464_ _4025_ VGND VGND VPWR VPWR _4030_ sky130_fd_sc_hd__mux2_1
X_5328_ RF.registers\[24\]\[1\] RF.registers\[25\]\[1\] RF.registers\[26\]\[1\] RF.registers\[27\]\[1\]
+ _1673_ _1690_ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__mux4_1
X_9096_ clknet_leaf_0_CLK _0256_ VGND VGND VPWR VPWR RF.registers\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8047_ _3993_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__clkbuf_1
X_5259_ _1777_ _2006_ _2010_ _2014_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_3_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8949_ clknet_leaf_44_CLK _0109_ VGND VGND VPWR VPWR RF.registers\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_4_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_634 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4630_ RF.registers\[24\]\[6\] RF.registers\[25\]\[6\] RF.registers\[26\]\[6\] RF.registers\[27\]\[6\]
+ _1219_ _1221_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4561_ RF.registers\[20\]\[31\] RF.registers\[21\]\[31\] RF.registers\[22\]\[31\]
+ RF.registers\[23\]\[31\] _1200_ _1202_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__mux4_1
XFILLER_0_80_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6300_ _3018_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7280_ _3081_ RF.registers\[29\]\[28\] _3577_ VGND VGND VPWR VPWR _3586_ sky130_fd_sc_hd__mux2_1
X_4492_ _1190_ _1247_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6231_ _2380_ _2383_ VGND VGND VPWR VPWR _2958_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6162_ _2891_ _2892_ VGND VGND VPWR VPWR _2893_ sky130_fd_sc_hd__or2_1
X_5113_ _1717_ _1868_ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _1512_ _1256_ _1635_ _2658_ _2741_ VGND VGND VPWR VPWR _2828_ sky130_fd_sc_hd__a41o_1
X_5044_ _1799_ VGND VGND VPWR VPWR _1800_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8803_ clknet_leaf_73_CLK _0987_ VGND VGND VPWR VPWR RF.registers\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6995_ _3419_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5946_ _2687_ _2688_ VGND VGND VPWR VPWR _2689_ sky130_fd_sc_hd__or2_1
X_8734_ clknet_leaf_69_CLK _0918_ VGND VGND VPWR VPWR RF.registers\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8665_ clknet_3_7__leaf_CLK _0849_ VGND VGND VPWR VPWR RF.registers\[0\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5877_ _2581_ _2622_ _1146_ VGND VGND VPWR VPWR _2623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7616_ _3764_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
X_4828_ RF.registers\[0\]\[16\] RF.registers\[1\]\[16\] RF.registers\[2\]\[16\] RF.registers\[3\]\[16\]
+ _1181_ _1183_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8596_ clknet_leaf_17_CLK _0780_ VGND VGND VPWR VPWR RF.registers\[22\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7547_ _3075_ RF.registers\[27\]\[25\] _3722_ VGND VGND VPWR VPWR _3728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4759_ _1513_ _1514_ _1035_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__mux2_1
X_7478_ _3691_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9217_ clknet_leaf_95_CLK _0377_ VGND VGND VPWR VPWR RF.registers\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6429_ RF.registers\[17\]\[7\] _3107_ _3093_ VGND VGND VPWR VPWR _3108_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9148_ clknet_leaf_23_CLK _0308_ VGND VGND VPWR VPWR RF.registers\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_9079_ clknet_leaf_30_CLK _0239_ VGND VGND VPWR VPWR RF.registers\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_7__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_3_7__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5800_ _2439_ _2424_ _2501_ VGND VGND VPWR VPWR _2550_ sky130_fd_sc_hd__mux2_1
X_6780_ _3305_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5731_ _2449_ _2451_ _2483_ VGND VGND VPWR VPWR _2484_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5662_ _2376_ _2407_ _2408_ _2416_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__o2bb2a_1
X_8450_ RF.registers\[11\]\[1\] net25 _4205_ VGND VGND VPWR VPWR _4207_ sky130_fd_sc_hd__mux2_1
X_4613_ _1214_ _1368_ _1239_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_100_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7401_ _3064_ RF.registers\[26\]\[20\] _3650_ VGND VGND VPWR VPWR _3651_ sky130_fd_sc_hd__mux2_1
X_5593_ _2343_ _2346_ _2347_ VGND VGND VPWR VPWR _2348_ sky130_fd_sc_hd__mux2_1
X_8381_ _4170_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4544_ RF.registers\[20\]\[27\] RF.registers\[21\]\[27\] RF.registers\[22\]\[27\]
+ RF.registers\[23\]\[27\] _1262_ _1263_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7332_ _3064_ RF.registers\[31\]\[20\] _3613_ VGND VGND VPWR VPWR _3614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7263_ _3554_ VGND VGND VPWR VPWR _3577_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4475_ RF.registers\[0\]\[28\] RF.registers\[1\]\[28\] RF.registers\[2\]\[28\] RF.registers\[3\]\[28\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6214_ _2426_ _2591_ VGND VGND VPWR VPWR _2942_ sky130_fd_sc_hd__nand2_1
X_9002_ clknet_leaf_2_CLK _0162_ VGND VGND VPWR VPWR RF.registers\[31\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7194_ RF.registers\[7\]\[20\] _3497_ _3539_ VGND VGND VPWR VPWR _3540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6145_ _2875_ _2876_ VGND VGND VPWR VPWR _2877_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6076_ _2773_ _2809_ _2810_ _2811_ VGND VGND VPWR VPWR _2812_ sky130_fd_sc_hd__o211a_1
X_5027_ RF.registers\[20\]\[20\] RF.registers\[21\]\[20\] RF.registers\[22\]\[20\]
+ RF.registers\[23\]\[20\] _1782_ _1680_ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_107_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6978_ _3409_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
X_8717_ clknet_leaf_84_CLK _0901_ VGND VGND VPWR VPWR RF.registers\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5929_ _2547_ _2672_ _1147_ VGND VGND VPWR VPWR _2673_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8648_ clknet_leaf_79_CLK _0832_ VGND VGND VPWR VPWR RF.registers\[0\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8579_ clknet_leaf_76_CLK _0763_ VGND VGND VPWR VPWR RF.registers\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7950_ _3941_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__clkbuf_1
X_7881_ _3139_ RF.registers\[23\]\[22\] _3902_ VGND VGND VPWR VPWR _3905_ sky130_fd_sc_hd__mux2_1
X_6901_ RF.registers\[5\]\[26\] _3002_ _3362_ VGND VGND VPWR VPWR _3369_ sky130_fd_sc_hd__mux2_1
X_6832_ _3332_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6763_ _3295_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9551_ clknet_leaf_11_CLK _0711_ VGND VGND VPWR VPWR RF.registers\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6694_ RF.registers\[8\]\[25\] _3145_ _3253_ VGND VGND VPWR VPWR _3259_ sky130_fd_sc_hd__mux2_1
X_8502_ RF.registers\[11\]\[26\] net32 _4227_ VGND VGND VPWR VPWR _4234_ sky130_fd_sc_hd__mux2_1
X_5714_ _2105_ _2462_ _2466_ VGND VGND VPWR VPWR _2467_ sky130_fd_sc_hd__o21a_1
X_9482_ clknet_leaf_10_CLK _0642_ VGND VGND VPWR VPWR RF.registers\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8433_ _4197_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5645_ _2398_ _2399_ VGND VGND VPWR VPWR _2400_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8364_ RF.registers\[16\]\[25\] _3508_ _4155_ VGND VGND VPWR VPWR _4161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5576_ _1669_ _1660_ VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__nand2_1
X_8295_ _4124_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__clkbuf_1
X_4527_ RF.registers\[28\]\[26\] RF.registers\[29\]\[26\] RF.registers\[30\]\[26\]
+ RF.registers\[31\]\[26\] _1181_ _1183_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7315_ _3048_ RF.registers\[31\]\[12\] _3602_ VGND VGND VPWR VPWR _3605_ sky130_fd_sc_hd__mux2_1
X_4458_ _1213_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__clkbuf_4
X_7246_ _3568_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7177_ RF.registers\[7\]\[12\] _3481_ _3528_ VGND VGND VPWR VPWR _3531_ sky130_fd_sc_hd__mux2_1
X_6128_ _2373_ _2572_ _2823_ _2569_ _2860_ VGND VGND VPWR VPWR _2861_ sky130_fd_sc_hd__a221o_1
X_4389_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__clkbuf_4
X_6059_ _2102_ _2488_ VGND VGND VPWR VPWR _2795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5430_ RF.registers\[8\]\[11\] RF.registers\[9\]\[11\] RF.registers\[10\]\[11\] RF.registers\[11\]\[11\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5361_ _1702_ VGND VGND VPWR VPWR _2117_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_130_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8080_ _4010_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5292_ _2046_ _2047_ _2044_ VGND VGND VPWR VPWR _2048_ sky130_fd_sc_hd__mux2_1
X_4312_ RF.registers\[24\]\[5\] RF.registers\[25\]\[5\] RF.registers\[26\]\[5\] RF.registers\[27\]\[5\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__mux4_1
X_7100_ _3484_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
X_7031_ _3438_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8982_ clknet_leaf_32_CLK _0142_ VGND VGND VPWR VPWR RF.registers\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7933_ _3932_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7864_ _3122_ RF.registers\[23\]\[14\] _3891_ VGND VGND VPWR VPWR _3896_ sky130_fd_sc_hd__mux2_1
X_6815_ _3323_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7795_ _3859_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6746_ _3286_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__clkbuf_1
X_9534_ clknet_leaf_71_CLK _0694_ VGND VGND VPWR VPWR RF.registers\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9465_ clknet_leaf_32_CLK _0625_ VGND VGND VPWR VPWR RF.registers\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6677_ RF.registers\[8\]\[17\] _3128_ _3242_ VGND VGND VPWR VPWR _3250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9396_ clknet_leaf_23_CLK _0556_ VGND VGND VPWR VPWR RF.registers\[24\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_5628_ _1668_ _1959_ VGND VGND VPWR VPWR _2383_ sky130_fd_sc_hd__nand2_1
X_8416_ _4188_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8347_ RF.registers\[16\]\[17\] _3491_ _4144_ VGND VGND VPWR VPWR _4152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5559_ RF.registers\[8\]\[5\] RF.registers\[9\]\[5\] RF.registers\[10\]\[5\] RF.registers\[11\]\[5\]
+ _1718_ _1721_ VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8278_ _4115_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__clkbuf_1
X_7229_ _3559_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4930_ _1685_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4861_ _1611_ _1613_ _1616_ _1214_ _1170_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6600_ _3209_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4792_ _1546_ _1547_ _1034_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__mux2_1
X_7580_ _3745_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_16 _4133_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ RF.registers\[0\]\[13\] _3120_ _3168_ VGND VGND VPWR VPWR _3172_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6462_ net23 VGND VGND VPWR VPWR _3130_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9250_ clknet_leaf_92_CLK _0410_ VGND VGND VPWR VPWR RF.registers\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6393_ _3082_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__clkbuf_1
X_9181_ clknet_leaf_15_CLK _0341_ VGND VGND VPWR VPWR RF.registers\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_8201_ RF.registers\[1\]\[12\] _3481_ _4072_ VGND VGND VPWR VPWR _4075_ sky130_fd_sc_hd__mux2_1
X_5413_ _2167_ _2168_ _1711_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5344_ _2083_ _2099_ _1148_ VGND VGND VPWR VPWR _2100_ sky130_fd_sc_hd__mux2_1
X_8132_ _4038_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5275_ _2029_ _2030_ _1901_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__mux2_1
X_8063_ RF.registers\[20\]\[11\] _3479_ _4000_ VGND VGND VPWR VPWR _4002_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7014_ _3429_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8965_ clknet_leaf_64_CLK _0125_ VGND VGND VPWR VPWR RF.registers\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_8896_ clknet_leaf_70_CLK _0056_ VGND VGND VPWR VPWR RF.registers\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_7916_ _3923_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7847_ _3105_ RF.registers\[23\]\[6\] _3880_ VGND VGND VPWR VPWR _3887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7778_ _3850_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__clkbuf_1
X_9517_ clknet_leaf_10_CLK _0677_ VGND VGND VPWR VPWR RF.registers\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6729_ _3277_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9448_ clknet_leaf_88_CLK _0608_ VGND VGND VPWR VPWR RF.registers\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9379_ clknet_leaf_74_CLK _0539_ VGND VGND VPWR VPWR RF.registers\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput36 WD3[2] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
Xinput25 WD3[1] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 WD3[0] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XFILLER_0_25_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput47 opcode[0] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5060_ RF.registers\[4\]\[18\] RF.registers\[5\]\[18\] RF.registers\[6\]\[18\] RF.registers\[7\]\[18\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_125_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8750_ clknet_leaf_15_CLK _0934_ VGND VGND VPWR VPWR RF.registers\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_5962_ _2675_ _2703_ _2347_ VGND VGND VPWR VPWR _2704_ sky130_fd_sc_hd__mux2_1
X_4913_ _1668_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__clkbuf_4
X_7701_ _3025_ RF.registers\[30\]\[1\] _3808_ VGND VGND VPWR VPWR _3810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5893_ _1528_ _1542_ _1558_ VGND VGND VPWR VPWR _2638_ sky130_fd_sc_hd__nand3b_1
X_8681_ clknet_leaf_87_CLK _0865_ VGND VGND VPWR VPWR RF.registers\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4844_ _1205_ _1599_ _1057_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__a21oi_1
X_7632_ _3773_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
X_4775_ RF.registers\[28\]\[9\] RF.registers\[29\]\[9\] RF.registers\[30\]\[9\] RF.registers\[31\]\[9\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__mux4_1
X_7563_ _3019_ RF.registers\[28\]\[0\] _3736_ VGND VGND VPWR VPWR _3737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9302_ clknet_leaf_47_CLK _0462_ VGND VGND VPWR VPWR RF.registers\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6514_ RF.registers\[0\]\[5\] _3103_ _3157_ VGND VGND VPWR VPWR _3163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9233_ clknet_leaf_13_CLK _0393_ VGND VGND VPWR VPWR RF.registers\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_7494_ _3699_ VGND VGND VPWR VPWR _3700_ sky130_fd_sc_hd__buf_6
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6445_ RF.registers\[17\]\[12\] _3118_ _3114_ VGND VGND VPWR VPWR _3119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6376_ net29 VGND VGND VPWR VPWR _3071_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9164_ clknet_leaf_84_CLK _0324_ VGND VGND VPWR VPWR RF.registers\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5327_ _2064_ _2082_ VGND VGND VPWR VPWR _2083_ sky130_fd_sc_hd__and2_1
X_9095_ clknet_leaf_58_CLK _0255_ VGND VGND VPWR VPWR RF.registers\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8115_ _4029_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8046_ RF.registers\[20\]\[3\] _3462_ _3989_ VGND VGND VPWR VPWR _3993_ sky130_fd_sc_hd__mux2_1
X_5258_ _1766_ _2013_ _1672_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__o21ai_1
X_5189_ RF.registers\[24\]\[28\] RF.registers\[25\]\[28\] RF.registers\[26\]\[28\]
+ RF.registers\[27\]\[28\] _1882_ _1884_ VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_3_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8948_ clknet_leaf_44_CLK _0108_ VGND VGND VPWR VPWR RF.registers\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8879_ clknet_leaf_13_CLK _0039_ VGND VGND VPWR VPWR RF.registers\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4560_ _1299_ _1315_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4491_ RF.registers\[8\]\[20\] RF.registers\[9\]\[20\] RF.registers\[10\]\[20\] RF.registers\[11\]\[20\]
+ _1201_ _1203_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6230_ _2503_ _2955_ _2956_ VGND VGND VPWR VPWR _2957_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6161_ _2015_ _2889_ VGND VGND VPWR VPWR _2892_ sky130_fd_sc_hd__nor2_1
X_5112_ _1866_ _1867_ _1713_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6092_ _2812_ _2817_ _2808_ VGND VGND VPWR VPWR _2827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5043_ _1167_ VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8802_ clknet_leaf_77_CLK _0986_ VGND VGND VPWR VPWR RF.registers\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_6994_ RF.registers\[3\]\[5\] _3103_ _3413_ VGND VGND VPWR VPWR _3419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8733_ clknet_leaf_15_CLK _0917_ VGND VGND VPWR VPWR RF.registers\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5945_ _2684_ _2686_ _2160_ VGND VGND VPWR VPWR _2688_ sky130_fd_sc_hd__a21oi_1
X_8664_ clknet_leaf_40_CLK _0848_ VGND VGND VPWR VPWR RF.registers\[0\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_5876_ _1839_ _2211_ _2248_ VGND VGND VPWR VPWR _2622_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7615_ _3075_ RF.registers\[28\]\[25\] _3758_ VGND VGND VPWR VPWR _3764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4827_ RF.registers\[4\]\[16\] RF.registers\[5\]\[16\] RF.registers\[6\]\[16\] RF.registers\[7\]\[16\]
+ _1181_ _1183_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8595_ clknet_leaf_27_CLK _0779_ VGND VGND VPWR VPWR RF.registers\[22\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7546_ _3727_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4758_ RF.registers\[16\]\[8\] RF.registers\[17\]\[8\] RF.registers\[18\]\[8\] RF.registers\[19\]\[8\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__mux4_1
X_7477_ _3073_ RF.registers\[25\]\[24\] _3686_ VGND VGND VPWR VPWR _3691_ sky130_fd_sc_hd__mux2_1
X_4689_ _1439_ _1441_ _1444_ _1254_ _1170_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9216_ clknet_leaf_71_CLK _0376_ VGND VGND VPWR VPWR RF.registers\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6428_ net43 VGND VGND VPWR VPWR _3107_ sky130_fd_sc_hd__buf_2
X_9147_ clknet_leaf_46_CLK _0307_ VGND VGND VPWR VPWR RF.registers\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6359_ _3059_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9078_ clknet_leaf_33_CLK _0238_ VGND VGND VPWR VPWR RF.registers\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_8029_ _3011_ RF.registers\[21\]\[28\] _3974_ VGND VGND VPWR VPWR _3983_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5730_ _2080_ _2448_ VGND VGND VPWR VPWR _2483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7400_ _3627_ VGND VGND VPWR VPWR _3650_ sky130_fd_sc_hd__clkbuf_8
X_5661_ _2332_ _2415_ VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4612_ _1366_ _1367_ _1199_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5592_ _1146_ VGND VGND VPWR VPWR _2347_ sky130_fd_sc_hd__clkbuf_4
X_8380_ RF.registers\[12\]\[0\] _3454_ _4169_ VGND VGND VPWR VPWR _4170_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7331_ _3590_ VGND VGND VPWR VPWR _3613_ sky130_fd_sc_hd__clkbuf_8
X_4543_ _1298_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7262_ _3576_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4474_ _1189_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__and2_1
X_6213_ _2934_ _2940_ VGND VGND VPWR VPWR _2941_ sky130_fd_sc_hd__xor2_1
X_9001_ clknet_leaf_1_CLK _0161_ VGND VGND VPWR VPWR RF.registers\[31\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7193_ _3516_ VGND VGND VPWR VPWR _3539_ sky130_fd_sc_hd__buf_4
X_6144_ _2033_ _2874_ VGND VGND VPWR VPWR _2876_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6075_ _1838_ _2783_ VGND VGND VPWR VPWR _2811_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5026_ _1733_ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_107_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6977_ RF.registers\[4\]\[30\] _3015_ _3375_ VGND VGND VPWR VPWR _3409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5928_ _2428_ _2288_ VGND VGND VPWR VPWR _2672_ sky130_fd_sc_hd__nor2_1
X_8716_ clknet_leaf_11_CLK _0900_ VGND VGND VPWR VPWR RF.registers\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5859_ _2404_ _2605_ _2591_ _2356_ VGND VGND VPWR VPWR _2606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8647_ clknet_leaf_59_CLK _0831_ VGND VGND VPWR VPWR RF.registers\[0\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8578_ clknet_leaf_92_CLK _0762_ VGND VGND VPWR VPWR RF.registers\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7529_ _3718_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6900_ _3368_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__clkbuf_1
X_7880_ _3904_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6831_ RF.registers\[6\]\[25\] _3145_ _3326_ VGND VGND VPWR VPWR _3332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9550_ clknet_leaf_14_CLK _0710_ VGND VGND VPWR VPWR RF.registers\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6762_ _3075_ RF.registers\[14\]\[25\] _3289_ VGND VGND VPWR VPWR _3295_ sky130_fd_sc_hd__mux2_1
X_8501_ _4233_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6693_ _3258_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5713_ _2255_ _2463_ _2465_ _2373_ VGND VGND VPWR VPWR _2466_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9481_ clknet_leaf_87_CLK _0641_ VGND VGND VPWR VPWR RF.registers\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8432_ RF.registers\[12\]\[25\] _3508_ _4191_ VGND VGND VPWR VPWR _4197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5644_ _1842_ _1838_ _1799_ VGND VGND VPWR VPWR _2399_ sky130_fd_sc_hd__o21ai_1
X_8363_ _4160_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5575_ _1669_ _1660_ VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__or2_1
X_7314_ _3604_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
X_8294_ _3143_ RF.registers\[13\]\[24\] _4119_ VGND VGND VPWR VPWR _4124_ sky130_fd_sc_hd__mux2_1
X_4526_ _1280_ _1281_ _1198_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4457_ _1038_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__buf_4
X_7245_ _3046_ RF.registers\[29\]\[11\] _3566_ VGND VGND VPWR VPWR _3568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7176_ _3530_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_113_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _2719_ _2731_ VGND VGND VPWR VPWR _2860_ sky130_fd_sc_hd__and2_1
X_4388_ _1025_ _1135_ _1139_ _1143_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__a2bb2o_1
X_6058_ _2373_ _2476_ _2789_ _2794_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5009_ _1761_ _1764_ _1697_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5360_ _1685_ _2115_ _1696_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_130_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5291_ RF.registers\[24\]\[3\] RF.registers\[25\]\[3\] RF.registers\[26\]\[3\] RF.registers\[27\]\[3\]
+ _1674_ _1691_ VGND VGND VPWR VPWR _2047_ sky130_fd_sc_hd__mux4_1
X_4311_ RF.registers\[28\]\[5\] RF.registers\[29\]\[5\] RF.registers\[30\]\[5\] RF.registers\[31\]\[5\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7030_ RF.registers\[3\]\[22\] _3139_ _3435_ VGND VGND VPWR VPWR _3438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8981_ clknet_leaf_25_CLK _0141_ VGND VGND VPWR VPWR RF.registers\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7932_ RF.registers\[18\]\[14\] _3485_ _3927_ VGND VGND VPWR VPWR _3932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7863_ _3895_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6814_ RF.registers\[6\]\[17\] _3128_ _3315_ VGND VGND VPWR VPWR _3323_ sky130_fd_sc_hd__mux2_1
X_7794_ RF.registers\[9\]\[13\] _3483_ _3855_ VGND VGND VPWR VPWR _3859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9533_ clknet_leaf_15_CLK _0693_ VGND VGND VPWR VPWR RF.registers\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6745_ _3058_ RF.registers\[14\]\[17\] _3278_ VGND VGND VPWR VPWR _3286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9464_ clknet_leaf_38_CLK _0624_ VGND VGND VPWR VPWR RF.registers\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6676_ _3249_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__clkbuf_1
X_8415_ RF.registers\[12\]\[17\] _3491_ _4180_ VGND VGND VPWR VPWR _4188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9395_ clknet_leaf_27_CLK _0555_ VGND VGND VPWR VPWR RF.registers\[24\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5627_ _2378_ _2381_ _1877_ VGND VGND VPWR VPWR _2382_ sky130_fd_sc_hd__mux2_1
X_8346_ _4151_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5558_ _2310_ _2313_ net4 VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__mux2_1
X_4509_ _1261_ _1264_ _1259_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__mux2_1
X_8277_ _3126_ RF.registers\[13\]\[16\] _4108_ VGND VGND VPWR VPWR _4115_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5489_ _1697_ _2240_ _2242_ _2244_ _1729_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__a221o_1
X_7228_ _3029_ RF.registers\[29\]\[3\] _3555_ VGND VGND VPWR VPWR _3559_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7159_ _3521_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4860_ _1614_ _1615_ _1189_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_17 _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4791_ RF.registers\[24\]\[10\] RF.registers\[25\]\[10\] RF.registers\[26\]\[10\]
+ RF.registers\[27\]\[10\] _1041_ _1043_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__mux4_1
X_6530_ _3171_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_99_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6461_ _3129_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6392_ _3081_ RF.registers\[22\]\[28\] _3065_ VGND VGND VPWR VPWR _3082_ sky130_fd_sc_hd__mux2_1
X_9180_ clknet_leaf_37_CLK _0340_ VGND VGND VPWR VPWR RF.registers\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8200_ _4074_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__clkbuf_1
X_5412_ RF.registers\[12\]\[12\] RF.registers\[13\]\[12\] RF.registers\[14\]\[12\]
+ RF.registers\[15\]\[12\] _2117_ _2118_ VGND VGND VPWR VPWR _2168_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5343_ _1167_ _2098_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8131_ RF.registers\[24\]\[11\] _3479_ _4036_ VGND VGND VPWR VPWR _4038_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_120_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5274_ RF.registers\[0\]\[24\] RF.registers\[1\]\[24\] RF.registers\[2\]\[24\] RF.registers\[3\]\[24\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8062_ _4001_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7013_ RF.registers\[3\]\[14\] _3122_ _3424_ VGND VGND VPWR VPWR _3429_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8964_ clknet_leaf_96_CLK _0124_ VGND VGND VPWR VPWR RF.registers\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_7915_ RF.registers\[18\]\[6\] _3468_ _3916_ VGND VGND VPWR VPWR _3923_ sky130_fd_sc_hd__mux2_1
X_8895_ clknet_leaf_72_CLK _0055_ VGND VGND VPWR VPWR RF.registers\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7846_ _3886_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4989_ _1686_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7777_ RF.registers\[9\]\[5\] _3466_ _3844_ VGND VGND VPWR VPWR _3850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9516_ clknet_leaf_87_CLK _0676_ VGND VGND VPWR VPWR RF.registers\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6728_ _3041_ RF.registers\[14\]\[9\] _3267_ VGND VGND VPWR VPWR _3277_ sky130_fd_sc_hd__mux2_1
X_6659_ _3240_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9447_ clknet_leaf_81_CLK _0607_ VGND VGND VPWR VPWR RF.registers\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9378_ clknet_leaf_92_CLK _0538_ VGND VGND VPWR VPWR RF.registers\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8329_ _4142_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 WD3[20] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput37 WD3[30] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 WD3[10] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput48 opcode[1] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5961_ _2161_ _2142_ VGND VGND VPWR VPWR _2703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4912_ _1667_ VGND VGND VPWR VPWR _1668_ sky130_fd_sc_hd__buf_2
X_7700_ _3809_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__clkbuf_1
X_8680_ clknet_leaf_88_CLK _0864_ VGND VGND VPWR VPWR RF.registers\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5892_ _2627_ _2629_ _2637_ _2621_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__o22a_1
X_7631_ RF.registers\[2\]\[0\] _3454_ _3772_ VGND VGND VPWR VPWR _3773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4843_ _1597_ _1598_ _1036_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7562_ _3735_ VGND VGND VPWR VPWR _3736_ sky130_fd_sc_hd__buf_6
X_4774_ RF.registers\[16\]\[9\] RF.registers\[17\]\[9\] RF.registers\[18\]\[9\] RF.registers\[19\]\[9\]
+ _1072_ _1073_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__mux4_1
X_9301_ clknet_leaf_28_CLK _0461_ VGND VGND VPWR VPWR RF.registers\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_7493_ _3193_ _3626_ VGND VGND VPWR VPWR _3699_ sky130_fd_sc_hd__nand2_4
X_6513_ _3162_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9232_ clknet_leaf_84_CLK _0392_ VGND VGND VPWR VPWR RF.registers\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_6444_ net17 VGND VGND VPWR VPWR _3118_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6375_ _3070_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__clkbuf_1
X_9163_ clknet_leaf_90_CLK _0323_ VGND VGND VPWR VPWR RF.registers\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5326_ _1168_ _2081_ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_54_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8114_ RF.registers\[24\]\[3\] _3462_ _4025_ VGND VGND VPWR VPWR _4029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9094_ clknet_leaf_64_CLK _0254_ VGND VGND VPWR VPWR RF.registers\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_5257_ _2011_ _2012_ _1745_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__mux2_1
X_8045_ _3992_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__clkbuf_1
X_5188_ _1800_ _1943_ VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8947_ clknet_leaf_50_CLK _0107_ VGND VGND VPWR VPWR RF.registers\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8878_ clknet_leaf_56_CLK _0038_ VGND VGND VPWR VPWR RF.registers\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7829_ RF.registers\[9\]\[30\] _3450_ _3843_ VGND VGND VPWR VPWR _3877_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4490_ _1242_ _1245_ _1187_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6160_ _2890_ VGND VGND VPWR VPWR _2891_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5111_ RF.registers\[12\]\[16\] RF.registers\[13\]\[16\] RF.registers\[14\]\[16\]
+ RF.registers\[15\]\[16\] _1720_ _1723_ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_127_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _2528_ _2823_ _2731_ _2824_ _2825_ VGND VGND VPWR VPWR _2826_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5042_ _1729_ _1789_ _1797_ VGND VGND VPWR VPWR _1798_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8801_ clknet_leaf_72_CLK _0985_ VGND VGND VPWR VPWR RF.registers\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6993_ _3418_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
X_8732_ clknet_leaf_16_CLK _0916_ VGND VGND VPWR VPWR RF.registers\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_5944_ _2160_ _2684_ _2686_ VGND VGND VPWR VPWR _2687_ sky130_fd_sc_hd__and3_1
X_8663_ clknet_leaf_49_CLK _0847_ VGND VGND VPWR VPWR RF.registers\[0\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5875_ _2607_ _2614_ _2620_ _2621_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__o22a_1
X_7614_ _3763_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
X_8594_ clknet_leaf_40_CLK _0778_ VGND VGND VPWR VPWR RF.registers\[22\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_4826_ _1213_ _1581_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7545_ _3073_ RF.registers\[27\]\[24\] _3722_ VGND VGND VPWR VPWR _3727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4757_ RF.registers\[20\]\[8\] RF.registers\[21\]\[8\] RF.registers\[22\]\[8\] RF.registers\[23\]\[8\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__mux4_1
X_7476_ _3690_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
X_4688_ _1442_ _1443_ _1211_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6427_ _3106_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__clkbuf_1
X_9215_ clknet_leaf_65_CLK _0375_ VGND VGND VPWR VPWR RF.registers\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_9146_ clknet_leaf_24_CLK _0306_ VGND VGND VPWR VPWR RF.registers\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6358_ _3058_ RF.registers\[22\]\[17\] _3044_ VGND VGND VPWR VPWR _3059_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5309_ RF.registers\[20\]\[2\] RF.registers\[21\]\[2\] RF.registers\[22\]\[2\] RF.registers\[23\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__mux4_1
X_9077_ clknet_leaf_25_CLK _0237_ VGND VGND VPWR VPWR RF.registers\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6289_ net34 VGND VGND VPWR VPWR _3011_ sky130_fd_sc_hd__buf_2
X_8028_ _3982_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5660_ _2413_ _2414_ VGND VGND VPWR VPWR _2415_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4611_ RF.registers\[0\]\[25\] RF.registers\[1\]\[25\] RF.registers\[2\]\[25\] RF.registers\[3\]\[25\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5591_ _2344_ _2345_ VGND VGND VPWR VPWR _2346_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4542_ _1170_ _1286_ _1297_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__a21o_1
X_7330_ _3612_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_90_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_90_CLK sky130_fd_sc_hd__clkbuf_8
X_4473_ RF.registers\[4\]\[28\] RF.registers\[5\]\[28\] RF.registers\[6\]\[28\] RF.registers\[7\]\[28\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__mux4_1
X_7261_ _3062_ RF.registers\[29\]\[19\] _3566_ VGND VGND VPWR VPWR _3576_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6212_ _2885_ _2936_ _2939_ VGND VGND VPWR VPWR _2940_ sky130_fd_sc_hd__a21bo_1
X_9000_ clknet_leaf_0_CLK _0160_ VGND VGND VPWR VPWR RF.registers\[31\]\[10\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7192_ _3538_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_6143_ _2033_ _2874_ VGND VGND VPWR VPWR _2875_ sky130_fd_sc_hd__nor2_1
X_6074_ _1838_ _2783_ _2768_ _1820_ VGND VGND VPWR VPWR _2810_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5025_ _1168_ _1780_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_107_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6976_ _3408_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5927_ _2669_ _2670_ VGND VGND VPWR VPWR _2671_ sky130_fd_sc_hd__nand2_1
X_8715_ clknet_leaf_90_CLK _0899_ VGND VGND VPWR VPWR RF.registers\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5858_ _1111_ _2102_ VGND VGND VPWR VPWR _2605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8646_ clknet_leaf_61_CLK _0830_ VGND VGND VPWR VPWR RF.registers\[0\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5789_ _2271_ _2538_ VGND VGND VPWR VPWR _2539_ sky130_fd_sc_hd__and2_1
X_8577_ clknet_leaf_93_CLK _0761_ VGND VGND VPWR VPWR RF.registers\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4809_ RF.registers\[12\]\[11\] RF.registers\[13\]\[11\] RF.registers\[14\]\[11\]
+ RF.registers\[15\]\[11\] _1052_ _1053_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__mux4_1
X_7528_ _3056_ RF.registers\[27\]\[16\] _3711_ VGND VGND VPWR VPWR _3718_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_81_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_81_CLK sky130_fd_sc_hd__clkbuf_8
X_7459_ _3681_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9129_ clknet_leaf_1_CLK _0289_ VGND VGND VPWR VPWR RF.registers\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_72_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6830_ _3331_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6761_ _3294_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8500_ RF.registers\[11\]\[25\] net31 _4227_ VGND VGND VPWR VPWR _4233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5712_ _1148_ _2368_ _2369_ _2464_ _2336_ VGND VGND VPWR VPWR _2465_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6692_ RF.registers\[8\]\[24\] _3143_ _3253_ VGND VGND VPWR VPWR _3258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9480_ clknet_leaf_96_CLK _0640_ VGND VGND VPWR VPWR RF.registers\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8431_ _4196_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5643_ _1842_ _1798_ _1667_ VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8362_ RF.registers\[16\]\[24\] _3506_ _4155_ VGND VGND VPWR VPWR _4160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5574_ _1666_ _2041_ _2103_ _2329_ VGND VGND VPWR VPWR _2330_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_63_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_63_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4525_ RF.registers\[16\]\[26\] RF.registers\[17\]\[26\] RF.registers\[18\]\[26\]
+ RF.registers\[19\]\[26\] _1181_ _1183_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__mux4_1
X_7313_ _3046_ RF.registers\[31\]\[11\] _3602_ VGND VGND VPWR VPWR _3604_ sky130_fd_sc_hd__mux2_1
X_8293_ _4123_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__clkbuf_1
X_4456_ _1209_ _1210_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7244_ _3567_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4387_ _1088_ _1142_ net8 VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__a21oi_1
X_7175_ RF.registers\[7\]\[11\] _3479_ _3528_ VGND VGND VPWR VPWR _3530_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _2791_ _2858_ _2501_ VGND VGND VPWR VPWR _2859_ sky130_fd_sc_hd__mux2_1
X_6057_ _2651_ _2731_ _2792_ _2496_ _2793_ VGND VGND VPWR VPWR _2794_ sky130_fd_sc_hd__a221o_1
X_5008_ _1762_ _1763_ _1726_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6959_ RF.registers\[4\]\[21\] _3137_ _3398_ VGND VGND VPWR VPWR _3400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8629_ clknet_leaf_29_CLK _0813_ VGND VGND VPWR VPWR RF.registers\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_54_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_15_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_45_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5290_ RF.registers\[28\]\[3\] RF.registers\[29\]\[3\] RF.registers\[30\]\[3\] RF.registers\[31\]\[3\]
+ _1674_ _1691_ VGND VGND VPWR VPWR _2046_ sky130_fd_sc_hd__mux4_1
X_4310_ A2[1] VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8980_ clknet_leaf_23_CLK _0140_ VGND VGND VPWR VPWR RF.registers\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_42_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7931_ _3931_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7862_ _3120_ RF.registers\[23\]\[13\] _3891_ VGND VGND VPWR VPWR _3895_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6813_ _3322_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__clkbuf_1
X_7793_ _3858_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9532_ clknet_leaf_16_CLK _0692_ VGND VGND VPWR VPWR RF.registers\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6744_ _3285_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__clkbuf_1
X_9463_ clknet_leaf_49_CLK _0623_ VGND VGND VPWR VPWR RF.registers\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6675_ RF.registers\[8\]\[16\] _3126_ _3242_ VGND VGND VPWR VPWR _3249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5626_ _2379_ _2380_ VGND VGND VPWR VPWR _2381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8414_ _4187_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_51_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_36_CLK sky130_fd_sc_hd__clkbuf_8
X_9394_ clknet_leaf_41_CLK _0554_ VGND VGND VPWR VPWR RF.registers\[24\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8345_ RF.registers\[16\]\[16\] _3489_ _4144_ VGND VGND VPWR VPWR _4151_ sky130_fd_sc_hd__mux2_1
X_5557_ _2311_ _2312_ _1684_ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__mux2_1
X_4508_ RF.registers\[24\]\[21\] RF.registers\[25\]\[21\] RF.registers\[26\]\[21\]
+ RF.registers\[27\]\[21\] _1262_ _1263_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__mux4_1
X_8276_ _4114_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5488_ _1712_ _2243_ _1716_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4439_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__buf_4
X_7227_ _3558_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7158_ RF.registers\[7\]\[3\] _3462_ _3517_ VGND VGND VPWR VPWR _3521_ sky130_fd_sc_hd__mux2_1
X_6109_ _2806_ _2841_ _2842_ VGND VGND VPWR VPWR _2843_ sky130_fd_sc_hd__a21oi_1
X_7089_ _3455_ VGND VGND VPWR VPWR _3477_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_27_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4790_ RF.registers\[28\]\[10\] RF.registers\[29\]\[10\] RF.registers\[30\]\[10\]
+ RF.registers\[31\]\[10\] _1041_ _1043_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_18_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6460_ RF.registers\[17\]\[17\] _3128_ _3114_ VGND VGND VPWR VPWR _3129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6391_ net34 VGND VGND VPWR VPWR _3081_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_99_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5411_ RF.registers\[8\]\[12\] RF.registers\[9\]\[12\] RF.registers\[10\]\[12\] RF.registers\[11\]\[12\]
+ _2117_ _2118_ VGND VGND VPWR VPWR _2167_ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5342_ _1638_ _2097_ VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8130_ _4037_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8061_ RF.registers\[20\]\[10\] _3476_ _4000_ VGND VGND VPWR VPWR _4001_ sky130_fd_sc_hd__mux2_1
X_5273_ RF.registers\[4\]\[24\] RF.registers\[5\]\[24\] RF.registers\[6\]\[24\] RF.registers\[7\]\[24\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7012_ _3428_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8963_ clknet_leaf_74_CLK _0123_ VGND VGND VPWR VPWR RF.registers\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7914_ _3922_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__clkbuf_1
X_8894_ clknet_leaf_68_CLK _0054_ VGND VGND VPWR VPWR RF.registers\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7845_ _3103_ RF.registers\[23\]\[5\] _3880_ VGND VGND VPWR VPWR _3886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4988_ _1740_ _1743_ _1697_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__mux2_1
X_7776_ _3849_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9515_ clknet_leaf_90_CLK _0675_ VGND VGND VPWR VPWR RF.registers\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6727_ _3276_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6658_ RF.registers\[8\]\[8\] _3109_ _3231_ VGND VGND VPWR VPWR _3240_ sky130_fd_sc_hd__mux2_1
X_9446_ clknet_leaf_61_CLK _0606_ VGND VGND VPWR VPWR RF.registers\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5609_ _2359_ _2362_ _2363_ VGND VGND VPWR VPWR _2364_ sky130_fd_sc_hd__mux2_1
X_9377_ clknet_leaf_93_CLK _0537_ VGND VGND VPWR VPWR RF.registers\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6589_ _3203_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__clkbuf_1
X_8328_ RF.registers\[16\]\[8\] _3472_ _4133_ VGND VGND VPWR VPWR _4142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8259_ _4105_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput27 WD3[21] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput16 WD3[11] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 WD3[31] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_7_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_125_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5960_ _2421_ _2690_ _2691_ _2695_ _2702_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__o32a_1
X_5891_ _2633_ _2636_ VGND VGND VPWR VPWR _2637_ sky130_fd_sc_hd__xor2_1
X_4911_ _1171_ _1153_ _1157_ _1161_ _1165_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__a32oi_4
XTAP_TAPCELL_ROW_44_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7630_ _3771_ VGND VGND VPWR VPWR _3772_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4842_ RF.registers\[0\]\[17\] RF.registers\[1\]\[17\] RF.registers\[2\]\[17\] RF.registers\[3\]\[17\]
+ _1181_ _1183_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7561_ _3155_ _3553_ VGND VGND VPWR VPWR _3735_ sky130_fd_sc_hd__nand2b_4
X_4773_ RF.registers\[20\]\[9\] RF.registers\[21\]\[9\] RF.registers\[22\]\[9\] RF.registers\[23\]\[9\]
+ _1290_ _1193_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9300_ clknet_leaf_24_CLK _0460_ VGND VGND VPWR VPWR RF.registers\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7492_ _3698_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6512_ RF.registers\[0\]\[4\] _3101_ _3157_ VGND VGND VPWR VPWR _3162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9231_ clknet_leaf_11_CLK _0391_ VGND VGND VPWR VPWR RF.registers\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6443_ _3117_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6374_ _3069_ RF.registers\[22\]\[22\] _3065_ VGND VGND VPWR VPWR _3070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9162_ clknet_leaf_85_CLK _0322_ VGND VGND VPWR VPWR RF.registers\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_5325_ _1638_ _2080_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8113_ _4028_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__clkbuf_1
X_9093_ clknet_leaf_59_CLK _0253_ VGND VGND VPWR VPWR RF.registers\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5256_ RF.registers\[0\]\[25\] RF.registers\[1\]\[25\] RF.registers\[2\]\[25\] RF.registers\[3\]\[25\]
+ _1767_ _1768_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8044_ RF.registers\[20\]\[2\] _3460_ _3989_ VGND VGND VPWR VPWR _3992_ sky130_fd_sc_hd__mux2_1
X_5187_ _1638_ _1942_ VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_3_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8946_ clknet_leaf_54_CLK _0106_ VGND VGND VPWR VPWR RF.registers\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8877_ clknet_leaf_83_CLK _0037_ VGND VGND VPWR VPWR RF.registers\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7828_ _3876_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7759_ _3083_ RF.registers\[30\]\[29\] _3830_ VGND VGND VPWR VPWR _3840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9429_ clknet_leaf_51_CLK _0589_ VGND VGND VPWR VPWR RF.registers\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_692 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ _2102_ _2523_ VGND VGND VPWR VPWR _2825_ sky130_fd_sc_hd__nor2_1
X_5110_ RF.registers\[8\]\[16\] RF.registers\[9\]\[16\] RF.registers\[10\]\[16\] RF.registers\[11\]\[16\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5041_ _1791_ _1793_ _1796_ _1697_ _1671_ VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_0_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8800_ clknet_leaf_71_CLK _0984_ VGND VGND VPWR VPWR RF.registers\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8731_ clknet_leaf_50_CLK _0915_ VGND VGND VPWR VPWR RF.registers\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6992_ RF.registers\[3\]\[4\] _3101_ _3413_ VGND VGND VPWR VPWR _3418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5943_ _2536_ _2657_ _2685_ _2683_ VGND VGND VPWR VPWR _2686_ sky130_fd_sc_hd__o211ai_1
X_8662_ clknet_leaf_48_CLK _0846_ VGND VGND VPWR VPWR RF.registers\[0\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5874_ _2333_ VGND VGND VPWR VPWR _2621_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7613_ _3073_ RF.registers\[28\]\[24\] _3758_ VGND VGND VPWR VPWR _3763_ sky130_fd_sc_hd__mux2_1
X_8593_ clknet_leaf_20_CLK _0777_ VGND VGND VPWR VPWR RF.registers\[22\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_4825_ _1579_ _1580_ _1287_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7544_ _3726_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_138_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4756_ _1495_ _1511_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_60_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7475_ _3071_ RF.registers\[25\]\[23\] _3686_ VGND VGND VPWR VPWR _3690_ sky130_fd_sc_hd__mux2_1
X_4687_ RF.registers\[0\]\[22\] RF.registers\[1\]\[22\] RF.registers\[2\]\[22\] RF.registers\[3\]\[22\]
+ _1173_ _1175_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9214_ clknet_leaf_67_CLK _0374_ VGND VGND VPWR VPWR RF.registers\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6426_ RF.registers\[17\]\[6\] _3105_ _3093_ VGND VGND VPWR VPWR _3106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9145_ clknet_leaf_27_CLK _0305_ VGND VGND VPWR VPWR RF.registers\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6357_ net22 VGND VGND VPWR VPWR _3058_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_8_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5308_ _1167_ _2063_ VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__or2_1
X_6288_ _3010_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__clkbuf_1
X_9076_ clknet_leaf_23_CLK _0236_ VGND VGND VPWR VPWR RF.registers\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_8027_ _3009_ RF.registers\[21\]\[27\] _3974_ VGND VGND VPWR VPWR _3982_ sky130_fd_sc_hd__mux2_1
X_5239_ _1773_ _1990_ _1992_ _1994_ _1672_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_67_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8929_ clknet_leaf_79_CLK _0089_ VGND VGND VPWR VPWR RF.registers\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4610_ RF.registers\[4\]\[25\] RF.registers\[5\]\[25\] RF.registers\[6\]\[25\] RF.registers\[7\]\[25\]
+ _1360_ _1361_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5590_ _2144_ _2160_ _1668_ VGND VGND VPWR VPWR _2345_ sky130_fd_sc_hd__a21o_1
X_4541_ _1289_ _1293_ _1296_ _1205_ _1025_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4472_ _1224_ _1227_ _1187_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__mux2_1
X_7260_ _3575_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6211_ _2891_ _2937_ _2935_ _2938_ _2916_ VGND VGND VPWR VPWR _2939_ sky130_fd_sc_hd__o311a_1
X_7191_ RF.registers\[7\]\[19\] _3495_ _3528_ VGND VGND VPWR VPWR _3538_ sky130_fd_sc_hd__mux2_1
X_6142_ _1384_ _2873_ VGND VGND VPWR VPWR _2874_ sky130_fd_sc_hd__xnor2_1
X_6073_ _2769_ _2784_ VGND VGND VPWR VPWR _2809_ sky130_fd_sc_hd__or2_1
X_5024_ _1758_ _1779_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_107_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ RF.registers\[4\]\[29\] _3013_ _3398_ VGND VGND VPWR VPWR _3408_ sky130_fd_sc_hd__mux2_1
X_5926_ _2663_ _2668_ VGND VGND VPWR VPWR _2670_ sky130_fd_sc_hd__nand2_1
X_8714_ clknet_leaf_85_CLK _0898_ VGND VGND VPWR VPWR RF.registers\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8645_ clknet_leaf_80_CLK _0829_ VGND VGND VPWR VPWR RF.registers\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5857_ _2390_ _2590_ VGND VGND VPWR VPWR _2604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5788_ _1399_ _2537_ VGND VGND VPWR VPWR _2538_ sky130_fd_sc_hd__xnor2_1
X_8576_ clknet_leaf_74_CLK _0760_ VGND VGND VPWR VPWR RF.registers\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4808_ RF.registers\[8\]\[11\] RF.registers\[9\]\[11\] RF.registers\[10\]\[11\] RF.registers\[11\]\[11\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__mux4_1
X_4739_ _1464_ _1480_ _1494_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__and3_1
X_7527_ _3717_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7458_ _3054_ RF.registers\[25\]\[15\] _3675_ VGND VGND VPWR VPWR _3681_ sky130_fd_sc_hd__mux2_1
X_6409_ _3094_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7389_ _3644_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
X_9128_ clknet_leaf_96_CLK _0288_ VGND VGND VPWR VPWR RF.registers\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9059_ clknet_leaf_74_CLK _0219_ VGND VGND VPWR VPWR RF.registers\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_88_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6760_ _3073_ RF.registers\[14\]\[24\] _3289_ VGND VGND VPWR VPWR _3294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5711_ _2178_ _2362_ VGND VGND VPWR VPWR _2464_ sky130_fd_sc_hd__and2b_1
X_6691_ _3257_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8430_ RF.registers\[12\]\[24\] _3506_ _4191_ VGND VGND VPWR VPWR _4196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5642_ _2393_ _2396_ _1146_ VGND VGND VPWR VPWR _2397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8361_ _4159_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__clkbuf_1
X_5573_ _2105_ _2253_ _2255_ _2328_ VGND VGND VPWR VPWR _2329_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4524_ RF.registers\[20\]\[26\] RF.registers\[21\]\[26\] RF.registers\[22\]\[26\]
+ RF.registers\[23\]\[26\] _1172_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__mux4_1
X_7312_ _3603_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8292_ _3141_ RF.registers\[13\]\[23\] _4119_ VGND VGND VPWR VPWR _4123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4455_ _1198_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__buf_4
X_7243_ _3043_ RF.registers\[29\]\[10\] _3566_ VGND VGND VPWR VPWR _3567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4386_ _1140_ _1141_ _1107_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__mux2_1
X_7174_ _3529_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _2820_ _2857_ _1147_ VGND VGND VPWR VPWR _2858_ sky130_fd_sc_hd__mux2_1
X_6056_ _2458_ _2738_ VGND VGND VPWR VPWR _2793_ sky130_fd_sc_hd__nor2_1
X_5007_ RF.registers\[24\]\[21\] RF.registers\[25\]\[21\] RF.registers\[26\]\[21\]
+ RF.registers\[27\]\[21\] _1676_ _1681_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6958_ _3399_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6889_ RF.registers\[5\]\[20\] _3134_ _3362_ VGND VGND VPWR VPWR _3363_ sky130_fd_sc_hd__mux2_1
X_5909_ _2468_ _2530_ _2475_ _2503_ VGND VGND VPWR VPWR _2654_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8628_ clknet_leaf_24_CLK _0812_ VGND VGND VPWR VPWR RF.registers\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8559_ _4263_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7930_ RF.registers\[18\]\[13\] _3483_ _3927_ VGND VGND VPWR VPWR _3931_ sky130_fd_sc_hd__mux2_1
X_7861_ _3894_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6812_ RF.registers\[6\]\[16\] _3126_ _3315_ VGND VGND VPWR VPWR _3322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7792_ RF.registers\[9\]\[12\] _3481_ _3855_ VGND VGND VPWR VPWR _3858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9531_ clknet_leaf_45_CLK _0691_ VGND VGND VPWR VPWR RF.registers\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6743_ _3056_ RF.registers\[14\]\[16\] _3278_ VGND VGND VPWR VPWR _3285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9462_ clknet_leaf_33_CLK _0622_ VGND VGND VPWR VPWR RF.registers\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6674_ _3248_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5625_ _1167_ _1943_ VGND VGND VPWR VPWR _2380_ sky130_fd_sc_hd__and2_1
X_8413_ RF.registers\[12\]\[16\] _3489_ _4180_ VGND VGND VPWR VPWR _4187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9393_ clknet_leaf_15_CLK _0553_ VGND VGND VPWR VPWR RF.registers\[24\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8344_ _4150_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__clkbuf_1
X_5556_ RF.registers\[24\]\[5\] RF.registers\[25\]\[5\] RF.registers\[26\]\[5\] RF.registers\[27\]\[5\]
+ _1702_ _1678_ VGND VGND VPWR VPWR _2312_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8275_ _3124_ RF.registers\[13\]\[15\] _4108_ VGND VGND VPWR VPWR _4114_ sky130_fd_sc_hd__mux2_1
X_4507_ _1221_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5487_ RF.registers\[0\]\[9\] RF.registers\[1\]\[9\] RF.registers\[2\]\[9\] RF.registers\[3\]\[9\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_57_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7226_ _3027_ RF.registers\[29\]\[2\] _3555_ VGND VGND VPWR VPWR _3558_ sky130_fd_sc_hd__mux2_1
X_4438_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7157_ _3520_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_4369_ _1024_ _1116_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__o21ai_4
X_6108_ _1779_ _2829_ VGND VGND VPWR VPWR _2842_ sky130_fd_sc_hd__and2b_1
X_7088_ net15 VGND VGND VPWR VPWR _3476_ sky130_fd_sc_hd__buf_2
X_6039_ _1669_ _1821_ _1860_ VGND VGND VPWR VPWR _2777_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_19 _1416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6390_ _3080_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5410_ _2162_ _2163_ _2164_ _2165_ _1711_ _1716_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5341_ _1640_ _2088_ _2096_ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__o21ai_2
X_8060_ _3988_ VGND VGND VPWR VPWR _4000_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5272_ _1901_ _2027_ _1717_ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__a21o_1
X_7011_ RF.registers\[3\]\[13\] _3120_ _3424_ VGND VGND VPWR VPWR _3428_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8962_ clknet_leaf_93_CLK _0122_ VGND VGND VPWR VPWR RF.registers\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_7913_ RF.registers\[18\]\[5\] _3466_ _3916_ VGND VGND VPWR VPWR _3922_ sky130_fd_sc_hd__mux2_1
X_8893_ clknet_leaf_16_CLK _0053_ VGND VGND VPWR VPWR RF.registers\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7844_ _3885_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__clkbuf_1
X_7775_ RF.registers\[9\]\[4\] _3464_ _3844_ VGND VGND VPWR VPWR _3849_ sky130_fd_sc_hd__mux2_1
X_4987_ _1741_ _1742_ _1739_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9514_ clknet_leaf_85_CLK _0674_ VGND VGND VPWR VPWR RF.registers\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6726_ _3039_ RF.registers\[14\]\[8\] _3267_ VGND VGND VPWR VPWR _3276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9445_ clknet_leaf_80_CLK _0605_ VGND VGND VPWR VPWR RF.registers\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6657_ _3239_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__clkbuf_1
X_5608_ _1877_ VGND VGND VPWR VPWR _2363_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9376_ clknet_leaf_74_CLK _0536_ VGND VGND VPWR VPWR RF.registers\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6588_ _3037_ RF.registers\[15\]\[7\] _3195_ VGND VGND VPWR VPWR _3203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5539_ _2293_ _2294_ _2044_ VGND VGND VPWR VPWR _2295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8327_ _4141_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8258_ _3107_ RF.registers\[13\]\[7\] _4097_ VGND VGND VPWR VPWR _4105_ sky130_fd_sc_hd__mux2_1
X_7209_ _3547_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
X_8189_ _4068_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput28 WD3[22] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 WD3[12] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput39 WD3[3] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_1
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4910_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__buf_2
X_5890_ _2598_ _2618_ _2617_ _2635_ VGND VGND VPWR VPWR _2636_ sky130_fd_sc_hd__a31o_1
X_4841_ RF.registers\[4\]\[17\] RF.registers\[5\]\[17\] RF.registers\[6\]\[17\] RF.registers\[7\]\[17\]
+ _1181_ _1183_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7560_ _3734_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4772_ _1025_ _1519_ _1527_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__o21a_2
X_7491_ _3087_ RF.registers\[25\]\[31\] _3663_ VGND VGND VPWR VPWR _3698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6511_ _3161_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9230_ clknet_leaf_14_CLK _0390_ VGND VGND VPWR VPWR RF.registers\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_6442_ RF.registers\[17\]\[11\] _3116_ _3114_ VGND VGND VPWR VPWR _3117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9161_ clknet_leaf_86_CLK _0321_ VGND VGND VPWR VPWR RF.registers\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6373_ net28 VGND VGND VPWR VPWR _3069_ sky130_fd_sc_hd__buf_2
X_8112_ RF.registers\[24\]\[2\] _3460_ _4025_ VGND VGND VPWR VPWR _4028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9092_ clknet_leaf_96_CLK _0252_ VGND VGND VPWR VPWR RF.registers\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_5324_ net5 _2071_ _2079_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__a21oi_2
X_5255_ RF.registers\[4\]\[25\] RF.registers\[5\]\[25\] RF.registers\[6\]\[25\] RF.registers\[7\]\[25\]
+ _1895_ _1897_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8043_ _3991_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5186_ _1777_ _1933_ _1941_ VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8945_ clknet_leaf_56_CLK _0105_ VGND VGND VPWR VPWR RF.registers\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8876_ clknet_leaf_84_CLK _0036_ VGND VGND VPWR VPWR RF.registers\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_7827_ RF.registers\[9\]\[29\] _3448_ _3866_ VGND VGND VPWR VPWR _3876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7758_ _3839_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7689_ RF.registers\[2\]\[28\] _3446_ _3794_ VGND VGND VPWR VPWR _3803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6709_ _3266_ VGND VGND VPWR VPWR _3267_ sky130_fd_sc_hd__clkbuf_8
X_9428_ clknet_leaf_44_CLK _0588_ VGND VGND VPWR VPWR RF.registers\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9359_ clknet_leaf_5_CLK _0519_ VGND VGND VPWR VPWR RF.registers\[20\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_2__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_3_2__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _1794_ _1795_ _1739_ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6991_ _3417_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
X_8730_ clknet_leaf_35_CLK _0914_ VGND VGND VPWR VPWR RF.registers\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5942_ _1464_ _2411_ VGND VGND VPWR VPWR _2685_ sky130_fd_sc_hd__or2_1
X_8661_ clknet_leaf_51_CLK _0845_ VGND VGND VPWR VPWR RF.registers\[0\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_105_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5873_ _2617_ _2619_ VGND VGND VPWR VPWR _2620_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7612_ _3762_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
X_4824_ RF.registers\[12\]\[16\] RF.registers\[13\]\[16\] RF.registers\[14\]\[16\]
+ RF.registers\[15\]\[16\] _1191_ _1174_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__mux4_1
X_8592_ clknet_leaf_7_CLK _0776_ VGND VGND VPWR VPWR RF.registers\[22\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7543_ _3071_ RF.registers\[27\]\[23\] _3722_ VGND VGND VPWR VPWR _3726_ sky130_fd_sc_hd__mux2_1
X_4755_ _1239_ _1502_ _1506_ _1510_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_56_671 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7474_ _3689_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
X_4686_ RF.registers\[4\]\[22\] RF.registers\[5\]\[22\] RF.registers\[6\]\[22\] RF.registers\[7\]\[22\]
+ _1173_ _1175_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__mux4_1
X_9213_ clknet_leaf_22_CLK _0373_ VGND VGND VPWR VPWR RF.registers\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6425_ net42 VGND VGND VPWR VPWR _3105_ sky130_fd_sc_hd__buf_2
X_9144_ clknet_leaf_38_CLK _0304_ VGND VGND VPWR VPWR RF.registers\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6356_ _3057_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9075_ clknet_leaf_26_CLK _0235_ VGND VGND VPWR VPWR RF.registers\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5307_ _1638_ _2062_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6287_ RF.registers\[10\]\[27\] _3009_ _3007_ VGND VGND VPWR VPWR _3010_ sky130_fd_sc_hd__mux2_1
X_8026_ _3981_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_126_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5238_ _1901_ _1993_ _1766_ VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__a21o_1
X_5169_ _1169_ _1924_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8928_ clknet_leaf_73_CLK _0088_ VGND VGND VPWR VPWR RF.registers\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_8859_ clknet_leaf_44_CLK _0019_ VGND VGND VPWR VPWR RF.registers\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_135_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4540_ _1294_ _1295_ _1287_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4471_ _1225_ _1226_ _1178_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6210_ _1996_ _2903_ _2917_ VGND VGND VPWR VPWR _2938_ sky130_fd_sc_hd__or3b_1
X_7190_ _3537_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6141_ _2595_ _2872_ VGND VGND VPWR VPWR _2873_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6072_ _2806_ _2807_ VGND VGND VPWR VPWR _2808_ sky130_fd_sc_hd__or2_1
X_5023_ _1672_ _1765_ _1772_ _1778_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6974_ _3407_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5925_ _2663_ _2668_ VGND VGND VPWR VPWR _2669_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8713_ clknet_leaf_86_CLK _0897_ VGND VGND VPWR VPWR RF.registers\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5856_ _2587_ _2589_ _2592_ _2603_ _2408_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_62_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8644_ clknet_leaf_77_CLK _0828_ VGND VGND VPWR VPWR RF.registers\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4807_ _1559_ _1560_ _1561_ _1562_ _1048_ _1050_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__mux4_1
X_5787_ _2506_ _2535_ _2536_ VGND VGND VPWR VPWR _2537_ sky130_fd_sc_hd__a21oi_1
X_8575_ clknet_leaf_71_CLK _0759_ VGND VGND VPWR VPWR RF.registers\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7526_ _3054_ RF.registers\[27\]\[15\] _3711_ VGND VGND VPWR VPWR _3717_ sky130_fd_sc_hd__mux2_1
X_4738_ _1215_ _1485_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4669_ _1214_ _1424_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7457_ _3680_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6408_ RF.registers\[17\]\[0\] _3089_ _3093_ VGND VGND VPWR VPWR _3094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9127_ clknet_leaf_58_CLK _0287_ VGND VGND VPWR VPWR RF.registers\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_7388_ _3052_ RF.registers\[26\]\[14\] _3639_ VGND VGND VPWR VPWR _3644_ sky130_fd_sc_hd__mux2_1
X_6339_ net16 VGND VGND VPWR VPWR _3046_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_73_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9058_ clknet_leaf_92_CLK _0218_ VGND VGND VPWR VPWR RF.registers\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_8009_ _3972_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5710_ _2354_ _2359_ _2178_ VGND VGND VPWR VPWR _2463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6690_ RF.registers\[8\]\[23\] _3141_ _3253_ VGND VGND VPWR VPWR _3257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5641_ _2394_ _2395_ VGND VGND VPWR VPWR _2396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8360_ RF.registers\[16\]\[23\] _3504_ _4155_ VGND VGND VPWR VPWR _4159_ sky130_fd_sc_hd__mux2_1
X_5572_ _2289_ _2326_ _2327_ VGND VGND VPWR VPWR _2328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8291_ _4122_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7311_ _3043_ RF.registers\[31\]\[10\] _3602_ VGND VGND VPWR VPWR _3603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4523_ _1073_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__buf_4
X_7242_ _3554_ VGND VGND VPWR VPWR _3566_ sky130_fd_sc_hd__buf_4
X_4454_ RF.registers\[0\]\[29\] RF.registers\[1\]\[29\] RF.registers\[2\]\[29\] RF.registers\[3\]\[29\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4385_ RF.registers\[0\]\[1\] RF.registers\[1\]\[1\] RF.registers\[2\]\[1\] RF.registers\[3\]\[1\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__mux4_1
X_7173_ RF.registers\[7\]\[10\] _3476_ _3528_ VGND VGND VPWR VPWR _3529_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _2394_ _2392_ VGND VGND VPWR VPWR _2857_ sky130_fd_sc_hd__nor2_1
X_6055_ _2718_ _2791_ _2501_ VGND VGND VPWR VPWR _2792_ sky130_fd_sc_hd__mux2_1
X_5006_ RF.registers\[28\]\[21\] RF.registers\[29\]\[21\] RF.registers\[30\]\[21\]
+ RF.registers\[31\]\[21\] _1676_ _1681_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6957_ RF.registers\[4\]\[20\] _3134_ _3398_ VGND VGND VPWR VPWR _3399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6888_ _3339_ VGND VGND VPWR VPWR _3362_ sky130_fd_sc_hd__buf_4
X_5908_ _1087_ _2652_ VGND VGND VPWR VPWR _2653_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8627_ clknet_leaf_27_CLK _0811_ VGND VGND VPWR VPWR RF.registers\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5839_ _2335_ _2586_ VGND VGND VPWR VPWR _2587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8558_ RF.registers\[10\]\[21\] net27 _4255_ VGND VGND VPWR VPWR _4263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7509_ _3037_ RF.registers\[27\]\[7\] _3700_ VGND VGND VPWR VPWR _3708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8489_ _4204_ VGND VGND VPWR VPWR _4227_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_75_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7860_ _3118_ RF.registers\[23\]\[12\] _3891_ VGND VGND VPWR VPWR _3894_ sky130_fd_sc_hd__mux2_1
X_6811_ _3321_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7791_ _3857_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__clkbuf_1
X_9530_ clknet_leaf_35_CLK _0690_ VGND VGND VPWR VPWR RF.registers\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6742_ _3284_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9461_ clknet_leaf_36_CLK _0621_ VGND VGND VPWR VPWR RF.registers\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6673_ RF.registers\[8\]\[15\] _3124_ _3242_ VGND VGND VPWR VPWR _3248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5624_ _1799_ _1924_ VGND VGND VPWR VPWR _2379_ sky130_fd_sc_hd__nor2_1
X_9392_ clknet_leaf_7_CLK _0552_ VGND VGND VPWR VPWR RF.registers\[24\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8412_ _4186_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8343_ RF.registers\[16\]\[15\] _3487_ _4144_ VGND VGND VPWR VPWR _4150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5555_ RF.registers\[28\]\[5\] RF.registers\[29\]\[5\] RF.registers\[30\]\[5\] RF.registers\[31\]\[5\]
+ _2050_ _1678_ VGND VGND VPWR VPWR _2311_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4506_ _1219_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__clkbuf_8
X_5486_ _1739_ _2241_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8274_ _4113_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7225_ _3557_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_4437_ _1066_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__clkbuf_4
X_7156_ RF.registers\[7\]\[2\] _3460_ _3517_ VGND VGND VPWR VPWR _3520_ sky130_fd_sc_hd__mux2_1
X_6107_ _2829_ _1779_ VGND VGND VPWR VPWR _2841_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_70_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4368_ _1118_ _1120_ _1123_ _1037_ net8 VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a221o_1
X_7087_ _3475_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
X_4299_ RF.registers\[12\]\[4\] RF.registers\[13\]\[4\] RF.registers\[14\]\[4\] RF.registers\[15\]\[4\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__mux4_1
X_6038_ _2102_ _2445_ VGND VGND VPWR VPWR _2776_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7989_ _3111_ RF.registers\[21\]\[9\] _3952_ VGND VGND VPWR VPWR _3962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_636 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5340_ _2090_ _2092_ _2095_ net4 net5 VGND VGND VPWR VPWR _2096_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5271_ RF.registers\[8\]\[24\] RF.registers\[9\]\[24\] RF.registers\[10\]\[24\] RF.registers\[11\]\[24\]
+ _1881_ _1883_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__mux4_1
X_7010_ _3427_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8961_ clknet_leaf_97_CLK _0121_ VGND VGND VPWR VPWR RF.registers\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7912_ _3921_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__clkbuf_1
X_8892_ clknet_leaf_37_CLK _0052_ VGND VGND VPWR VPWR RF.registers\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7843_ _3101_ RF.registers\[23\]\[4\] _3880_ VGND VGND VPWR VPWR _3885_ sky130_fd_sc_hd__mux2_1
X_4986_ RF.registers\[24\]\[22\] RF.registers\[25\]\[22\] RF.registers\[26\]\[22\]
+ RF.registers\[27\]\[22\] _1734_ _1735_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7774_ _3848_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6725_ _3275_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__clkbuf_1
X_9513_ clknet_leaf_86_CLK _0673_ VGND VGND VPWR VPWR RF.registers\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9444_ clknet_leaf_89_CLK _0604_ VGND VGND VPWR VPWR RF.registers\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_6656_ RF.registers\[8\]\[7\] _3107_ _3231_ VGND VGND VPWR VPWR _3239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5607_ _2360_ _2361_ VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__and2_1
X_6587_ _3202_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__clkbuf_1
X_9375_ clknet_leaf_72_CLK _0535_ VGND VGND VPWR VPWR RF.registers\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5538_ RF.registers\[24\]\[4\] RF.registers\[25\]\[4\] RF.registers\[26\]\[4\] RF.registers\[27\]\[4\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2294_ sky130_fd_sc_hd__mux4_1
X_8326_ RF.registers\[16\]\[7\] _3470_ _4133_ VGND VGND VPWR VPWR _4141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8257_ _4104_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7208_ RF.registers\[7\]\[27\] _3444_ _3539_ VGND VGND VPWR VPWR _3547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5469_ RF.registers\[4\]\[8\] RF.registers\[5\]\[8\] RF.registers\[6\]\[8\] RF.registers\[7\]\[8\]
+ _1734_ _1735_ VGND VGND VPWR VPWR _2225_ sky130_fd_sc_hd__mux4_1
X_8188_ RF.registers\[1\]\[6\] _3468_ _4061_ VGND VGND VPWR VPWR _4068_ sky130_fd_sc_hd__mux2_1
X_7139_ _3510_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 WD3[13] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_37_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput29 WD3[23] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4840_ _1213_ _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6510_ RF.registers\[0\]\[3\] _3099_ _3157_ VGND VGND VPWR VPWR _3161_ sky130_fd_sc_hd__mux2_1
X_4771_ _1521_ _1523_ _1526_ _1050_ net8 VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__a221o_1
X_7490_ _3697_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6441_ net16 VGND VGND VPWR VPWR _3116_ sky130_fd_sc_hd__buf_2
XFILLER_0_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6372_ _3068_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9160_ clknet_leaf_78_CLK _0320_ VGND VGND VPWR VPWR RF.registers\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5323_ _2073_ _2075_ _2078_ net4 _1640_ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__o221a_1
X_8111_ _4027_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_54_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9091_ clknet_leaf_75_CLK _0251_ VGND VGND VPWR VPWR RF.registers\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5254_ _1773_ _2009_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__nor2_1
X_8042_ RF.registers\[20\]\[1\] _3458_ _3989_ VGND VGND VPWR VPWR _3991_ sky130_fd_sc_hd__mux2_1
X_5185_ _1935_ _1937_ _1940_ _1773_ _1671_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8944_ clknet_leaf_57_CLK _0104_ VGND VGND VPWR VPWR RF.registers\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_8875_ clknet_leaf_90_CLK _0035_ VGND VGND VPWR VPWR RF.registers\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7826_ _3875_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4969_ RF.registers\[0\]\[23\] RF.registers\[1\]\[23\] RF.registers\[2\]\[23\] RF.registers\[3\]\[23\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__mux4_1
X_7757_ _3081_ RF.registers\[30\]\[28\] _3830_ VGND VGND VPWR VPWR _3839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7688_ _3802_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6708_ _3020_ _3192_ VGND VGND VPWR VPWR _3266_ sky130_fd_sc_hd__nand2_4
X_9427_ clknet_leaf_50_CLK _0587_ VGND VGND VPWR VPWR RF.registers\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6639_ _3229_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9358_ clknet_leaf_20_CLK _0518_ VGND VGND VPWR VPWR RF.registers\[20\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_8309_ _4131_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__clkbuf_1
X_9289_ clknet_leaf_9_CLK _0449_ VGND VGND VPWR VPWR RF.registers\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6990_ RF.registers\[3\]\[3\] _3099_ _3413_ VGND VGND VPWR VPWR _3417_ sky130_fd_sc_hd__mux2_1
X_5941_ _1464_ _2657_ _2411_ _2683_ VGND VGND VPWR VPWR _2684_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8660_ clknet_leaf_53_CLK _0844_ VGND VGND VPWR VPWR RF.registers\[0\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5872_ _2229_ _2597_ _2598_ _2618_ VGND VGND VPWR VPWR _2619_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7611_ _3071_ RF.registers\[28\]\[23\] _3758_ VGND VGND VPWR VPWR _3762_ sky130_fd_sc_hd__mux2_1
X_4823_ RF.registers\[8\]\[16\] RF.registers\[9\]\[16\] RF.registers\[10\]\[16\] RF.registers\[11\]\[16\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__mux4_1
X_8591_ clknet_leaf_5_CLK _0775_ VGND VGND VPWR VPWR RF.registers\[22\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7542_ _3725_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
X_4754_ _1254_ _1509_ _1170_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_93_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_93_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7473_ _3069_ RF.registers\[25\]\[22\] _3686_ VGND VGND VPWR VPWR _3689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4685_ _1199_ _1440_ _1213_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__o21a_1
X_9212_ clknet_leaf_23_CLK _0372_ VGND VGND VPWR VPWR RF.registers\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6424_ _3104_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9143_ clknet_leaf_31_CLK _0303_ VGND VGND VPWR VPWR RF.registers\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_6355_ _3056_ RF.registers\[22\]\[16\] _3044_ VGND VGND VPWR VPWR _3057_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6286_ net33 VGND VGND VPWR VPWR _3009_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9074_ clknet_leaf_40_CLK _0234_ VGND VGND VPWR VPWR RF.registers\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5306_ _1729_ _2049_ _2057_ _2061_ VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__o2bb2a_2
X_8025_ _3002_ RF.registers\[21\]\[26\] _3974_ VGND VGND VPWR VPWR _3981_ sky130_fd_sc_hd__mux2_1
X_5237_ RF.registers\[0\]\[26\] RF.registers\[1\]\[26\] RF.registers\[2\]\[26\] RF.registers\[3\]\[26\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__mux4_1
X_5168_ _1639_ _1923_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5099_ RF.registers\[0\]\[17\] RF.registers\[1\]\[17\] RF.registers\[2\]\[17\] RF.registers\[3\]\[17\]
+ _1822_ _1823_ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_67_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8927_ clknet_leaf_65_CLK _0087_ VGND VGND VPWR VPWR RF.registers\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8858_ clknet_leaf_42_CLK _0018_ VGND VGND VPWR VPWR RF.registers\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8789_ clknet_leaf_44_CLK _0973_ VGND VGND VPWR VPWR RF.registers\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_7809_ RF.registers\[9\]\[20\] _3497_ _3866_ VGND VGND VPWR VPWR _3867_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_84_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_84_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_75_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_75_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_100_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4470_ RF.registers\[24\]\[28\] RF.registers\[25\]\[28\] RF.registers\[26\]\[28\]
+ RF.registers\[27\]\[28\] _1220_ _1222_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6140_ _1447_ _2871_ VGND VGND VPWR VPWR _2872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6071_ _1798_ _2805_ VGND VGND VPWR VPWR _2807_ sky130_fd_sc_hd__and2_1
X_5022_ _1773_ _1776_ _1777_ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6973_ RF.registers\[4\]\[28\] _3011_ _3398_ VGND VGND VPWR VPWR _3407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5924_ _2602_ _2665_ _2667_ VGND VGND VPWR VPWR _2668_ sky130_fd_sc_hd__o21a_1
X_8712_ clknet_leaf_89_CLK _0896_ VGND VGND VPWR VPWR RF.registers\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_5855_ _2598_ _2602_ VGND VGND VPWR VPWR _2603_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_62_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8643_ clknet_leaf_73_CLK _0827_ VGND VGND VPWR VPWR RF.registers\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4806_ RF.registers\[20\]\[11\] RF.registers\[21\]\[11\] RF.registers\[22\]\[11\]
+ RF.registers\[23\]\[11\] _1072_ _1073_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5786_ _2411_ VGND VGND VPWR VPWR _2536_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8574_ clknet_leaf_68_CLK _0758_ VGND VGND VPWR VPWR RF.registers\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_66_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_66_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_32_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4737_ _1487_ _1489_ _1492_ _1213_ _1057_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7525_ _3716_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
X_4668_ _1422_ _1423_ _1190_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7456_ _3052_ RF.registers\[25\]\[14\] _3675_ VGND VGND VPWR VPWR _3680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6407_ _3092_ VGND VGND VPWR VPWR _3093_ sky130_fd_sc_hd__buf_6
X_4599_ _1353_ _1354_ _1199_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7387_ _3643_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
X_9126_ clknet_leaf_66_CLK _0286_ VGND VGND VPWR VPWR RF.registers\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_6338_ _3045_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__clkbuf_1
X_6269_ _2992_ _2993_ VGND VGND VPWR VPWR _2994_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9057_ clknet_leaf_94_CLK _0217_ VGND VGND VPWR VPWR RF.registers\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8008_ _3130_ RF.registers\[21\]\[18\] _3963_ VGND VGND VPWR VPWR _3972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_57_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_57_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_48_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_48_CLK sky130_fd_sc_hd__clkbuf_8
X_5640_ _1668_ _1780_ VGND VGND VPWR VPWR _2395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5571_ _1803_ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8290_ _3139_ RF.registers\[13\]\[22\] _4119_ VGND VGND VPWR VPWR _4122_ sky130_fd_sc_hd__mux2_1
X_4522_ _1256_ _1277_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__nand2_1
X_7310_ _3590_ VGND VGND VPWR VPWR _3602_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4453_ RF.registers\[4\]\[29\] RF.registers\[5\]\[29\] RF.registers\[6\]\[29\] RF.registers\[7\]\[29\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__mux4_1
XFILLER_0_80_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7241_ _3565_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7172_ _3516_ VGND VGND VPWR VPWR _3528_ sky130_fd_sc_hd__buf_4
X_4384_ RF.registers\[4\]\[1\] RF.registers\[5\]\[1\] RF.registers\[6\]\[1\] RF.registers\[7\]\[1\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_113_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ _2854_ _2855_ VGND VGND VPWR VPWR _2856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6054_ _2752_ _2790_ _1147_ VGND VGND VPWR VPWR _2791_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5005_ _1759_ _1760_ _1726_ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6956_ _3375_ VGND VGND VPWR VPWR _3398_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_37_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5907_ _2458_ _2487_ _2651_ _2530_ VGND VGND VPWR VPWR _2652_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6887_ _3361_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8626_ clknet_leaf_43_CLK _0810_ VGND VGND VPWR VPWR RF.registers\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_39_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_39_CLK sky130_fd_sc_hd__clkbuf_8
X_5838_ _2105_ _2584_ _2487_ _2585_ VGND VGND VPWR VPWR _2586_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8557_ _4262_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__clkbuf_1
X_5769_ _2518_ _2519_ VGND VGND VPWR VPWR _2520_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7508_ _3707_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8488_ _4226_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7439_ _3035_ RF.registers\[25\]\[6\] _3664_ VGND VGND VPWR VPWR _3671_ sky130_fd_sc_hd__mux2_1
X_9109_ clknet_leaf_25_CLK _0269_ VGND VGND VPWR VPWR RF.registers\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6810_ RF.registers\[6\]\[15\] _3124_ _3315_ VGND VGND VPWR VPWR _3321_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_11_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7790_ RF.registers\[9\]\[11\] _3479_ _3855_ VGND VGND VPWR VPWR _3857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6741_ _3054_ RF.registers\[14\]\[15\] _3278_ VGND VGND VPWR VPWR _3284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9460_ clknet_leaf_43_CLK _0620_ VGND VGND VPWR VPWR RF.registers\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6672_ _3247_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5623_ _2377_ VGND VGND VPWR VPWR _2378_ sky130_fd_sc_hd__inv_2
X_9391_ clknet_leaf_4_CLK _0551_ VGND VGND VPWR VPWR RF.registers\[24\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8411_ RF.registers\[12\]\[15\] _3487_ _4180_ VGND VGND VPWR VPWR _4186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8342_ _4149_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5554_ _2308_ _2309_ _1684_ VGND VGND VPWR VPWR _2310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_667 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4505_ RF.registers\[28\]\[21\] RF.registers\[29\]\[21\] RF.registers\[30\]\[21\]
+ RF.registers\[31\]\[21\] _1220_ _1222_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5485_ RF.registers\[4\]\[9\] RF.registers\[5\]\[9\] RF.registers\[6\]\[9\] RF.registers\[7\]\[9\]
+ _1734_ _1735_ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__mux4_1
X_8273_ _3122_ RF.registers\[13\]\[14\] _4108_ VGND VGND VPWR VPWR _4113_ sky130_fd_sc_hd__mux2_1
X_4436_ _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_57_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7224_ _3025_ RF.registers\[29\]\[1\] _3555_ VGND VGND VPWR VPWR _3557_ sky130_fd_sc_hd__mux2_1
X_4367_ _1121_ _1122_ _1047_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__mux2_1
X_7155_ _3519_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
X_6106_ _2838_ _2839_ VGND VGND VPWR VPWR _2840_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_70_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7086_ RF.registers\[19\]\[9\] _3474_ _3456_ VGND VGND VPWR VPWR _3475_ sky130_fd_sc_hd__mux2_1
X_4298_ RF.registers\[8\]\[4\] RF.registers\[9\]\[4\] RF.registers\[10\]\[4\] RF.registers\[11\]\[4\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__mux4_1
X_6037_ _2769_ _2774_ VGND VGND VPWR VPWR _2775_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7988_ _3961_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6939_ _3389_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8609_ clknet_leaf_94_CLK _0793_ VGND VGND VPWR VPWR RF.registers\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_9589_ clknet_leaf_35_CLK _0749_ VGND VGND VPWR VPWR RF.registers\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5270_ _1889_ _2025_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8960_ clknet_leaf_69_CLK _0120_ VGND VGND VPWR VPWR RF.registers\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_7911_ RF.registers\[18\]\[4\] _3464_ _3916_ VGND VGND VPWR VPWR _3921_ sky130_fd_sc_hd__mux2_1
X_8891_ clknet_leaf_44_CLK _0051_ VGND VGND VPWR VPWR RF.registers\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7842_ _3884_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__clkbuf_1
X_4985_ RF.registers\[28\]\[22\] RF.registers\[29\]\[22\] RF.registers\[30\]\[22\]
+ RF.registers\[31\]\[22\] _1734_ _1735_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7773_ RF.registers\[9\]\[3\] _3462_ _3844_ VGND VGND VPWR VPWR _3848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9512_ clknet_leaf_87_CLK _0672_ VGND VGND VPWR VPWR RF.registers\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6724_ _3037_ RF.registers\[14\]\[7\] _3267_ VGND VGND VPWR VPWR _3275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9443_ clknet_leaf_75_CLK _0603_ VGND VGND VPWR VPWR RF.registers\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6655_ _3238_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5606_ _1667_ _2272_ VGND VGND VPWR VPWR _2361_ sky130_fd_sc_hd__nand2_1
X_9374_ clknet_leaf_69_CLK _0534_ VGND VGND VPWR VPWR RF.registers\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6586_ _3035_ RF.registers\[15\]\[6\] _3195_ VGND VGND VPWR VPWR _3202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5537_ RF.registers\[28\]\[4\] RF.registers\[29\]\[4\] RF.registers\[30\]\[4\] RF.registers\[31\]\[4\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2293_ sky130_fd_sc_hd__mux4_1
X_8325_ _4140_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8256_ _3105_ RF.registers\[13\]\[6\] _4097_ VGND VGND VPWR VPWR _4104_ sky130_fd_sc_hd__mux2_1
X_7207_ _3546_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_5468_ _1697_ _2223_ VGND VGND VPWR VPWR _2224_ sky130_fd_sc_hd__nand2_1
X_4419_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__buf_4
X_8187_ _4067_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5399_ _1711_ _2154_ _1655_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__o21a_1
X_7138_ RF.registers\[19\]\[26\] _3442_ _3498_ VGND VGND VPWR VPWR _3510_ sky130_fd_sc_hd__mux2_1
X_7069_ _3463_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 WD3[14] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_125_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4770_ _1524_ _1525_ _1035_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6440_ _3115_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6371_ _3067_ RF.registers\[22\]\[21\] _3065_ VGND VGND VPWR VPWR _3068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5322_ _2076_ _2077_ _1684_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8110_ RF.registers\[24\]\[1\] _3458_ _4025_ VGND VGND VPWR VPWR _4027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9090_ clknet_leaf_92_CLK _0250_ VGND VGND VPWR VPWR RF.registers\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5253_ _2007_ _2008_ _1713_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__mux2_1
X_8041_ _3990_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__clkbuf_1
X_5184_ _1938_ _1939_ _1713_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8943_ clknet_leaf_84_CLK _0103_ VGND VGND VPWR VPWR RF.registers\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_8874_ clknet_leaf_85_CLK _0034_ VGND VGND VPWR VPWR RF.registers\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_7825_ RF.registers\[9\]\[28\] _3446_ _3866_ VGND VGND VPWR VPWR _3875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7756_ _3838_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__clkbuf_1
X_4968_ RF.registers\[4\]\[23\] RF.registers\[5\]\[23\] RF.registers\[6\]\[23\] RF.registers\[7\]\[23\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7687_ RF.registers\[2\]\[27\] _3444_ _3794_ VGND VGND VPWR VPWR _3802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6707_ _3265_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4899_ net4 VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9426_ clknet_leaf_54_CLK _0586_ VGND VGND VPWR VPWR RF.registers\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_6638_ _3087_ RF.registers\[15\]\[31\] _3194_ VGND VGND VPWR VPWR _3229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9357_ clknet_leaf_8_CLK _0517_ VGND VGND VPWR VPWR RF.registers\[20\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6569_ _3191_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__clkbuf_1
X_8308_ _3017_ RF.registers\[13\]\[31\] _4096_ VGND VGND VPWR VPWR _4131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9288_ clknet_leaf_1_CLK _0448_ VGND VGND VPWR VPWR RF.registers\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_8239_ _4094_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5940_ _1480_ VGND VGND VPWR VPWR _2683_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7610_ _3761_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5871_ _2600_ _2601_ VGND VGND VPWR VPWR _2618_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8590_ clknet_leaf_21_CLK _0774_ VGND VGND VPWR VPWR RF.registers\[22\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_4822_ _1574_ _1575_ _1576_ _1577_ _1287_ _1078_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__mux4_2
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7541_ _3069_ RF.registers\[27\]\[22\] _3722_ VGND VGND VPWR VPWR _3725_ sky130_fd_sc_hd__mux2_1
X_4753_ _1507_ _1508_ _1211_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7472_ _3688_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9211_ clknet_leaf_34_CLK _0371_ VGND VGND VPWR VPWR RF.registers\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_4684_ RF.registers\[12\]\[22\] RF.registers\[13\]\[22\] RF.registers\[14\]\[22\]
+ RF.registers\[15\]\[22\] _1192_ _1195_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6423_ RF.registers\[17\]\[5\] _3103_ _3093_ VGND VGND VPWR VPWR _3104_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9142_ clknet_leaf_33_CLK _0302_ VGND VGND VPWR VPWR RF.registers\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_6354_ net21 VGND VGND VPWR VPWR _3056_ sky130_fd_sc_hd__buf_2
XFILLER_0_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6285_ _3008_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__clkbuf_1
X_9073_ clknet_leaf_7_CLK _0233_ VGND VGND VPWR VPWR RF.registers\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5305_ _1699_ _2060_ _1670_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__o21ai_1
X_8024_ _3980_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__clkbuf_1
X_5236_ _1889_ _1991_ VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5167_ _1777_ _1912_ _1916_ _1922_ VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__o2bb2a_2
X_5098_ RF.registers\[4\]\[17\] RF.registers\[5\]\[17\] RF.registers\[6\]\[17\] RF.registers\[7\]\[17\]
+ _1822_ _1823_ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_3_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8926_ clknet_leaf_67_CLK _0086_ VGND VGND VPWR VPWR RF.registers\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8857_ clknet_leaf_50_CLK _0017_ VGND VGND VPWR VPWR RF.registers\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8788_ clknet_leaf_53_CLK _0972_ VGND VGND VPWR VPWR RF.registers\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7808_ _3843_ VGND VGND VPWR VPWR _3866_ sky130_fd_sc_hd__buf_4
X_7739_ _3829_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9409_ clknet_leaf_79_CLK _0569_ VGND VGND VPWR VPWR RF.registers\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_49_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6070_ _1798_ _2805_ VGND VGND VPWR VPWR _2806_ sky130_fd_sc_hd__nor2_1
X_5021_ _1729_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6972_ _3406_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
X_8711_ clknet_leaf_59_CLK _0895_ VGND VGND VPWR VPWR RF.registers\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5923_ _2645_ _2642_ _2664_ _2635_ _2666_ VGND VGND VPWR VPWR _2667_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_48_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5854_ _2600_ _2601_ VGND VGND VPWR VPWR _2602_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8642_ clknet_leaf_76_CLK _0826_ VGND VGND VPWR VPWR RF.registers\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8573_ clknet_leaf_15_CLK _0757_ VGND VGND VPWR VPWR RF.registers\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4805_ RF.registers\[16\]\[11\] RF.registers\[17\]\[11\] RF.registers\[18\]\[11\]
+ RF.registers\[19\]\[11\] _1072_ _1073_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__mux4_1
X_5785_ _1059_ _1083_ VGND VGND VPWR VPWR _2535_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7524_ _3052_ RF.registers\[27\]\[14\] _3711_ VGND VGND VPWR VPWR _3716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4736_ _1490_ _1491_ _1287_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4667_ RF.registers\[12\]\[23\] RF.registers\[13\]\[23\] RF.registers\[14\]\[23\]
+ RF.registers\[15\]\[23\] _1267_ _1268_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7455_ _3679_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6406_ _3090_ _3091_ VGND VGND VPWR VPWR _3092_ sky130_fd_sc_hd__nor2_2
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7386_ _3050_ RF.registers\[26\]\[13\] _3639_ VGND VGND VPWR VPWR _3643_ sky130_fd_sc_hd__mux2_1
X_4598_ RF.registers\[16\]\[25\] RF.registers\[17\]\[25\] RF.registers\[18\]\[25\]
+ RF.registers\[19\]\[25\] _1351_ _1352_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__mux4_1
X_6337_ _3043_ RF.registers\[22\]\[10\] _3044_ VGND VGND VPWR VPWR _3045_ sky130_fd_sc_hd__mux2_1
X_9125_ clknet_leaf_64_CLK _0285_ VGND VGND VPWR VPWR RF.registers\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6268_ _1334_ _1904_ VGND VGND VPWR VPWR _2993_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_73_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9056_ clknet_leaf_74_CLK _0216_ VGND VGND VPWR VPWR RF.registers\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_5219_ RF.registers\[0\]\[27\] RF.registers\[1\]\[27\] RF.registers\[2\]\[27\] RF.registers\[3\]\[27\]
+ _1895_ _1897_ VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__mux4_1
X_6199_ _2475_ _2591_ _2652_ _2737_ _2927_ VGND VGND VPWR VPWR _2928_ sky130_fd_sc_hd__a221o_1
X_8007_ _3971_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8909_ clknet_leaf_4_CLK _0069_ VGND VGND VPWR VPWR RF.registers\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5570_ _2307_ _2325_ VGND VGND VPWR VPWR _2326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4521_ _1239_ _1266_ _1272_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_81_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4452_ _1174_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__clkbuf_4
X_7240_ _3041_ RF.registers\[29\]\[9\] _3555_ VGND VGND VPWR VPWR _3565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_84_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7171_ _3527_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4383_ _1038_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__nand2_1
X_6122_ _2840_ _2844_ _2838_ VGND VGND VPWR VPWR _2855_ sky130_fd_sc_hd__o21ai_1
X_6053_ _1800_ _1821_ _2399_ VGND VGND VPWR VPWR _2790_ sky130_fd_sc_hd__o21a_1
X_5004_ RF.registers\[16\]\[21\] RF.registers\[17\]\[21\] RF.registers\[18\]\[21\]
+ RF.registers\[19\]\[21\] _1676_ _1681_ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6955_ _3397_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_37_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5906_ _2648_ _2650_ _2501_ VGND VGND VPWR VPWR _2651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8625_ clknet_leaf_18_CLK _0809_ VGND VGND VPWR VPWR RF.registers\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6886_ RF.registers\[5\]\[19\] _3132_ _3351_ VGND VGND VPWR VPWR _3361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5837_ _1758_ _2331_ _1148_ VGND VGND VPWR VPWR _2585_ sky130_fd_sc_hd__or3b_1
XFILLER_0_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8556_ RF.registers\[10\]\[20\] net26 _4255_ VGND VGND VPWR VPWR _4262_ sky130_fd_sc_hd__mux2_1
X_5768_ _2511_ _2512_ _2509_ VGND VGND VPWR VPWR _2519_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8487_ RF.registers\[11\]\[19\] net24 _4216_ VGND VGND VPWR VPWR _4226_ sky130_fd_sc_hd__mux2_1
X_4719_ _1213_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7507_ _3035_ RF.registers\[27\]\[6\] _3700_ VGND VGND VPWR VPWR _3707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5699_ _2449_ _2451_ VGND VGND VPWR VPWR _2453_ sky130_fd_sc_hd__or2_1
X_7438_ _3670_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7369_ _3033_ RF.registers\[26\]\[5\] _3628_ VGND VGND VPWR VPWR _3634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9108_ clknet_leaf_23_CLK _0268_ VGND VGND VPWR VPWR RF.registers\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_9039_ clknet_leaf_5_CLK _0199_ VGND VGND VPWR VPWR RF.registers\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6740_ _3283_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6671_ RF.registers\[8\]\[14\] _3122_ _3242_ VGND VGND VPWR VPWR _3247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5622_ _1168_ _1905_ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__and2_1
X_9390_ clknet_leaf_20_CLK _0550_ VGND VGND VPWR VPWR RF.registers\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8410_ _4185_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5553_ RF.registers\[16\]\[5\] RF.registers\[17\]\[5\] RF.registers\[18\]\[5\] RF.registers\[19\]\[5\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2309_ sky130_fd_sc_hd__mux4_1
X_8341_ RF.registers\[16\]\[14\] _3485_ _4144_ VGND VGND VPWR VPWR _4149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4504_ _1257_ _1258_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_8272_ _4112_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__clkbuf_1
X_5484_ _2238_ _2239_ _1685_ VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7223_ _3556_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4435_ _1072_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4366_ RF.registers\[12\]\[2\] RF.registers\[13\]\[2\] RF.registers\[14\]\[2\] RF.registers\[15\]\[2\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__mux4_1
X_7154_ RF.registers\[7\]\[1\] _3458_ _3517_ VGND VGND VPWR VPWR _3519_ sky130_fd_sc_hd__mux2_1
X_6105_ _1754_ _2837_ VGND VGND VPWR VPWR _2839_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_70_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4297_ _1043_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__buf_4
X_7085_ net45 VGND VGND VPWR VPWR _3474_ sky130_fd_sc_hd__buf_2
X_6036_ _2749_ _2771_ _2773_ VGND VGND VPWR VPWR _2774_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7987_ _3109_ RF.registers\[21\]\[8\] _3952_ VGND VGND VPWR VPWR _3961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6938_ RF.registers\[4\]\[11\] _3116_ _3387_ VGND VGND VPWR VPWR _3389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6869_ _3352_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9588_ clknet_leaf_42_CLK _0748_ VGND VGND VPWR VPWR RF.registers\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8608_ clknet_leaf_70_CLK _0792_ VGND VGND VPWR VPWR RF.registers\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8539_ RF.registers\[10\]\[12\] net17 _4244_ VGND VGND VPWR VPWR _4253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8890_ clknet_leaf_34_CLK _0050_ VGND VGND VPWR VPWR RF.registers\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_7910_ _3920_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__clkbuf_1
X_7841_ _3099_ RF.registers\[23\]\[3\] _3880_ VGND VGND VPWR VPWR _3884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4984_ _1736_ _1737_ _1739_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7772_ _3847_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6723_ _3274_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__clkbuf_1
X_9511_ clknet_leaf_81_CLK _0671_ VGND VGND VPWR VPWR RF.registers\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9442_ clknet_leaf_91_CLK _0602_ VGND VGND VPWR VPWR RF.registers\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6654_ RF.registers\[8\]\[6\] _3105_ _3231_ VGND VGND VPWR VPWR _3238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5605_ _1668_ _2324_ VGND VGND VPWR VPWR _2360_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9373_ clknet_leaf_18_CLK _0533_ VGND VGND VPWR VPWR RF.registers\[20\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6585_ _3201_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5536_ _2290_ _2291_ _2044_ VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__mux2_1
X_8324_ RF.registers\[16\]\[6\] _3468_ _4133_ VGND VGND VPWR VPWR _4140_ sky130_fd_sc_hd__mux2_1
X_5467_ _2221_ _2222_ _1712_ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__mux2_1
X_8255_ _4103_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7206_ RF.registers\[7\]\[26\] _3442_ _3539_ VGND VGND VPWR VPWR _3546_ sky130_fd_sc_hd__mux2_1
X_4418_ _1073_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__buf_4
X_8186_ RF.registers\[1\]\[5\] _3466_ _4061_ VGND VGND VPWR VPWR _4067_ sky130_fd_sc_hd__mux2_1
X_5398_ RF.registers\[0\]\[13\] RF.registers\[1\]\[13\] RF.registers\[2\]\[13\] RF.registers\[3\]\[13\]
+ _1702_ _1678_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__mux4_1
X_7137_ _3509_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
X_4349_ _1043_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__clkbuf_4
X_7068_ RF.registers\[19\]\[3\] _3462_ _3456_ VGND VGND VPWR VPWR _3463_ sky130_fd_sc_hd__mux2_1
X_6019_ _1127_ _2524_ _2737_ _2503_ VGND VGND VPWR VPWR _2758_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6370_ net27 VGND VGND VPWR VPWR _3067_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5321_ RF.registers\[0\]\[2\] RF.registers\[1\]\[2\] RF.registers\[2\]\[2\] RF.registers\[3\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8040_ RF.registers\[20\]\[0\] _3454_ _3989_ VGND VGND VPWR VPWR _3990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5252_ RF.registers\[12\]\[25\] RF.registers\[13\]\[25\] RF.registers\[14\]\[25\]
+ RF.registers\[15\]\[25\] _1895_ _1897_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5183_ RF.registers\[12\]\[29\] RF.registers\[13\]\[29\] RF.registers\[14\]\[29\]
+ RF.registers\[15\]\[29\] _1767_ _1768_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8942_ clknet_leaf_13_CLK _0102_ VGND VGND VPWR VPWR RF.registers\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8873_ clknet_leaf_86_CLK _0033_ VGND VGND VPWR VPWR RF.registers\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_7824_ _3874_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7755_ _3079_ RF.registers\[30\]\[27\] _3830_ VGND VGND VPWR VPWR _3838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4967_ _1722_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7686_ _3801_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__clkbuf_1
X_6706_ RF.registers\[8\]\[31\] _3017_ _3230_ VGND VGND VPWR VPWR _3265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4898_ net4 _1653_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6637_ _3228_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__clkbuf_1
X_9425_ clknet_leaf_55_CLK _0585_ VGND VGND VPWR VPWR RF.registers\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6568_ RF.registers\[0\]\[31\] _3017_ _3156_ VGND VGND VPWR VPWR _3191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9356_ clknet_leaf_2_CLK _0516_ VGND VGND VPWR VPWR RF.registers\[20\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8307_ _4130_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5519_ RF.registers\[16\]\[7\] RF.registers\[17\]\[7\] RF.registers\[18\]\[7\] RF.registers\[19\]\[7\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__mux4_1
XFILLER_0_131_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6499_ net13 net12 net11 VGND VGND VPWR VPWR _3153_ sky130_fd_sc_hd__or3_4
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9287_ clknet_leaf_83_CLK _0447_ VGND VGND VPWR VPWR RF.registers\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8238_ RF.registers\[1\]\[30\] _3450_ _4060_ VGND VGND VPWR VPWR _4094_ sky130_fd_sc_hd__mux2_1
X_8169_ _4057_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_93_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5870_ _2246_ _2616_ VGND VGND VPWR VPWR _2617_ sky130_fd_sc_hd__xor2_2
X_4821_ RF.registers\[20\]\[16\] RF.registers\[21\]\[16\] RF.registers\[22\]\[16\]
+ RF.registers\[23\]\[16\] _1291_ _1194_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7540_ _3724_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
X_4752_ RF.registers\[0\]\[15\] RF.registers\[1\]\[15\] RF.registers\[2\]\[15\] RF.registers\[3\]\[15\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7471_ _3067_ RF.registers\[25\]\[21\] _3686_ VGND VGND VPWR VPWR _3688_ sky130_fd_sc_hd__mux2_1
X_4683_ _1189_ _1438_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9210_ clknet_leaf_25_CLK _0370_ VGND VGND VPWR VPWR RF.registers\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6422_ net41 VGND VGND VPWR VPWR _3103_ sky130_fd_sc_hd__buf_2
X_9141_ clknet_leaf_28_CLK _0301_ VGND VGND VPWR VPWR RF.registers\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6353_ _3055_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6284_ RF.registers\[10\]\[26\] _3002_ _3007_ VGND VGND VPWR VPWR _3008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9072_ clknet_leaf_8_CLK _0232_ VGND VGND VPWR VPWR RF.registers\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_5304_ _2058_ _2059_ _1685_ VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__mux2_1
X_8023_ _3145_ RF.registers\[21\]\[25\] _3974_ VGND VGND VPWR VPWR _3980_ sky130_fd_sc_hd__mux2_1
X_5235_ RF.registers\[4\]\[26\] RF.registers\[5\]\[26\] RF.registers\[6\]\[26\] RF.registers\[7\]\[26\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5166_ _1766_ _1921_ _1672_ VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__o21ai_1
X_5097_ _1700_ _1852_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__nand2_1
X_8925_ clknet_leaf_18_CLK _0085_ VGND VGND VPWR VPWR RF.registers\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8856_ clknet_leaf_40_CLK _0016_ VGND VGND VPWR VPWR RF.registers\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_8787_ clknet_leaf_50_CLK _0971_ VGND VGND VPWR VPWR RF.registers\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7807_ _3865_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__clkbuf_1
X_5999_ _2585_ _2738_ _2333_ VGND VGND VPWR VPWR _2739_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7738_ _3062_ RF.registers\[30\]\[19\] _3819_ VGND VGND VPWR VPWR _3829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7669_ _3792_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
X_9408_ clknet_leaf_69_CLK _0568_ VGND VGND VPWR VPWR RF.registers\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9339_ clknet_leaf_45_CLK _0499_ VGND VGND VPWR VPWR RF.registers\[21\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_113_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_122_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5020_ _1774_ _1775_ _1726_ VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_131_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6971_ RF.registers\[4\]\[27\] _3009_ _3398_ VGND VGND VPWR VPWR _3406_ sky130_fd_sc_hd__mux2_1
X_8710_ clknet_leaf_61_CLK _0894_ VGND VGND VPWR VPWR RF.registers\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5922_ _2193_ _2640_ _2641_ VGND VGND VPWR VPWR _2666_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5853_ _2539_ _2559_ _2560_ VGND VGND VPWR VPWR _2601_ sky130_fd_sc_hd__o21ai_2
X_8641_ clknet_leaf_72_CLK _0825_ VGND VGND VPWR VPWR RF.registers\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_8572_ clknet_leaf_16_CLK _0756_ VGND VGND VPWR VPWR RF.registers\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5784_ _2534_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_1
X_4804_ RF.registers\[28\]\[11\] RF.registers\[29\]\[11\] RF.registers\[30\]\[11\]
+ RF.registers\[31\]\[11\] _1042_ _1044_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__mux4_1
X_7523_ _3715_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_32_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4735_ RF.registers\[12\]\[14\] RF.registers\[13\]\[14\] RF.registers\[14\]\[14\]
+ RF.registers\[15\]\[14\] _1172_ _1279_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4666_ RF.registers\[8\]\[23\] RF.registers\[9\]\[23\] RF.registers\[10\]\[23\] RF.registers\[11\]\[23\]
+ _1267_ _1268_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7454_ _3050_ RF.registers\[25\]\[13\] _3675_ VGND VGND VPWR VPWR _3679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4597_ RF.registers\[20\]\[25\] RF.registers\[21\]\[25\] RF.registers\[22\]\[25\]
+ RF.registers\[23\]\[25\] _1351_ _1352_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__mux4_1
X_6405_ net10 net9 net46 VGND VGND VPWR VPWR _3091_ sky130_fd_sc_hd__nand3b_4
X_7385_ _3642_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6336_ _3022_ VGND VGND VPWR VPWR _3044_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9124_ clknet_leaf_94_CLK _0284_ VGND VGND VPWR VPWR RF.registers\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_9055_ clknet_leaf_73_CLK _0215_ VGND VGND VPWR VPWR RF.registers\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6267_ _1348_ _2981_ _2741_ VGND VGND VPWR VPWR _2992_ sky130_fd_sc_hd__a21o_1
X_5218_ RF.registers\[4\]\[27\] RF.registers\[5\]\[27\] RF.registers\[6\]\[27\] RF.registers\[7\]\[27\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__mux4_1
X_6198_ _2530_ _2792_ _2922_ _2926_ VGND VGND VPWR VPWR _2927_ sky130_fd_sc_hd__o211a_1
X_8006_ _3128_ RF.registers\[21\]\[17\] _3963_ VGND VGND VPWR VPWR _3971_ sky130_fd_sc_hd__mux2_1
X_5149_ _1842_ _1904_ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8908_ clknet_leaf_3_CLK _0068_ VGND VGND VPWR VPWR RF.registers\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8839_ clknet_leaf_60_CLK _1023_ VGND VGND VPWR VPWR RF.registers\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4520_ _1254_ _1275_ _1171_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4451_ _1191_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7170_ RF.registers\[7\]\[9\] _3474_ _3517_ VGND VGND VPWR VPWR _3527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6121_ _1731_ _2853_ VGND VGND VPWR VPWR _2854_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_59_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4382_ _1136_ _1137_ _1047_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6052_ _2421_ _2788_ VGND VGND VPWR VPWR _2789_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5003_ RF.registers\[20\]\[21\] RF.registers\[21\]\[21\] RF.registers\[22\]\[21\]
+ RF.registers\[23\]\[21\] _1676_ _1681_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__mux4_1
X_6954_ RF.registers\[4\]\[19\] _3132_ _3387_ VGND VGND VPWR VPWR _3397_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5905_ _2609_ _2649_ _1803_ VGND VGND VPWR VPWR _2650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6885_ _3360_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__clkbuf_1
X_8624_ clknet_leaf_7_CLK _0808_ VGND VGND VPWR VPWR RF.registers\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5836_ _2579_ _2583_ _2252_ VGND VGND VPWR VPWR _2584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8555_ _4261_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5767_ _2516_ _2517_ VGND VGND VPWR VPWR _2518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8486_ _4225_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__clkbuf_1
X_5698_ _2449_ _2451_ VGND VGND VPWR VPWR _2452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7506_ _3706_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4718_ _1472_ _1473_ _1287_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7437_ _3033_ RF.registers\[25\]\[5\] _3664_ VGND VGND VPWR VPWR _3670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4649_ _1403_ _1404_ _1107_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7368_ _3633_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
X_9107_ clknet_leaf_26_CLK _0267_ VGND VGND VPWR VPWR RF.registers\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6319_ _3032_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__clkbuf_1
X_7299_ _3596_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_9038_ clknet_leaf_21_CLK _0198_ VGND VGND VPWR VPWR RF.registers\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6670_ _3246_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5621_ _2335_ _2337_ _2340_ _2375_ _2333_ VGND VGND VPWR VPWR _2376_ sky130_fd_sc_hd__o311a_1
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5552_ RF.registers\[20\]\[5\] RF.registers\[21\]\[5\] RF.registers\[22\]\[5\] RF.registers\[23\]\[5\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2308_ sky130_fd_sc_hd__mux4_1
X_8340_ _4148_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4503_ _1036_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8271_ _3120_ RF.registers\[13\]\[13\] _4108_ VGND VGND VPWR VPWR _4112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5483_ RF.registers\[8\]\[9\] RF.registers\[9\]\[9\] RF.registers\[10\]\[9\] RF.registers\[11\]\[9\]
+ _1782_ _1692_ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4434_ _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_57_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7222_ _3019_ RF.registers\[29\]\[0\] _3555_ VGND VGND VPWR VPWR _3556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7153_ _3518_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_4365_ RF.registers\[8\]\[2\] RF.registers\[9\]\[2\] RF.registers\[10\]\[2\] RF.registers\[11\]\[2\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__mux4_1
X_6104_ _1754_ _2837_ VGND VGND VPWR VPWR _2838_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7084_ _3473_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
X_6035_ _1858_ _2762_ _2772_ VGND VGND VPWR VPWR _2773_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_70_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _1041_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7986_ _3960_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6937_ _3388_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6868_ RF.registers\[5\]\[10\] _3113_ _3351_ VGND VGND VPWR VPWR _3352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9587_ clknet_leaf_29_CLK _0747_ VGND VGND VPWR VPWR RF.registers\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_5819_ _2458_ _2567_ _1126_ VGND VGND VPWR VPWR _2568_ sky130_fd_sc_hd__mux2_1
X_8607_ clknet_leaf_71_CLK _0791_ VGND VGND VPWR VPWR RF.registers\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6799_ _3303_ VGND VGND VPWR VPWR _3315_ sky130_fd_sc_hd__buf_4
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8538_ _4252_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8469_ RF.registers\[11\]\[10\] net15 _4216_ VGND VGND VPWR VPWR _4217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7840_ _3883_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4983_ _1738_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__clkbuf_8
X_7771_ RF.registers\[9\]\[2\] _3460_ _3844_ VGND VGND VPWR VPWR _3847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6722_ _3035_ RF.registers\[14\]\[6\] _3267_ VGND VGND VPWR VPWR _3274_ sky130_fd_sc_hd__mux2_1
X_9510_ clknet_leaf_63_CLK _0670_ VGND VGND VPWR VPWR RF.registers\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9441_ clknet_leaf_93_CLK _0601_ VGND VGND VPWR VPWR RF.registers\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6653_ _3237_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5604_ _2357_ _2358_ VGND VGND VPWR VPWR _2359_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9372_ clknet_leaf_16_CLK _0532_ VGND VGND VPWR VPWR RF.registers\[20\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6584_ _3033_ RF.registers\[15\]\[5\] _3195_ VGND VGND VPWR VPWR _3201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5535_ RF.registers\[16\]\[4\] RF.registers\[17\]\[4\] RF.registers\[18\]\[4\] RF.registers\[19\]\[4\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__mux4_1
X_8323_ _4139_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8254_ _3103_ RF.registers\[13\]\[5\] _4097_ VGND VGND VPWR VPWR _4103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5466_ RF.registers\[12\]\[8\] RF.registers\[13\]\[8\] RF.registers\[14\]\[8\] RF.registers\[15\]\[8\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__mux4_1
X_7205_ _3545_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4417_ _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8185_ _4066_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5397_ _1684_ _2152_ VGND VGND VPWR VPWR _2153_ sky130_fd_sc_hd__or2_1
X_7136_ RF.registers\[19\]\[25\] _3508_ _3498_ VGND VGND VPWR VPWR _3509_ sky130_fd_sc_hd__mux2_1
X_4348_ _1041_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__buf_4
X_7067_ net39 VGND VGND VPWR VPWR _3462_ sky130_fd_sc_hd__clkbuf_4
X_4279_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_87_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6018_ _2527_ _2756_ _2426_ VGND VGND VPWR VPWR _2757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7969_ _3021_ _3552_ VGND VGND VPWR VPWR _3951_ sky130_fd_sc_hd__nand2_4
XFILLER_0_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5320_ RF.registers\[4\]\[2\] RF.registers\[5\]\[2\] RF.registers\[6\]\[2\] RF.registers\[7\]\[2\]
+ _1701_ _1677_ VGND VGND VPWR VPWR _2076_ sky130_fd_sc_hd__mux4_1
X_5251_ RF.registers\[8\]\[25\] RF.registers\[9\]\[25\] RF.registers\[10\]\[25\] RF.registers\[11\]\[25\]
+ _1895_ _1897_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_54_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5182_ RF.registers\[8\]\[29\] RF.registers\[9\]\[29\] RF.registers\[10\]\[29\] RF.registers\[11\]\[29\]
+ _1767_ _1768_ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8941_ clknet_leaf_83_CLK _0101_ VGND VGND VPWR VPWR RF.registers\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8872_ clknet_leaf_78_CLK _0032_ VGND VGND VPWR VPWR RF.registers\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_7823_ RF.registers\[9\]\[27\] _3444_ _3866_ VGND VGND VPWR VPWR _3874_ sky130_fd_sc_hd__mux2_1
X_7754_ _3837_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_96_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_96_CLK sky130_fd_sc_hd__clkbuf_8
X_6705_ _3264_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4966_ _1721_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__buf_4
X_7685_ RF.registers\[2\]\[26\] _3442_ _3794_ VGND VGND VPWR VPWR _3801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4897_ _1651_ _1652_ net3 VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6636_ _3085_ RF.registers\[15\]\[30\] _3194_ VGND VGND VPWR VPWR _3228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9424_ clknet_leaf_57_CLK _0584_ VGND VGND VPWR VPWR RF.registers\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6567_ _3190_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9355_ clknet_leaf_1_CLK _0515_ VGND VGND VPWR VPWR RF.registers\[20\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8306_ _3015_ RF.registers\[13\]\[30\] _4096_ VGND VGND VPWR VPWR _4130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5518_ RF.registers\[28\]\[7\] RF.registers\[29\]\[7\] RF.registers\[30\]\[7\] RF.registers\[31\]\[7\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2274_ sky130_fd_sc_hd__mux4_1
X_6498_ _3152_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__clkbuf_1
X_9286_ clknet_leaf_62_CLK _0446_ VGND VGND VPWR VPWR RF.registers\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8237_ _4093_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__clkbuf_1
X_5449_ _1699_ _2204_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__nand2_1
X_8168_ RF.registers\[24\]\[29\] _3448_ _4047_ VGND VGND VPWR VPWR _4057_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_20_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7119_ net26 VGND VGND VPWR VPWR _3497_ sky130_fd_sc_hd__buf_2
X_8099_ _4020_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_87_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_87_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_11_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_127_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4820_ RF.registers\[16\]\[16\] RF.registers\[17\]\[16\] RF.registers\[18\]\[16\]
+ RF.registers\[19\]\[16\] _1291_ _1194_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_78_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_78_CLK sky130_fd_sc_hd__clkbuf_8
X_4751_ RF.registers\[4\]\[15\] RF.registers\[5\]\[15\] RF.registers\[6\]\[15\] RF.registers\[7\]\[15\]
+ _1192_ _1195_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4682_ RF.registers\[8\]\[22\] RF.registers\[9\]\[22\] RF.registers\[10\]\[22\] RF.registers\[11\]\[22\]
+ _1207_ _1208_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__mux4_1
X_7470_ _3687_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6421_ _3102_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9140_ clknet_leaf_24_CLK _0300_ VGND VGND VPWR VPWR RF.registers\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6352_ _3054_ RF.registers\[22\]\[15\] _3044_ VGND VGND VPWR VPWR _3055_ sky130_fd_sc_hd__mux2_1
X_6283_ _3006_ VGND VGND VPWR VPWR _3007_ sky130_fd_sc_hd__buf_6
X_9071_ clknet_leaf_4_CLK _0231_ VGND VGND VPWR VPWR RF.registers\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_5303_ RF.registers\[0\]\[3\] RF.registers\[1\]\[3\] RF.registers\[2\]\[3\] RF.registers\[3\]\[3\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__mux4_1
X_8022_ _3979_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__clkbuf_1
X_5234_ _1988_ _1989_ _1901_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__mux2_1
X_5165_ _1917_ _1920_ _1901_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5096_ _1850_ _1851_ _1713_ VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__mux2_1
X_8924_ clknet_leaf_18_CLK _0084_ VGND VGND VPWR VPWR RF.registers\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8855_ clknet_leaf_49_CLK _0015_ VGND VGND VPWR VPWR RF.registers\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7806_ RF.registers\[9\]\[19\] _3495_ _3855_ VGND VGND VPWR VPWR _3865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8786_ clknet_leaf_43_CLK _0970_ VGND VGND VPWR VPWR RF.registers\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5998_ _1127_ _2737_ VGND VGND VPWR VPWR _2738_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_69_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_69_CLK sky130_fd_sc_hd__clkbuf_8
X_4949_ _1704_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__buf_6
X_7737_ _3828_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7668_ RF.registers\[2\]\[18\] _3493_ _3783_ VGND VGND VPWR VPWR _3792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6619_ _3219_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9407_ clknet_leaf_66_CLK _0567_ VGND VGND VPWR VPWR RF.registers\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_95_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7599_ _3755_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9338_ clknet_leaf_37_CLK _0498_ VGND VGND VPWR VPWR RF.registers\[21\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9269_ clknet_leaf_28_CLK _0429_ VGND VGND VPWR VPWR RF.registers\[23\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_CLK clknet_3_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6970_ _3405_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
X_5921_ _2598_ _2617_ _2664_ VGND VGND VPWR VPWR _2665_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_49_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5852_ _2511_ _2512_ _2518_ _2542_ _2599_ VGND VGND VPWR VPWR _2600_ sky130_fd_sc_hd__a311o_1
X_8640_ clknet_leaf_69_CLK _0824_ VGND VGND VPWR VPWR RF.registers\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8571_ clknet_leaf_45_CLK _0755_ VGND VGND VPWR VPWR RF.registers\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5783_ _2521_ _2529_ _2533_ VGND VGND VPWR VPWR _2534_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_62_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ RF.registers\[24\]\[11\] RF.registers\[25\]\[11\] RF.registers\[26\]\[11\]
+ RF.registers\[27\]\[11\] _1072_ _1073_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__mux4_1
X_4734_ RF.registers\[8\]\[14\] RF.registers\[9\]\[14\] RF.registers\[10\]\[14\] RF.registers\[11\]\[14\]
+ _1172_ _1279_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__mux4_1
X_7522_ _3050_ RF.registers\[27\]\[13\] _3711_ VGND VGND VPWR VPWR _3715_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4665_ _1417_ _1418_ _1419_ _1420_ _1190_ _1205_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__mux4_2
XFILLER_0_71_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7453_ _3678_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4596_ _1325_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6404_ net12 net11 net13 VGND VGND VPWR VPWR _3090_ sky130_fd_sc_hd__or3b_2
X_7384_ _3048_ RF.registers\[26\]\[12\] _3639_ VGND VGND VPWR VPWR _3642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9123_ clknet_leaf_74_CLK _0283_ VGND VGND VPWR VPWR RF.registers\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_6335_ net15 VGND VGND VPWR VPWR _3043_ sky130_fd_sc_hd__clkbuf_2
X_9054_ clknet_leaf_69_CLK _0214_ VGND VGND VPWR VPWR RF.registers\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6266_ _2952_ _2986_ _2987_ _2984_ VGND VGND VPWR VPWR _2991_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_90_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8005_ _3970_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__clkbuf_1
X_5217_ _1773_ _1972_ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__nor2_1
X_6197_ _2337_ _2925_ _1086_ VGND VGND VPWR VPWR _2926_ sky130_fd_sc_hd__o21a_1
X_5148_ _1777_ _1890_ _1894_ _1903_ VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__o2bb2a_2
X_5079_ RF.registers\[0\]\[19\] RF.registers\[1\]\[19\] RF.registers\[2\]\[19\] RF.registers\[3\]\[19\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__mux4_1
X_8907_ clknet_leaf_98_CLK _0067_ VGND VGND VPWR VPWR RF.registers\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8838_ clknet_leaf_61_CLK _1022_ VGND VGND VPWR VPWR RF.registers\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8769_ clknet_leaf_79_CLK _0953_ VGND VGND VPWR VPWR RF.registers\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4450_ _1199_ _1204_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4381_ RF.registers\[12\]\[1\] RF.registers\[13\]\[1\] RF.registers\[14\]\[1\] RF.registers\[15\]\[1\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6120_ _1430_ _2852_ VGND VGND VPWR VPWR _2853_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_59_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6051_ _2784_ _2787_ VGND VGND VPWR VPWR _2788_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_72_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _1639_ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__buf_2
XFILLER_0_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6953_ _3396_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_37_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6884_ RF.registers\[5\]\[18\] _3130_ _3351_ VGND VGND VPWR VPWR _3360_ sky130_fd_sc_hd__mux2_1
X_5904_ _2352_ _2350_ VGND VGND VPWR VPWR _2649_ sky130_fd_sc_hd__and2_1
X_5835_ _2547_ _2582_ _2363_ VGND VGND VPWR VPWR _2583_ sky130_fd_sc_hd__mux2_1
X_8623_ clknet_leaf_4_CLK _0807_ VGND VGND VPWR VPWR RF.registers\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8554_ RF.registers\[10\]\[19\] net24 _4255_ VGND VGND VPWR VPWR _4261_ sky130_fd_sc_hd__mux2_1
X_5766_ _2323_ _2515_ VGND VGND VPWR VPWR _2517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8485_ RF.registers\[11\]\[18\] net23 _4216_ VGND VGND VPWR VPWR _4225_ sky130_fd_sc_hd__mux2_1
X_5697_ _2450_ _2414_ _2413_ VGND VGND VPWR VPWR _2451_ sky130_fd_sc_hd__o21bai_1
X_7505_ _3033_ RF.registers\[27\]\[5\] _3700_ VGND VGND VPWR VPWR _3706_ sky130_fd_sc_hd__mux2_1
X_4717_ RF.registers\[12\]\[13\] RF.registers\[13\]\[13\] RF.registers\[14\]\[13\]
+ RF.registers\[15\]\[13\] _1291_ _1194_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__mux4_1
X_7436_ _3669_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4648_ RF.registers\[24\]\[7\] RF.registers\[25\]\[7\] RF.registers\[26\]\[7\] RF.registers\[27\]\[7\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__mux4_1
X_9106_ clknet_leaf_41_CLK _0266_ VGND VGND VPWR VPWR RF.registers\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_4579_ RF.registers\[24\]\[30\] RF.registers\[25\]\[30\] RF.registers\[26\]\[30\]
+ RF.registers\[27\]\[30\] _1267_ _1268_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__mux4_1
X_7367_ _3031_ RF.registers\[26\]\[4\] _3628_ VGND VGND VPWR VPWR _3633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6318_ _3031_ RF.registers\[22\]\[4\] _3023_ VGND VGND VPWR VPWR _3032_ sky130_fd_sc_hd__mux2_1
X_7298_ _3031_ RF.registers\[31\]\[4\] _3591_ VGND VGND VPWR VPWR _3596_ sky130_fd_sc_hd__mux2_1
X_6249_ _1148_ _1925_ VGND VGND VPWR VPWR _2975_ sky130_fd_sc_hd__nand2_1
X_9037_ clknet_leaf_4_CLK _0197_ VGND VGND VPWR VPWR RF.registers\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5620_ _2105_ _2356_ _2374_ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5551_ _1799_ _2306_ VGND VGND VPWR VPWR _2307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4502_ RF.registers\[16\]\[21\] RF.registers\[17\]\[21\] RF.registers\[18\]\[21\]
+ RF.registers\[19\]\[21\] _1220_ _1222_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8270_ _4111_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7221_ _3554_ VGND VGND VPWR VPWR _3555_ sky130_fd_sc_hd__buf_6
XFILLER_0_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5482_ RF.registers\[12\]\[9\] RF.registers\[13\]\[9\] RF.registers\[14\]\[9\] RF.registers\[15\]\[9\]
+ _1782_ _1680_ VGND VGND VPWR VPWR _2238_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4433_ _1048_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__clkbuf_8
X_4364_ _1047_ _1119_ _1050_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__o21a_1
X_7152_ RF.registers\[7\]\[0\] _3454_ _3517_ VGND VGND VPWR VPWR _3518_ sky130_fd_sc_hd__mux2_1
X_6103_ _1446_ _2836_ VGND VGND VPWR VPWR _2837_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4295_ _1048_ _1049_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__o21a_1
X_7083_ RF.registers\[19\]\[8\] _3472_ _3456_ VGND VGND VPWR VPWR _3473_ sky130_fd_sc_hd__mux2_1
X_6034_ _1874_ _2743_ _2762_ _1858_ VGND VGND VPWR VPWR _2772_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7985_ _3107_ RF.registers\[21\]\[7\] _3952_ VGND VGND VPWR VPWR _3960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6936_ RF.registers\[4\]\[10\] _3113_ _3387_ VGND VGND VPWR VPWR _3388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6867_ _3339_ VGND VGND VPWR VPWR _3351_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9586_ clknet_leaf_56_CLK _0746_ VGND VGND VPWR VPWR RF.registers\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_5818_ _2525_ _2566_ _1146_ VGND VGND VPWR VPWR _2567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8606_ clknet_leaf_68_CLK _0790_ VGND VGND VPWR VPWR RF.registers\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_6798_ _3314_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5749_ _1126_ VGND VGND VPWR VPWR _2501_ sky130_fd_sc_hd__clkbuf_4
X_8537_ RF.registers\[10\]\[11\] net16 _4244_ VGND VGND VPWR VPWR _4252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8468_ _4204_ VGND VGND VPWR VPWR _4216_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_20_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7419_ _3083_ RF.registers\[26\]\[29\] _3650_ VGND VGND VPWR VPWR _3660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8399_ _4179_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput80 net80 VGND VGND VPWR VPWR ALU_result[9] sky130_fd_sc_hd__buf_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4982_ _1684_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__buf_4
X_7770_ _3846_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6721_ _3273_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__clkbuf_1
X_9440_ clknet_leaf_73_CLK _0600_ VGND VGND VPWR VPWR RF.registers\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_6652_ RF.registers\[8\]\[5\] _3103_ _3231_ VGND VGND VPWR VPWR _3237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9371_ clknet_leaf_42_CLK _0531_ VGND VGND VPWR VPWR RF.registers\[20\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_5603_ _1839_ _2230_ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8322_ RF.registers\[16\]\[5\] _3466_ _4133_ VGND VGND VPWR VPWR _4139_ sky130_fd_sc_hd__mux2_1
X_6583_ _3200_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5534_ RF.registers\[20\]\[4\] RF.registers\[21\]\[4\] RF.registers\[22\]\[4\] RF.registers\[23\]\[4\]
+ _2050_ _2052_ VGND VGND VPWR VPWR _2290_ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5465_ RF.registers\[8\]\[8\] RF.registers\[9\]\[8\] RF.registers\[10\]\[8\] RF.registers\[11\]\[8\]
+ _1719_ _1722_ VGND VGND VPWR VPWR _2221_ sky130_fd_sc_hd__mux4_1
X_8253_ _4102_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__clkbuf_1
X_7204_ RF.registers\[7\]\[25\] _3508_ _3539_ VGND VGND VPWR VPWR _3545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8184_ RF.registers\[1\]\[4\] _3464_ _4061_ VGND VGND VPWR VPWR _4066_ sky130_fd_sc_hd__mux2_1
X_4416_ _1072_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__buf_4
X_7135_ net31 VGND VGND VPWR VPWR _3508_ sky130_fd_sc_hd__buf_2
XFILLER_0_100_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5396_ RF.registers\[4\]\[13\] RF.registers\[5\]\[13\] RF.registers\[6\]\[13\] RF.registers\[7\]\[13\]
+ _1702_ _1678_ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__mux4_1
X_4347_ RF.registers\[4\]\[3\] RF.registers\[5\]\[3\] RF.registers\[6\]\[3\] RF.registers\[7\]\[3\]
+ _1089_ _1090_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__mux4_1
X_7066_ _3461_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
X_4278_ net6 VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6017_ _2565_ _2609_ _1148_ VGND VGND VPWR VPWR _2756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7968_ _3950_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__clkbuf_1
X_7899_ _3017_ RF.registers\[23\]\[31\] _3879_ VGND VGND VPWR VPWR _3914_ sky130_fd_sc_hd__mux2_1
X_6919_ RF.registers\[4\]\[2\] _3097_ _3376_ VGND VGND VPWR VPWR _3379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9569_ clknet_leaf_95_CLK _0729_ VGND VGND VPWR VPWR RF.registers\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5250_ _2002_ _2005_ _1700_ VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5181_ _1745_ _1936_ _1697_ VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8940_ clknet_leaf_84_CLK _0100_ VGND VGND VPWR VPWR RF.registers\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8871_ clknet_leaf_59_CLK _0031_ VGND VGND VPWR VPWR RF.registers\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_7822_ _3873_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__clkbuf_1
X_7753_ _3077_ RF.registers\[30\]\[26\] _3830_ VGND VGND VPWR VPWR _3837_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4965_ _1678_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6704_ RF.registers\[8\]\[30\] _3015_ _3230_ VGND VGND VPWR VPWR _3264_ sky130_fd_sc_hd__mux2_1
X_7684_ _3800_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9423_ clknet_leaf_13_CLK _0583_ VGND VGND VPWR VPWR RF.registers\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_4896_ RF.registers\[12\]\[0\] RF.registers\[13\]\[0\] RF.registers\[14\]\[0\] RF.registers\[15\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_22_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6635_ _3227_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6566_ RF.registers\[0\]\[30\] _3015_ _3156_ VGND VGND VPWR VPWR _3190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9354_ clknet_leaf_9_CLK _0514_ VGND VGND VPWR VPWR RF.registers\[20\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8305_ _4129_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__clkbuf_1
X_9285_ clknet_leaf_63_CLK _0445_ VGND VGND VPWR VPWR RF.registers\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_5517_ RF.registers\[24\]\[7\] RF.registers\[25\]\[7\] RF.registers\[26\]\[7\] RF.registers\[27\]\[7\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2273_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8236_ RF.registers\[1\]\[29\] _3448_ _4083_ VGND VGND VPWR VPWR _4093_ sky130_fd_sc_hd__mux2_1
X_6497_ RF.registers\[17\]\[31\] _3017_ _3092_ VGND VGND VPWR VPWR _3152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5448_ _2202_ _2203_ _1711_ VGND VGND VPWR VPWR _2204_ sky130_fd_sc_hd__mux2_1
X_8167_ _4056_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5379_ _1699_ _2134_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__nand2_1
X_8098_ RF.registers\[20\]\[28\] _3446_ _4011_ VGND VGND VPWR VPWR _4020_ sky130_fd_sc_hd__mux2_1
X_7118_ _3496_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_7049_ _3449_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4750_ _1214_ _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4681_ _1433_ _1436_ _1187_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6420_ RF.registers\[17\]\[4\] _3101_ _3093_ VGND VGND VPWR VPWR _3102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6351_ net20 VGND VGND VPWR VPWR _3054_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5302_ RF.registers\[4\]\[3\] RF.registers\[5\]\[3\] RF.registers\[6\]\[3\] RF.registers\[7\]\[3\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__mux4_1
XFILLER_0_122_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6282_ _3003_ _3005_ VGND VGND VPWR VPWR _3006_ sky130_fd_sc_hd__nor2_4
X_9070_ clknet_leaf_5_CLK _0230_ VGND VGND VPWR VPWR RF.registers\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8021_ _3143_ RF.registers\[21\]\[24\] _3974_ VGND VGND VPWR VPWR _3979_ sky130_fd_sc_hd__mux2_1
X_5233_ RF.registers\[8\]\[26\] RF.registers\[9\]\[26\] RF.registers\[10\]\[26\] RF.registers\[11\]\[26\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5164_ RF.registers\[0\]\[30\] RF.registers\[1\]\[30\] RF.registers\[2\]\[30\] RF.registers\[3\]\[30\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__mux4_1
XFILLER_0_79_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5095_ RF.registers\[12\]\[17\] RF.registers\[13\]\[17\] RF.registers\[14\]\[17\]
+ RF.registers\[15\]\[17\] _1720_ _1723_ VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__mux4_1
X_8923_ clknet_leaf_46_CLK _0083_ VGND VGND VPWR VPWR RF.registers\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8854_ clknet_leaf_49_CLK _0014_ VGND VGND VPWR VPWR RF.registers\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7805_ _3864_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5997_ _1060_ _1085_ VGND VGND VPWR VPWR _2737_ sky130_fd_sc_hd__nor2b_2
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8785_ clknet_leaf_56_CLK _0969_ VGND VGND VPWR VPWR RF.registers\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7736_ _3060_ RF.registers\[30\]\[18\] _3819_ VGND VGND VPWR VPWR _3828_ sky130_fd_sc_hd__mux2_1
X_4948_ _1703_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__clkbuf_8
X_4879_ _1602_ _1618_ _1634_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7667_ _3791_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
X_6618_ _3067_ RF.registers\[15\]\[21\] _3217_ VGND VGND VPWR VPWR _3219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9406_ clknet_leaf_67_CLK _0566_ VGND VGND VPWR VPWR RF.registers\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_95_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7598_ _3058_ RF.registers\[28\]\[17\] _3747_ VGND VGND VPWR VPWR _3755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9337_ clknet_leaf_31_CLK _0497_ VGND VGND VPWR VPWR RF.registers\[21\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6549_ _3181_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_95_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9268_ clknet_leaf_37_CLK _0428_ VGND VGND VPWR VPWR RF.registers\[23\]\[22\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8219_ _4084_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__clkbuf_1
X_9199_ clknet_leaf_5_CLK _0359_ VGND VGND VPWR VPWR RF.registers\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_27_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5920_ _2633_ _2642_ _2643_ VGND VGND VPWR VPWR _2664_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_45_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5851_ _2562_ _2560_ _2559_ VGND VGND VPWR VPWR _2599_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8570_ clknet_leaf_36_CLK _0754_ VGND VGND VPWR VPWR RF.registers\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5782_ _2530_ _2531_ _2532_ _2373_ VGND VGND VPWR VPWR _2533_ sky130_fd_sc_hd__o211a_1
X_4802_ _1024_ _1549_ _1553_ _1557_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_90_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4733_ _1287_ _1488_ _1078_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7521_ _3714_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7452_ _3048_ RF.registers\[25\]\[12\] _3675_ VGND VGND VPWR VPWR _3678_ sky130_fd_sc_hd__mux2_1
X_4664_ RF.registers\[20\]\[23\] RF.registers\[21\]\[23\] RF.registers\[22\]\[23\]
+ RF.registers\[23\]\[23\] _1351_ _1352_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_54_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6403_ net14 VGND VGND VPWR VPWR _3089_ sky130_fd_sc_hd__buf_2
X_4595_ _1324_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7383_ _3641_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6334_ _3042_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9122_ clknet_leaf_92_CLK _0282_ VGND VGND VPWR VPWR RF.registers\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6265_ _2966_ _2980_ _2408_ _2990_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__o2bb2a_1
X_9053_ clknet_leaf_22_CLK _0213_ VGND VGND VPWR VPWR RF.registers\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5216_ _1970_ _1971_ _1889_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8004_ _3126_ RF.registers\[21\]\[16\] _3963_ VGND VGND VPWR VPWR _3970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6196_ _2895_ _2924_ _2363_ VGND VGND VPWR VPWR _2925_ sky130_fd_sc_hd__mux2_1
X_5147_ _1766_ _1902_ _1672_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__o21ai_1
X_5078_ RF.registers\[4\]\[19\] RF.registers\[5\]\[19\] RF.registers\[6\]\[19\] RF.registers\[7\]\[19\]
+ _1704_ _1707_ VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__mux4_1
X_8906_ clknet_leaf_7_CLK _0066_ VGND VGND VPWR VPWR RF.registers\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8837_ clknet_leaf_81_CLK _1021_ VGND VGND VPWR VPWR RF.registers\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8768_ clknet_leaf_73_CLK _0952_ VGND VGND VPWR VPWR RF.registers\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7719_ _3807_ VGND VGND VPWR VPWR _3819_ sky130_fd_sc_hd__buf_4
X_8699_ clknet_leaf_45_CLK _0883_ VGND VGND VPWR VPWR RF.registers\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4380_ RF.registers\[8\]\[1\] RF.registers\[9\]\[1\] RF.registers\[10\]\[1\] RF.registers\[11\]\[1\]
+ _1052_ _1053_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_59_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _2785_ _2774_ _2786_ VGND VGND VPWR VPWR _2787_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5001_ _1669_ _1732_ _1756_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_72_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6952_ RF.registers\[4\]\[18\] _3130_ _3387_ VGND VGND VPWR VPWR _3396_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5903_ _2567_ VGND VGND VPWR VPWR _2648_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6883_ _3359_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8622_ clknet_leaf_21_CLK _0806_ VGND VGND VPWR VPWR RF.registers\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_5834_ _2581_ VGND VGND VPWR VPWR _2582_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_62_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8553_ _4260_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__clkbuf_1
X_5765_ _2323_ _2515_ VGND VGND VPWR VPWR _2516_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8484_ _4224_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__clkbuf_1
X_5696_ _1667_ _1660_ VGND VGND VPWR VPWR _2450_ sky130_fd_sc_hd__and2_1
X_7504_ _3705_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
X_4716_ RF.registers\[8\]\[13\] RF.registers\[9\]\[13\] RF.registers\[10\]\[13\] RF.registers\[11\]\[13\]
+ _1291_ _1194_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7435_ _3031_ RF.registers\[25\]\[4\] _3664_ VGND VGND VPWR VPWR _3669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4647_ RF.registers\[28\]\[7\] RF.registers\[29\]\[7\] RF.registers\[30\]\[7\] RF.registers\[31\]\[7\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7366_ _3632_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4578_ _1171_ _1323_ _1333_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__a21o_1
X_9105_ clknet_leaf_7_CLK _0265_ VGND VGND VPWR VPWR RF.registers\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_6317_ net40 VGND VGND VPWR VPWR _3031_ sky130_fd_sc_hd__clkbuf_2
X_7297_ _3595_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_71_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6248_ _2969_ _2973_ _2530_ VGND VGND VPWR VPWR _2974_ sky130_fd_sc_hd__mux2_1
X_9036_ clknet_leaf_3_CLK _0196_ VGND VGND VPWR VPWR RF.registers\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_6179_ _2017_ _1998_ VGND VGND VPWR VPWR _2909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5550_ _1842_ _2305_ VGND VGND VPWR VPWR _2306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4501_ RF.registers\[20\]\[21\] RF.registers\[21\]\[21\] RF.registers\[22\]\[21\]
+ RF.registers\[23\]\[21\] _1220_ _1222_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__mux4_1
X_5481_ _2233_ _2236_ _1828_ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4432_ _1179_ _1186_ _1187_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__mux2_1
X_7220_ _3552_ _3553_ VGND VGND VPWR VPWR _3554_ sky130_fd_sc_hd__nand2_4
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7151_ _3516_ VGND VGND VPWR VPWR _3517_ sky130_fd_sc_hd__clkbuf_8
X_4363_ RF.registers\[0\]\[2\] RF.registers\[1\]\[2\] RF.registers\[2\]\[2\] RF.registers\[3\]\[2\]
+ _1026_ _1061_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6102_ _1512_ _2835_ _1635_ _2658_ _2536_ VGND VGND VPWR VPWR _2836_ sky130_fd_sc_hd__a41o_1
X_4294_ net7 VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_1_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7082_ net44 VGND VGND VPWR VPWR _3472_ sky130_fd_sc_hd__buf_2
X_6033_ _2770_ VGND VGND VPWR VPWR _2771_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7984_ _3959_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6935_ _3375_ VGND VGND VPWR VPWR _3387_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6866_ _3350_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__clkbuf_1
X_8605_ clknet_leaf_18_CLK _0789_ VGND VGND VPWR VPWR RF.registers\[22\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_9585_ clknet_leaf_13_CLK _0745_ VGND VGND VPWR VPWR RF.registers\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_5817_ _2565_ VGND VGND VPWR VPWR _2566_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6797_ RF.registers\[6\]\[9\] _3111_ _3304_ VGND VGND VPWR VPWR _3314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5748_ _2418_ _2499_ _1147_ VGND VGND VPWR VPWR _2500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8536_ _4251_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5679_ _2307_ _2325_ _1148_ VGND VGND VPWR VPWR _2433_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_20_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8467_ _4215_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7418_ _3659_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__clkbuf_1
X_8398_ RF.registers\[12\]\[9\] _3474_ _4169_ VGND VGND VPWR VPWR _4179_ sky130_fd_sc_hd__mux2_1
X_7349_ _3622_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
X_9019_ clknet_leaf_34_CLK _0179_ VGND VGND VPWR VPWR RF.registers\[31\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput70 net70 VGND VGND VPWR VPWR ALU_result[29] sky130_fd_sc_hd__buf_1
XFILLER_0_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4981_ RF.registers\[16\]\[22\] RF.registers\[17\]\[22\] RF.registers\[18\]\[22\]
+ RF.registers\[19\]\[22\] _1734_ _1735_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6720_ _3033_ RF.registers\[14\]\[5\] _3267_ VGND VGND VPWR VPWR _3273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6651_ _3236_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9370_ clknet_leaf_36_CLK _0530_ VGND VGND VPWR VPWR RF.registers\[20\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5602_ _1667_ _2287_ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__or2_1
X_6582_ _3031_ RF.registers\[15\]\[4\] _3195_ VGND VGND VPWR VPWR _3200_ sky130_fd_sc_hd__mux2_1
X_5533_ _1169_ _2272_ _2288_ VGND VGND VPWR VPWR _2289_ sky130_fd_sc_hd__a21oi_1
X_8321_ _4138_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8252_ _3101_ RF.registers\[13\]\[4\] _4097_ VGND VGND VPWR VPWR _4102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5464_ _2216_ _2219_ _1699_ VGND VGND VPWR VPWR _2220_ sky130_fd_sc_hd__mux2_1
X_7203_ _3544_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4415_ _1170_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__buf_6
XFILLER_0_1_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5395_ _2147_ _2150_ net4 VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__mux2_1
X_8183_ _4065_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__clkbuf_1
X_7134_ _3507_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
X_4346_ _1071_ _1101_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__nand2_1
X_4277_ RF.registers\[24\]\[4\] RF.registers\[25\]\[4\] RF.registers\[26\]\[4\] RF.registers\[27\]\[4\]
+ _1027_ _1029_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__mux4_1
X_7065_ RF.registers\[19\]\[2\] _3460_ _3456_ VGND VGND VPWR VPWR _3461_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6016_ _2496_ _2754_ VGND VGND VPWR VPWR _2755_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7967_ RF.registers\[18\]\[31\] _3452_ _3915_ VGND VGND VPWR VPWR _3950_ sky130_fd_sc_hd__mux2_1
X_7898_ _3913_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__clkbuf_1
X_6918_ _3378_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6849_ RF.registers\[5\]\[1\] _3095_ _3340_ VGND VGND VPWR VPWR _3342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_666 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9568_ clknet_leaf_72_CLK _0728_ VGND VGND VPWR VPWR RF.registers\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9499_ clknet_leaf_46_CLK _0659_ VGND VGND VPWR VPWR RF.registers\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_114_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8519_ _4242_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5180_ RF.registers\[0\]\[29\] RF.registers\[1\]\[29\] RF.registers\[2\]\[29\] RF.registers\[3\]\[29\]
+ _1895_ _1897_ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_8870_ clknet_leaf_61_CLK _0030_ VGND VGND VPWR VPWR RF.registers\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7821_ RF.registers\[9\]\[26\] _3442_ _3866_ VGND VGND VPWR VPWR _3873_ sky130_fd_sc_hd__mux2_1
X_7752_ _3836_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_82_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4964_ _1719_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6703_ _3263_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7683_ RF.registers\[2\]\[25\] _3508_ _3794_ VGND VGND VPWR VPWR _3800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9422_ clknet_leaf_39_CLK _0582_ VGND VGND VPWR VPWR RF.registers\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4895_ RF.registers\[8\]\[0\] RF.registers\[9\]\[0\] RF.registers\[10\]\[0\] RF.registers\[11\]\[0\]
+ _1641_ _1642_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_22_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6634_ _3083_ RF.registers\[15\]\[29\] _3217_ VGND VGND VPWR VPWR _3227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6565_ _3189_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9353_ clknet_leaf_87_CLK _0513_ VGND VGND VPWR VPWR RF.registers\[20\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8304_ _3013_ RF.registers\[13\]\[29\] _4119_ VGND VGND VPWR VPWR _4129_ sky130_fd_sc_hd__mux2_1
X_6496_ _3151_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__clkbuf_1
X_5516_ _1638_ _2271_ VGND VGND VPWR VPWR _2272_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9284_ clknet_leaf_95_CLK _0444_ VGND VGND VPWR VPWR RF.registers\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_8235_ _4092_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__clkbuf_1
X_5447_ RF.registers\[12\]\[10\] RF.registers\[13\]\[10\] RF.registers\[14\]\[10\]
+ RF.registers\[15\]\[10\] _2117_ _2118_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8166_ RF.registers\[24\]\[28\] _3446_ _4047_ VGND VGND VPWR VPWR _4056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5378_ _2132_ _2133_ _1711_ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__mux2_1
X_8097_ _4019_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__clkbuf_1
X_7117_ RF.registers\[19\]\[19\] _3495_ _3477_ VGND VGND VPWR VPWR _3496_ sky130_fd_sc_hd__mux2_1
X_4329_ net47 _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7048_ RF.registers\[3\]\[29\] _3448_ _3435_ VGND VGND VPWR VPWR _3449_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8999_ clknet_leaf_58_CLK _0159_ VGND VGND VPWR VPWR RF.registers\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4680_ _1434_ _1435_ _1178_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6350_ _3053_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5301_ _1828_ _2056_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6281_ net9 _3004_ VGND VGND VPWR VPWR _3005_ sky130_fd_sc_hd__or2_4
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8020_ _3978_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__clkbuf_1
X_5232_ RF.registers\[12\]\[26\] RF.registers\[13\]\[26\] RF.registers\[14\]\[26\]
+ RF.registers\[15\]\[26\] _1896_ _1898_ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5163_ _1823_ VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5094_ RF.registers\[8\]\[17\] RF.registers\[9\]\[17\] RF.registers\[10\]\[17\] RF.registers\[11\]\[17\]
+ _1720_ _1723_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__mux4_1
X_8922_ clknet_leaf_24_CLK _0082_ VGND VGND VPWR VPWR RF.registers\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8853_ clknet_leaf_53_CLK _0013_ VGND VGND VPWR VPWR RF.registers\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7804_ RF.registers\[9\]\[18\] _3493_ _3855_ VGND VGND VPWR VPWR _3864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5996_ _2733_ _2735_ _1879_ VGND VGND VPWR VPWR _2736_ sky130_fd_sc_hd__mux2_1
X_8784_ clknet_leaf_58_CLK _0968_ VGND VGND VPWR VPWR RF.registers\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7735_ _3827_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__clkbuf_1
X_4947_ _1702_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7666_ RF.registers\[2\]\[17\] _3491_ _3783_ VGND VGND VPWR VPWR _3791_ sky130_fd_sc_hd__mux2_1
X_4878_ _1239_ _1625_ _1629_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_62_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6617_ _3218_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__clkbuf_1
X_9405_ clknet_leaf_18_CLK _0565_ VGND VGND VPWR VPWR RF.registers\[24\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9336_ clknet_leaf_39_CLK _0496_ VGND VGND VPWR VPWR RF.registers\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_7597_ _3754_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6548_ RF.registers\[0\]\[21\] _3137_ _3179_ VGND VGND VPWR VPWR _3181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9267_ clknet_leaf_30_CLK _0427_ VGND VGND VPWR VPWR RF.registers\[23\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_6479_ RF.registers\[17\]\[23\] _3141_ _3135_ VGND VGND VPWR VPWR _3142_ sky130_fd_sc_hd__mux2_1
X_8218_ RF.registers\[1\]\[20\] _3497_ _4083_ VGND VGND VPWR VPWR _4084_ sky130_fd_sc_hd__mux2_1
X_9198_ clknet_leaf_20_CLK _0358_ VGND VGND VPWR VPWR RF.registers\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8149_ _4024_ VGND VGND VPWR VPWR _4047_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_122_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5850_ _2229_ _2597_ VGND VGND VPWR VPWR _2598_ sky130_fd_sc_hd__xor2_2
XFILLER_0_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5781_ _2255_ _2355_ _2364_ _2337_ VGND VGND VPWR VPWR _2532_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4801_ _1088_ _1556_ net8 VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4732_ RF.registers\[0\]\[14\] RF.registers\[1\]\[14\] RF.registers\[2\]\[14\] RF.registers\[3\]\[14\]
+ _1191_ _1174_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__mux4_1
X_7520_ _3048_ RF.registers\[27\]\[12\] _3711_ VGND VGND VPWR VPWR _3714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4663_ RF.registers\[16\]\[23\] RF.registers\[17\]\[23\] RF.registers\[18\]\[23\]
+ RF.registers\[19\]\[23\] _1351_ _1352_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7451_ _3677_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6402_ _3088_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4594_ _1238_ _1278_ _1316_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7382_ _3046_ RF.registers\[26\]\[11\] _3639_ VGND VGND VPWR VPWR _3641_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6333_ _3041_ RF.registers\[22\]\[9\] _3023_ VGND VGND VPWR VPWR _3042_ sky130_fd_sc_hd__mux2_1
X_9121_ clknet_leaf_96_CLK _0281_ VGND VGND VPWR VPWR RF.registers\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_6264_ _2988_ _2989_ VGND VGND VPWR VPWR _2990_ sky130_fd_sc_hd__nor2_1
X_9052_ clknet_leaf_22_CLK _0212_ VGND VGND VPWR VPWR RF.registers\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5215_ RF.registers\[12\]\[27\] RF.registers\[13\]\[27\] RF.registers\[14\]\[27\]
+ RF.registers\[15\]\[27\] _1918_ _1919_ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_90_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8003_ _3969_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__clkbuf_1
X_6195_ _2923_ _2384_ VGND VGND VPWR VPWR _2924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5146_ _1899_ _1900_ _1901_ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__mux2_1
X_5077_ _1700_ _1832_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__nand2_1
X_8905_ clknet_leaf_9_CLK _0065_ VGND VGND VPWR VPWR RF.registers\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8836_ clknet_leaf_78_CLK _1020_ VGND VGND VPWR VPWR RF.registers\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_5979_ _2569_ _2719_ _2104_ VGND VGND VPWR VPWR _2720_ sky130_fd_sc_hd__mux2_1
X_8767_ clknet_leaf_65_CLK _0951_ VGND VGND VPWR VPWR RF.registers\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7718_ _3818_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8698_ clknet_leaf_36_CLK _0882_ VGND VGND VPWR VPWR RF.registers\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7649_ RF.registers\[2\]\[9\] _3474_ _3772_ VGND VGND VPWR VPWR _3782_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9319_ clknet_leaf_58_CLK _0479_ VGND VGND VPWR VPWR RF.registers\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _1668_ _1755_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_72_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6951_ _3395_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_37_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5902_ _2644_ _2646_ VGND VGND VPWR VPWR _2647_ sky130_fd_sc_hd__xnor2_1
X_6882_ RF.registers\[5\]\[17\] _3128_ _3351_ VGND VGND VPWR VPWR _3359_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5833_ _2230_ _2580_ _1839_ VGND VGND VPWR VPWR _2581_ sky130_fd_sc_hd__mux2_1
X_8621_ clknet_leaf_6_CLK _0805_ VGND VGND VPWR VPWR RF.registers\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8552_ RF.registers\[10\]\[18\] net23 _4255_ VGND VGND VPWR VPWR _4260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5764_ _1083_ _2514_ VGND VGND VPWR VPWR _2515_ sky130_fd_sc_hd__xnor2_1
X_7503_ _3031_ RF.registers\[27\]\[4\] _3700_ VGND VGND VPWR VPWR _3705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8483_ RF.registers\[11\]\[17\] net22 _4216_ VGND VGND VPWR VPWR _4224_ sky130_fd_sc_hd__mux2_1
X_5695_ _2080_ _2448_ VGND VGND VPWR VPWR _2449_ sky130_fd_sc_hd__xor2_1
X_4715_ _1467_ _1470_ _1071_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__mux2_1
X_7434_ _3668_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4646_ _1400_ _1401_ _1107_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4577_ _1327_ _1329_ _1332_ _1187_ _1215_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7365_ _3029_ RF.registers\[26\]\[3\] _3628_ VGND VGND VPWR VPWR _3632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9104_ clknet_leaf_6_CLK _0264_ VGND VGND VPWR VPWR RF.registers\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6316_ _3030_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_3__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_3_3__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7296_ _3029_ RF.registers\[31\]\[3\] _3591_ VGND VGND VPWR VPWR _3595_ sky130_fd_sc_hd__mux2_1
X_6247_ _2972_ VGND VGND VPWR VPWR _2973_ sky130_fd_sc_hd__inv_2
X_9035_ clknet_leaf_98_CLK _0195_ VGND VGND VPWR VPWR RF.registers\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_6178_ _2444_ _2864_ VGND VGND VPWR VPWR _2908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5129_ RF.registers\[24\]\[31\] RF.registers\[25\]\[31\] RF.registers\[26\]\[31\]
+ RF.registers\[27\]\[31\] _1882_ _1884_ VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8819_ clknet_leaf_51_CLK _1003_ VGND VGND VPWR VPWR RF.registers\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4500_ _1239_ _1246_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__o21ai_2
X_5480_ _2234_ _2235_ _1685_ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 _1421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4431_ _1071_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7150_ _3411_ _3302_ VGND VGND VPWR VPWR _3516_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4362_ _1107_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__or2_1
X_6101_ _1256_ _1277_ VGND VGND VPWR VPWR _2835_ sky130_fd_sc_hd__and2_1
X_4293_ RF.registers\[0\]\[4\] RF.registers\[1\]\[4\] RF.registers\[2\]\[4\] RF.registers\[3\]\[4\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7081_ _3471_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
X_6032_ _2744_ _2763_ VGND VGND VPWR VPWR _2770_ sky130_fd_sc_hd__nand2_1
X_7983_ _3105_ RF.registers\[21\]\[6\] _3952_ VGND VGND VPWR VPWR _3959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6934_ _3386_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8604_ clknet_leaf_18_CLK _0788_ VGND VGND VPWR VPWR RF.registers\[22\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_6865_ RF.registers\[5\]\[9\] _3111_ _3340_ VGND VGND VPWR VPWR _3350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_9584_ clknet_leaf_12_CLK _0744_ VGND VGND VPWR VPWR RF.registers\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_5816_ _2361_ _2357_ VGND VGND VPWR VPWR _2565_ sky130_fd_sc_hd__and2_1
X_6796_ _3313_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5747_ _2498_ VGND VGND VPWR VPWR _2499_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8535_ RF.registers\[10\]\[10\] net15 _4244_ VGND VGND VPWR VPWR _4251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8466_ RF.registers\[11\]\[9\] net45 _4205_ VGND VGND VPWR VPWR _4215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7417_ _3081_ RF.registers\[26\]\[28\] _3650_ VGND VGND VPWR VPWR _3659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5678_ _2083_ VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__inv_2
X_4629_ _1370_ _1384_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__nand2_1
X_8397_ _4178_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_50_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_50_CLK sky130_fd_sc_hd__clkbuf_8
X_7348_ _3081_ RF.registers\[31\]\[28\] _3613_ VGND VGND VPWR VPWR _3622_ sky130_fd_sc_hd__mux2_1
X_7279_ _3585_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9018_ clknet_leaf_25_CLK _0178_ VGND VGND VPWR VPWR RF.registers\[31\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_41_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_41_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_56_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput60 net60 VGND VGND VPWR VPWR ALU_result[1] sky130_fd_sc_hd__buf_1
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput71 net71 VGND VGND VPWR VPWR ALU_result[2] sky130_fd_sc_hd__buf_1
XFILLER_0_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4980_ RF.registers\[20\]\[22\] RF.registers\[21\]\[22\] RF.registers\[22\]\[22\]
+ RF.registers\[23\]\[22\] _1734_ _1735_ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_47_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6650_ RF.registers\[8\]\[4\] _3101_ _3231_ VGND VGND VPWR VPWR _3236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5601_ _2348_ _2355_ _1879_ VGND VGND VPWR VPWR _2356_ sky130_fd_sc_hd__mux2_1
X_6581_ _3199_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__clkbuf_1
X_5532_ _1800_ _2287_ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8320_ RF.registers\[16\]\[4\] _3464_ _4133_ VGND VGND VPWR VPWR _4138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8251_ _4101_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__clkbuf_1
X_5463_ _2217_ _2218_ _1685_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_32_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_32_CLK sky130_fd_sc_hd__clkbuf_8
X_7202_ RF.registers\[7\]\[24\] _3506_ _3539_ VGND VGND VPWR VPWR _3544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4414_ _1057_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__buf_4
X_5394_ _2148_ _2149_ _1684_ VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__mux2_1
X_8182_ RF.registers\[1\]\[3\] _3462_ _4061_ VGND VGND VPWR VPWR _4065_ sky130_fd_sc_hd__mux2_1
X_7133_ RF.registers\[19\]\[24\] _3506_ _3498_ VGND VGND VPWR VPWR _3507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4345_ _1099_ _1100_ _1048_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4276_ RF.registers\[28\]\[4\] RF.registers\[29\]\[4\] RF.registers\[30\]\[4\] RF.registers\[31\]\[4\]
+ _1027_ _1029_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__mux4_1
X_7064_ net36 VGND VGND VPWR VPWR _3460_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_129_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6015_ _2751_ _2753_ _2252_ VGND VGND VPWR VPWR _2754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7966_ _3949_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7897_ _3015_ RF.registers\[23\]\[30\] _3879_ VGND VGND VPWR VPWR _3913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6917_ RF.registers\[4\]\[1\] _3095_ _3376_ VGND VGND VPWR VPWR _3378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6848_ _3341_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9567_ clknet_leaf_64_CLK _0727_ VGND VGND VPWR VPWR RF.registers\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_138_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8518_ RF.registers\[10\]\[2\] net36 _3007_ VGND VGND VPWR VPWR _4242_ sky130_fd_sc_hd__mux2_1
X_6779_ RF.registers\[6\]\[0\] _3089_ _3304_ VGND VGND VPWR VPWR _3305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9498_ clknet_leaf_28_CLK _0658_ VGND VGND VPWR VPWR RF.registers\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_98_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8449_ _4206_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_23_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_14_CLK clknet_3_4__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_14_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7820_ _3872_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7751_ _3075_ RF.registers\[30\]\[25\] _3830_ VGND VGND VPWR VPWR _3836_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4963_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__clkbuf_8
X_7682_ _3799_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__clkbuf_1
X_6702_ RF.registers\[8\]\[29\] _3013_ _3253_ VGND VGND VPWR VPWR _3263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6633_ _3226_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__clkbuf_1
X_9421_ clknet_leaf_83_CLK _0581_ VGND VGND VPWR VPWR RF.registers\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_4894_ _1646_ _1649_ net4 VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6564_ RF.registers\[0\]\[29\] _3013_ _3179_ VGND VGND VPWR VPWR _3189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9352_ clknet_leaf_88_CLK _0512_ VGND VGND VPWR VPWR RF.registers\[20\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8303_ _4128_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__clkbuf_1
X_6495_ RF.registers\[17\]\[30\] _3015_ _3092_ VGND VGND VPWR VPWR _3151_ sky130_fd_sc_hd__mux2_1
X_9283_ clknet_leaf_76_CLK _0443_ VGND VGND VPWR VPWR RF.registers\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_5515_ _1670_ _2262_ _2266_ _2270_ VGND VGND VPWR VPWR _2271_ sky130_fd_sc_hd__a2bb2o_2
X_8234_ RF.registers\[1\]\[28\] _3446_ _4083_ VGND VGND VPWR VPWR _4092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5446_ RF.registers\[8\]\[10\] RF.registers\[9\]\[10\] RF.registers\[10\]\[10\] RF.registers\[11\]\[10\]
+ _1703_ _1706_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8165_ _4055_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5377_ RF.registers\[12\]\[14\] RF.registers\[13\]\[14\] RF.registers\[14\]\[14\]
+ RF.registers\[15\]\[14\] _2113_ _2114_ VGND VGND VPWR VPWR _2133_ sky130_fd_sc_hd__mux4_1
X_8096_ RF.registers\[20\]\[27\] _3444_ _4011_ VGND VGND VPWR VPWR _4019_ sky130_fd_sc_hd__mux2_1
X_7116_ net24 VGND VGND VPWR VPWR _3495_ sky130_fd_sc_hd__clkbuf_4
X_4328_ net48 _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__nand2_1
X_7047_ net35 VGND VGND VPWR VPWR _3448_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_2_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8998_ clknet_leaf_65_CLK _0158_ VGND VGND VPWR VPWR RF.registers\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_7949_ RF.registers\[18\]\[22\] _3502_ _3938_ VGND VGND VPWR VPWR _3941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_CLK clknet_3_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_3_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5300_ _2054_ _2055_ _1712_ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6280_ net10 net46 VGND VGND VPWR VPWR _3004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5231_ _1983_ _1986_ _1766_ VGND VGND VPWR VPWR _1987_ sky130_fd_sc_hd__mux2_1
X_5162_ _1822_ VGND VGND VPWR VPWR _1918_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5093_ _1845_ _1848_ _1697_ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__mux2_1
X_8921_ clknet_leaf_27_CLK _0081_ VGND VGND VPWR VPWR RF.registers\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8852_ clknet_leaf_53_CLK _0012_ VGND VGND VPWR VPWR RF.registers\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7803_ _3863_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__clkbuf_1
X_8783_ clknet_leaf_84_CLK _0967_ VGND VGND VPWR VPWR RF.registers\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5995_ _2703_ _2734_ _2347_ VGND VGND VPWR VPWR _2735_ sky130_fd_sc_hd__mux2_1
X_7734_ _3058_ RF.registers\[30\]\[17\] _3819_ VGND VGND VPWR VPWR _3827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4946_ _1701_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__buf_4
X_7665_ _3790_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
X_4877_ _1254_ _1632_ _1170_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6616_ _3064_ RF.registers\[15\]\[20\] _3217_ VGND VGND VPWR VPWR _3218_ sky130_fd_sc_hd__mux2_1
X_9404_ clknet_leaf_23_CLK _0564_ VGND VGND VPWR VPWR RF.registers\[24\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_7596_ _3056_ RF.registers\[28\]\[16\] _3747_ VGND VGND VPWR VPWR _3754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9335_ clknet_leaf_32_CLK _0495_ VGND VGND VPWR VPWR RF.registers\[21\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6547_ _3180_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6478_ net29 VGND VGND VPWR VPWR _3141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9266_ clknet_leaf_40_CLK _0426_ VGND VGND VPWR VPWR RF.registers\[23\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_8217_ _4060_ VGND VGND VPWR VPWR _4083_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_7_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5429_ RF.registers\[12\]\[11\] RF.registers\[13\]\[11\] RF.registers\[14\]\[11\]
+ RF.registers\[15\]\[11\] _1704_ _1707_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__mux4_1
X_9197_ clknet_leaf_3_CLK _0357_ VGND VGND VPWR VPWR RF.registers\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_8148_ _4046_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8079_ RF.registers\[20\]\[19\] _3495_ _4000_ VGND VGND VPWR VPWR _4010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4800_ _1554_ _1555_ _1107_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5780_ _2403_ _2348_ _1879_ VGND VGND VPWR VPWR _2531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4731_ _1198_ _1486_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4662_ RF.registers\[28\]\[23\] RF.registers\[29\]\[23\] RF.registers\[30\]\[23\]
+ RF.registers\[31\]\[23\] _1267_ _1268_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7450_ _3046_ RF.registers\[25\]\[11\] _3675_ VGND VGND VPWR VPWR _3677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6401_ _3087_ RF.registers\[22\]\[31\] _3022_ VGND VGND VPWR VPWR _3088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4593_ _1334_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__or2b_1
X_9120_ clknet_leaf_69_CLK _0280_ VGND VGND VPWR VPWR RF.registers\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7381_ _3640_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6332_ net45 VGND VGND VPWR VPWR _3041_ sky130_fd_sc_hd__clkbuf_2
X_9051_ clknet_leaf_35_CLK _0211_ VGND VGND VPWR VPWR RF.registers\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6263_ _2952_ _2987_ _2986_ VGND VGND VPWR VPWR _2989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5214_ RF.registers\[8\]\[27\] RF.registers\[9\]\[27\] RF.registers\[10\]\[27\] RF.registers\[11\]\[27\]
+ _1918_ _1919_ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8002_ _3124_ RF.registers\[21\]\[15\] _3963_ VGND VGND VPWR VPWR _3969_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6194_ _1669_ _1997_ VGND VGND VPWR VPWR _2923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5145_ _1726_ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5076_ _1830_ _1831_ _1686_ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8904_ clknet_leaf_1_CLK _0064_ VGND VGND VPWR VPWR RF.registers\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8835_ clknet_leaf_73_CLK _1019_ VGND VGND VPWR VPWR RF.registers\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5978_ _2650_ _2718_ _2251_ VGND VGND VPWR VPWR _2719_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8766_ clknet_leaf_67_CLK _0950_ VGND VGND VPWR VPWR RF.registers\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_8697_ clknet_leaf_31_CLK _0881_ VGND VGND VPWR VPWR RF.registers\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7717_ _3041_ RF.registers\[30\]\[9\] _3808_ VGND VGND VPWR VPWR _3818_ sky130_fd_sc_hd__mux2_1
X_4929_ _1684_ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7648_ _3781_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_119_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7579_ _3039_ RF.registers\[28\]\[8\] _3736_ VGND VGND VPWR VPWR _3745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9318_ clknet_leaf_61_CLK _0478_ VGND VGND VPWR VPWR RF.registers\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9249_ clknet_leaf_93_CLK _0409_ VGND VGND VPWR VPWR RF.registers\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_773 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6950_ RF.registers\[4\]\[17\] _3128_ _3387_ VGND VGND VPWR VPWR _3395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5901_ _2633_ _2636_ _2645_ VGND VGND VPWR VPWR _2646_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_37_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6881_ _3358_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5832_ _2287_ VGND VGND VPWR VPWR _2580_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8620_ clknet_leaf_3_CLK _0804_ VGND VGND VPWR VPWR RF.registers\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_8551_ _4259_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5763_ _1060_ _2506_ _2411_ VGND VGND VPWR VPWR _2514_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7502_ _3704_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
X_4714_ _1468_ _1469_ _1036_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8482_ _4223_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__clkbuf_1
X_5694_ _1125_ _2447_ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7433_ _3029_ RF.registers\[25\]\[3\] _3664_ VGND VGND VPWR VPWR _3668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4645_ RF.registers\[16\]\[7\] RF.registers\[17\]\[7\] RF.registers\[18\]\[7\] RF.registers\[19\]\[7\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__mux4_1
X_4576_ _1330_ _1331_ _1259_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__mux2_1
X_7364_ _3631_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9103_ clknet_leaf_5_CLK _0263_ VGND VGND VPWR VPWR RF.registers\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6315_ _3029_ RF.registers\[22\]\[3\] _3023_ VGND VGND VPWR VPWR _3030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7295_ _3594_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_9034_ clknet_leaf_8_CLK _0194_ VGND VGND VPWR VPWR RF.registers\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_6246_ _2970_ _2971_ _1126_ VGND VGND VPWR VPWR _2972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_110_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6177_ _2626_ _2797_ VGND VGND VPWR VPWR _2907_ sky130_fd_sc_hd__nor2_1
X_5128_ _1883_ VGND VGND VPWR VPWR _1884_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5059_ _1700_ _1814_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__nand2_1
X_8818_ clknet_leaf_54_CLK _1002_ VGND VGND VPWR VPWR RF.registers\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8749_ clknet_leaf_10_CLK _0933_ VGND VGND VPWR VPWR RF.registers\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_762 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4430_ _1180_ _1185_ _1178_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__mux2_1
XANTENNA_2 _1471_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6100_ _2496_ _2822_ _2826_ _2834_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__a211o_1
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4361_ RF.registers\[4\]\[2\] RF.registers\[5\]\[2\] RF.registers\[6\]\[2\] RF.registers\[7\]\[2\]
+ _1065_ _1066_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4292_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__buf_4
X_7080_ RF.registers\[19\]\[7\] _3470_ _3456_ VGND VGND VPWR VPWR _3471_ sky130_fd_sc_hd__mux2_1
X_6031_ _1820_ _2768_ VGND VGND VPWR VPWR _2769_ sky130_fd_sc_hd__xnor2_1
X_7982_ _3958_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__clkbuf_1
X_6933_ RF.registers\[4\]\[9\] _3111_ _3376_ VGND VGND VPWR VPWR _3386_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6864_ _3349_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8603_ clknet_leaf_46_CLK _0787_ VGND VGND VPWR VPWR RF.registers\[22\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5815_ _2561_ _2563_ VGND VGND VPWR VPWR _2564_ sky130_fd_sc_hd__xnor2_1
X_9583_ clknet_leaf_11_CLK _0743_ VGND VGND VPWR VPWR RF.registers\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_6795_ RF.registers\[6\]\[8\] _3109_ _3304_ VGND VGND VPWR VPWR _3313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5746_ _2064_ _2307_ VGND VGND VPWR VPWR _2498_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8534_ _4250_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5677_ _2430_ _2289_ _2363_ VGND VGND VPWR VPWR _2431_ sky130_fd_sc_hd__mux2_1
X_8465_ _4214_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4628_ _1171_ _1375_ _1379_ _1383_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__o2bb2a_2
X_7416_ _3658_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_116_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8396_ RF.registers\[12\]\[8\] _3472_ _4169_ VGND VGND VPWR VPWR _4178_ sky130_fd_sc_hd__mux2_1
X_7347_ _3621_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
X_4559_ _1171_ _1306_ _1310_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__o2bb2a_1
X_7278_ _3079_ RF.registers\[29\]\[27\] _3577_ VGND VGND VPWR VPWR _3585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9017_ clknet_leaf_26_CLK _0177_ VGND VGND VPWR VPWR RF.registers\[31\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6229_ _2953_ _2954_ VGND VGND VPWR VPWR _2956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput61 net61 VGND VGND VPWR VPWR ALU_result[20] sky130_fd_sc_hd__buf_1
Xoutput50 net50 VGND VGND VPWR VPWR ALU_result[10] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_56_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput72 net72 VGND VGND VPWR VPWR ALU_result[30] sky130_fd_sc_hd__buf_1
XFILLER_0_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5600_ _2351_ _2354_ _2347_ VGND VGND VPWR VPWR _2355_ sky130_fd_sc_hd__mux2_1
X_6580_ _3029_ RF.registers\[15\]\[3\] _3195_ VGND VGND VPWR VPWR _3199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5531_ _1638_ _2286_ VGND VGND VPWR VPWR _2287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8250_ _3099_ RF.registers\[13\]\[3\] _4097_ VGND VGND VPWR VPWR _4101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7201_ _3543_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5462_ RF.registers\[24\]\[8\] RF.registers\[25\]\[8\] RF.registers\[26\]\[8\] RF.registers\[27\]\[8\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4413_ _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8181_ _4064_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__clkbuf_1
X_5393_ RF.registers\[24\]\[13\] RF.registers\[25\]\[13\] RF.registers\[26\]\[13\]
+ RF.registers\[27\]\[13\] _1673_ _1690_ VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__mux4_1
X_7132_ net30 VGND VGND VPWR VPWR _3506_ sky130_fd_sc_hd__buf_2
X_4344_ RF.registers\[12\]\[3\] RF.registers\[13\]\[3\] RF.registers\[14\]\[3\] RF.registers\[15\]\[3\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7063_ _3459_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6014_ _2717_ _2752_ _1146_ VGND VGND VPWR VPWR _2753_ sky130_fd_sc_hd__mux2_1
X_4275_ RF.registers\[16\]\[4\] RF.registers\[17\]\[4\] RF.registers\[18\]\[4\] RF.registers\[19\]\[4\]
+ _1027_ _1029_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7965_ RF.registers\[18\]\[30\] _3450_ _3915_ VGND VGND VPWR VPWR _3949_ sky130_fd_sc_hd__mux2_1
X_7896_ _3912_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6916_ _3377_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6847_ RF.registers\[5\]\[0\] _3089_ _3340_ VGND VGND VPWR VPWR _3341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6778_ _3303_ VGND VGND VPWR VPWR _3304_ sky130_fd_sc_hd__clkbuf_8
X_9566_ clknet_leaf_71_CLK _0726_ VGND VGND VPWR VPWR RF.registers\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_5729_ _2480_ _2481_ VGND VGND VPWR VPWR _2482_ sky130_fd_sc_hd__or2b_1
X_8517_ _4241_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__clkbuf_1
X_9497_ clknet_leaf_30_CLK _0657_ VGND VGND VPWR VPWR RF.registers\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_98_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8448_ RF.registers\[11\]\[0\] net14 _4205_ VGND VGND VPWR VPWR _4206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8379_ _4168_ VGND VGND VPWR VPWR _4169_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7750_ _3835_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_82_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4962_ _1702_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__buf_4
X_7681_ RF.registers\[2\]\[24\] _3506_ _3794_ VGND VGND VPWR VPWR _3799_ sky130_fd_sc_hd__mux2_1
X_6701_ _3262_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4893_ _1647_ _1648_ _1645_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__mux2_1
X_6632_ _3081_ RF.registers\[15\]\[28\] _3217_ VGND VGND VPWR VPWR _3226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9420_ clknet_leaf_84_CLK _0580_ VGND VGND VPWR VPWR RF.registers\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6563_ _3188_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__clkbuf_1
X_9351_ clknet_leaf_59_CLK _0511_ VGND VGND VPWR VPWR RF.registers\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6494_ _3150_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__clkbuf_1
X_8302_ _3011_ RF.registers\[13\]\[28\] _4119_ VGND VGND VPWR VPWR _4128_ sky130_fd_sc_hd__mux2_1
X_9282_ clknet_leaf_92_CLK _0442_ VGND VGND VPWR VPWR RF.registers\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_5514_ _1828_ _2269_ _1728_ VGND VGND VPWR VPWR _2270_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8233_ _4091_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5445_ _2197_ _2200_ _1716_ VGND VGND VPWR VPWR _2201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8164_ RF.registers\[24\]\[27\] _3444_ _4047_ VGND VGND VPWR VPWR _4055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7115_ _3494_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
X_5376_ RF.registers\[8\]\[14\] RF.registers\[9\]\[14\] RF.registers\[10\]\[14\] RF.registers\[11\]\[14\]
+ _2113_ _2114_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__mux4_1
X_8095_ _4018_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__clkbuf_1
X_4327_ _1025_ _1070_ _1077_ _1082_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7046_ _3447_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8997_ clknet_leaf_80_CLK _0157_ VGND VGND VPWR VPWR RF.registers\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_7948_ _3940_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7879_ _3137_ RF.registers\[23\]\[21\] _3902_ VGND VGND VPWR VPWR _3904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_9549_ clknet_leaf_11_CLK _0709_ VGND VGND VPWR VPWR RF.registers\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5230_ _1984_ _1985_ _1901_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__mux2_1
X_5161_ RF.registers\[4\]\[30\] RF.registers\[5\]\[30\] RF.registers\[6\]\[30\] RF.registers\[7\]\[30\]
+ _1881_ _1883_ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5092_ _1846_ _1847_ _1686_ VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__mux2_1
X_8920_ clknet_leaf_38_CLK _0080_ VGND VGND VPWR VPWR RF.registers\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8851_ clknet_leaf_50_CLK _0011_ VGND VGND VPWR VPWR RF.registers\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5994_ _1169_ _2124_ _1875_ VGND VGND VPWR VPWR _2734_ sky130_fd_sc_hd__o21a_1
X_8782_ clknet_leaf_40_CLK _0966_ VGND VGND VPWR VPWR RF.registers\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7802_ RF.registers\[9\]\[17\] _3491_ _3855_ VGND VGND VPWR VPWR _3863_ sky130_fd_sc_hd__mux2_1
X_7733_ _3826_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__clkbuf_1
X_4945_ net1 VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7664_ RF.registers\[2\]\[16\] _3489_ _3783_ VGND VGND VPWR VPWR _3790_ sky130_fd_sc_hd__mux2_1
X_4876_ _1630_ _1631_ _1178_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__mux2_1
X_9403_ clknet_leaf_46_CLK _0563_ VGND VGND VPWR VPWR RF.registers\[24\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_6615_ _3194_ VGND VGND VPWR VPWR _3217_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7595_ _3753_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
X_9334_ clknet_leaf_48_CLK _0494_ VGND VGND VPWR VPWR RF.registers\[21\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6546_ RF.registers\[0\]\[20\] _3134_ _3179_ VGND VGND VPWR VPWR _3180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6477_ _3140_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__clkbuf_1
X_9265_ clknet_leaf_19_CLK _0425_ VGND VGND VPWR VPWR RF.registers\[23\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_8216_ _4082_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9196_ clknet_leaf_2_CLK _0356_ VGND VGND VPWR VPWR RF.registers\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_5428_ _2180_ _2181_ _2182_ _2183_ _1712_ _1716_ VGND VGND VPWR VPWR _2184_ sky130_fd_sc_hd__mux4_1
X_8147_ RF.registers\[24\]\[19\] _3495_ _4036_ VGND VGND VPWR VPWR _4046_ sky130_fd_sc_hd__mux2_1
X_5359_ RF.registers\[12\]\[15\] RF.registers\[13\]\[15\] RF.registers\[14\]\[15\]
+ RF.registers\[15\]\[15\] _2113_ _2114_ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__mux4_1
X_8078_ _4009_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7029_ _3437_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4730_ RF.registers\[4\]\[14\] RF.registers\[5\]\[14\] RF.registers\[6\]\[14\] RF.registers\[7\]\[14\]
+ _1172_ _1279_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4661_ RF.registers\[24\]\[23\] RF.registers\[25\]\[23\] RF.registers\[26\]\[23\]
+ RF.registers\[27\]\[23\] _1351_ _1352_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6400_ net38 VGND VGND VPWR VPWR _3087_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7380_ _3043_ RF.registers\[26\]\[10\] _3639_ VGND VGND VPWR VPWR _3640_ sky130_fd_sc_hd__mux2_1
X_4592_ _1171_ _1339_ _1347_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_12_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6331_ _3040_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9050_ clknet_leaf_25_CLK _0210_ VGND VGND VPWR VPWR RF.registers\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_6262_ _2952_ _2986_ _2987_ VGND VGND VPWR VPWR _2988_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5213_ _1965_ _1968_ _1700_ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6193_ _2254_ _2858_ VGND VGND VPWR VPWR _2922_ sky130_fd_sc_hd__or2_1
X_8001_ _3968_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5144_ RF.registers\[0\]\[31\] RF.registers\[1\]\[31\] RF.registers\[2\]\[31\] RF.registers\[3\]\[31\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5075_ RF.registers\[8\]\[19\] RF.registers\[9\]\[19\] RF.registers\[10\]\[19\] RF.registers\[11\]\[19\]
+ _1689_ _1693_ VGND VGND VPWR VPWR _1831_ sky130_fd_sc_hd__mux4_1
X_8903_ clknet_leaf_83_CLK _0063_ VGND VGND VPWR VPWR RF.registers\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8834_ clknet_leaf_76_CLK _1018_ VGND VGND VPWR VPWR RF.registers\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_32_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8765_ clknet_leaf_18_CLK _0949_ VGND VGND VPWR VPWR RF.registers\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_5977_ _2697_ _2717_ _1803_ VGND VGND VPWR VPWR _2718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8696_ clknet_leaf_38_CLK _0880_ VGND VGND VPWR VPWR RF.registers\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_4928_ _1645_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__buf_4
X_7716_ _3817_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7647_ RF.registers\[2\]\[8\] _3472_ _3772_ VGND VGND VPWR VPWR _3781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4859_ RF.registers\[12\]\[19\] RF.registers\[13\]\[19\] RF.registers\[14\]\[19\]
+ RF.registers\[15\]\[19\] _1173_ _1175_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7578_ _3744_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9317_ clknet_leaf_63_CLK _0477_ VGND VGND VPWR VPWR RF.registers\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_6529_ RF.registers\[0\]\[12\] _3118_ _3168_ VGND VGND VPWR VPWR _3171_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9248_ clknet_leaf_73_CLK _0408_ VGND VGND VPWR VPWR RF.registers\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9179_ clknet_leaf_44_CLK _0339_ VGND VGND VPWR VPWR RF.registers\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5900_ _2210_ _2632_ VGND VGND VPWR VPWR _2645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6880_ RF.registers\[5\]\[16\] _3126_ _3351_ VGND VGND VPWR VPWR _3358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5831_ _2578_ VGND VGND VPWR VPWR _2579_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8550_ RF.registers\[10\]\[17\] net22 _4255_ VGND VGND VPWR VPWR _4259_ sky130_fd_sc_hd__mux2_1
X_5762_ _2489_ _2494_ _2505_ _2513_ _2408_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__o32a_1
XFILLER_0_57_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7501_ _3029_ RF.registers\[27\]\[3\] _3700_ VGND VGND VPWR VPWR _3704_ sky130_fd_sc_hd__mux2_1
X_4713_ RF.registers\[24\]\[13\] RF.registers\[25\]\[13\] RF.registers\[26\]\[13\]
+ RF.registers\[27\]\[13\] _1027_ _1029_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8481_ RF.registers\[11\]\[16\] net21 _4216_ VGND VGND VPWR VPWR _4223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5693_ _1145_ _1166_ _2411_ VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7432_ _3667_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__clkbuf_1
X_4644_ RF.registers\[20\]\[7\] RF.registers\[21\]\[7\] RF.registers\[22\]\[7\] RF.registers\[23\]\[7\]
+ _1104_ _1105_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4575_ RF.registers\[0\]\[31\] RF.registers\[1\]\[31\] RF.registers\[2\]\[31\] RF.registers\[3\]\[31\]
+ _1324_ _1325_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__mux4_1
X_7363_ _3027_ RF.registers\[26\]\[2\] _3628_ VGND VGND VPWR VPWR _3631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9102_ clknet_leaf_21_CLK _0262_ VGND VGND VPWR VPWR RF.registers\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_7294_ _3027_ RF.registers\[31\]\[2\] _3591_ VGND VGND VPWR VPWR _3594_ sky130_fd_sc_hd__mux2_1
X_6314_ net39 VGND VGND VPWR VPWR _3029_ sky130_fd_sc_hd__clkbuf_2
X_6245_ _2675_ _2703_ _1803_ VGND VGND VPWR VPWR _2971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9033_ clknet_leaf_1_CLK _0193_ VGND VGND VPWR VPWR RF.registers\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_6176_ _2904_ _2905_ VGND VGND VPWR VPWR _2906_ sky130_fd_sc_hd__xnor2_1
X_5127_ _1723_ VGND VGND VPWR VPWR _1883_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5058_ _1812_ _1813_ _1713_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8817_ clknet_leaf_55_CLK _1001_ VGND VGND VPWR VPWR RF.registers\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8748_ clknet_leaf_9_CLK _0932_ VGND VGND VPWR VPWR RF.registers\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8679_ clknet_leaf_81_CLK _0863_ VGND VGND VPWR VPWR RF.registers\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_3 _1690_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4360_ _1112_ _1113_ _1114_ _1115_ _1047_ _1050_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__mux4_2
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4291_ net6 VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__buf_4
X_6030_ _1634_ _2767_ VGND VGND VPWR VPWR _2768_ sky130_fd_sc_hd__xor2_2
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7981_ _3103_ RF.registers\[21\]\[5\] _3952_ VGND VGND VPWR VPWR _3958_ sky130_fd_sc_hd__mux2_1
X_6932_ _3385_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6863_ RF.registers\[5\]\[8\] _3109_ _3340_ VGND VGND VPWR VPWR _3349_ sky130_fd_sc_hd__mux2_1
X_8602_ clknet_leaf_29_CLK _0786_ VGND VGND VPWR VPWR RF.registers\[22\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_5814_ _2539_ _2543_ _2562_ VGND VGND VPWR VPWR _2563_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9582_ clknet_leaf_14_CLK _0742_ VGND VGND VPWR VPWR RF.registers\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6794_ _3312_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5745_ _2327_ _1169_ _1661_ VGND VGND VPWR VPWR _2497_ sky130_fd_sc_hd__and3_1
X_8533_ RF.registers\[10\]\[9\] net45 _4244_ VGND VGND VPWR VPWR _4250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5676_ _2428_ _2429_ VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8464_ RF.registers\[11\]\[8\] net44 _4205_ VGND VGND VPWR VPWR _4214_ sky130_fd_sc_hd__mux2_1
X_7415_ _3079_ RF.registers\[26\]\[27\] _3650_ VGND VGND VPWR VPWR _3658_ sky130_fd_sc_hd__mux2_1
X_4627_ _1254_ _1382_ _1239_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_116_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8395_ _4177_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__clkbuf_1
X_7346_ _3079_ RF.registers\[31\]\[27\] _3613_ VGND VGND VPWR VPWR _3621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4558_ _1214_ _1313_ _1239_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7277_ _3584_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
X_4489_ _1243_ _1244_ _1211_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_9016_ clknet_leaf_38_CLK _0176_ VGND VGND VPWR VPWR RF.registers\[31\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_6228_ _2953_ _2954_ VGND VGND VPWR VPWR _2955_ sky130_fd_sc_hd__or2_1
X_6159_ _2015_ _2889_ VGND VGND VPWR VPWR _2890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput51 net51 VGND VGND VPWR VPWR ALU_result[11] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_56_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput73 net73 VGND VGND VPWR VPWR ALU_result[31] sky130_fd_sc_hd__buf_1
Xoutput62 net62 VGND VGND VPWR VPWR ALU_result[21] sky130_fd_sc_hd__buf_1
XFILLER_0_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5530_ _1670_ _2277_ _2281_ _2285_ VGND VGND VPWR VPWR _2286_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5461_ RF.registers\[28\]\[8\] RF.registers\[29\]\[8\] RF.registers\[30\]\[8\] RF.registers\[31\]\[8\]
+ _2051_ _2053_ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7200_ RF.registers\[7\]\[23\] _3504_ _3539_ VGND VGND VPWR VPWR _3543_ sky130_fd_sc_hd__mux2_1
X_4412_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8180_ RF.registers\[1\]\[2\] _3460_ _4061_ VGND VGND VPWR VPWR _4064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5392_ RF.registers\[28\]\[13\] RF.registers\[29\]\[13\] RF.registers\[30\]\[13\]
+ RF.registers\[31\]\[13\] _1673_ _1690_ VGND VGND VPWR VPWR _2148_ sky130_fd_sc_hd__mux4_1
X_7131_ _3505_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4343_ RF.registers\[8\]\[3\] RF.registers\[9\]\[3\] RF.registers\[10\]\[3\] RF.registers\[11\]\[3\]
+ _1042_ _1044_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__mux4_1
X_4274_ RF.registers\[20\]\[4\] RF.registers\[21\]\[4\] RF.registers\[22\]\[4\] RF.registers\[23\]\[4\]
+ _1027_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__mux4_1
X_7062_ RF.registers\[19\]\[1\] _3458_ _3456_ VGND VGND VPWR VPWR _3459_ sky130_fd_sc_hd__mux2_1
X_6013_ _2341_ _2401_ VGND VGND VPWR VPWR _2752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7964_ _3948_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_6_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6915_ RF.registers\[4\]\[0\] _3089_ _3376_ VGND VGND VPWR VPWR _3377_ sky130_fd_sc_hd__mux2_1
X_7895_ _3013_ RF.registers\[23\]\[29\] _3902_ VGND VGND VPWR VPWR _3912_ sky130_fd_sc_hd__mux2_1
X_6846_ _3339_ VGND VGND VPWR VPWR _3340_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9565_ clknet_leaf_15_CLK _0725_ VGND VGND VPWR VPWR RF.registers\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_6777_ _3005_ _3302_ VGND VGND VPWR VPWR _3303_ sky130_fd_sc_hd__nor2_2
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5728_ _2062_ _2479_ VGND VGND VPWR VPWR _2481_ sky130_fd_sc_hd__nand2_1
X_8516_ RF.registers\[10\]\[1\] net25 _3007_ VGND VGND VPWR VPWR _4241_ sky130_fd_sc_hd__mux2_1
X_9496_ clknet_leaf_42_CLK _0656_ VGND VGND VPWR VPWR RF.registers\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5659_ _2097_ _2410_ _2412_ VGND VGND VPWR VPWR _2414_ sky130_fd_sc_hd__and3_1
X_8447_ _4204_ VGND VGND VPWR VPWR _4205_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_8378_ _3155_ _3192_ VGND VGND VPWR VPWR _4168_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_130_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7329_ _3062_ RF.registers\[31\]\[19\] _3602_ VGND VGND VPWR VPWR _3612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4961_ _1716_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__clkbuf_8
X_7680_ _3798_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__clkbuf_1
X_6700_ RF.registers\[8\]\[28\] _3011_ _3253_ VGND VGND VPWR VPWR _3262_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4892_ RF.registers\[24\]\[0\] RF.registers\[25\]\[0\] RF.registers\[26\]\[0\] RF.registers\[27\]\[0\]
+ net1 net2 VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6631_ _3225_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_9350_ clknet_leaf_62_CLK _0510_ VGND VGND VPWR VPWR RF.registers\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_8301_ _4127_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__clkbuf_1
X_6562_ RF.registers\[0\]\[28\] _3011_ _3179_ VGND VGND VPWR VPWR _3188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6493_ RF.registers\[17\]\[29\] _3013_ _3135_ VGND VGND VPWR VPWR _3150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9281_ clknet_leaf_94_CLK _0441_ VGND VGND VPWR VPWR RF.registers\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_5513_ _2267_ _2268_ _1738_ VGND VGND VPWR VPWR _2269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_8232_ RF.registers\[1\]\[27\] _3444_ _4083_ VGND VGND VPWR VPWR _4091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5444_ _2198_ _2199_ _2044_ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8163_ _4054_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7114_ RF.registers\[19\]\[18\] _3493_ _3477_ VGND VGND VPWR VPWR _3494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5375_ _2127_ _2130_ _1696_ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8094_ RF.registers\[20\]\[26\] _3442_ _4011_ VGND VGND VPWR VPWR _4018_ sky130_fd_sc_hd__mux2_1
X_4326_ _1078_ _1081_ _1057_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7045_ RF.registers\[3\]\[28\] _3446_ _3435_ VGND VGND VPWR VPWR _3447_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8996_ clknet_leaf_96_CLK _0156_ VGND VGND VPWR VPWR RF.registers\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_7947_ RF.registers\[18\]\[21\] _3500_ _3938_ VGND VGND VPWR VPWR _3940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7878_ _3903_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__clkbuf_1
X_6829_ RF.registers\[6\]\[24\] _3143_ _3326_ VGND VGND VPWR VPWR _3331_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9548_ clknet_leaf_10_CLK _0708_ VGND VGND VPWR VPWR RF.registers\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9479_ clknet_leaf_81_CLK _0639_ VGND VGND VPWR VPWR RF.registers\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_78_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5160_ _1773_ _1915_ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_87_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5091_ RF.registers\[24\]\[17\] RF.registers\[25\]\[17\] RF.registers\[26\]\[17\]
+ RF.registers\[27\]\[17\] _1689_ _1693_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__mux4_1
X_8850_ clknet_leaf_54_CLK _0010_ VGND VGND VPWR VPWR RF.registers\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7801_ _3862_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__clkbuf_1
X_5993_ _2327_ _2675_ _2732_ VGND VGND VPWR VPWR _2733_ sky130_fd_sc_hd__a21o_1
X_8781_ clknet_leaf_57_CLK _0965_ VGND VGND VPWR VPWR RF.registers\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4944_ _1699_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__buf_4
X_7732_ _3056_ RF.registers\[30\]\[16\] _3819_ VGND VGND VPWR VPWR _3826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_9402_ clknet_leaf_24_CLK _0562_ VGND VGND VPWR VPWR RF.registers\[24\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_4875_ RF.registers\[0\]\[18\] RF.registers\[1\]\[18\] RF.registers\[2\]\[18\] RF.registers\[3\]\[18\]
+ _1173_ _1175_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__mux4_1
X_7663_ _3789_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6614_ _3216_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7594_ _3054_ RF.registers\[28\]\[15\] _3747_ VGND VGND VPWR VPWR _3753_ sky130_fd_sc_hd__mux2_1
X_9333_ clknet_leaf_29_CLK _0493_ VGND VGND VPWR VPWR RF.registers\[21\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_6545_ _3156_ VGND VGND VPWR VPWR _3179_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9264_ clknet_leaf_7_CLK _0424_ VGND VGND VPWR VPWR RF.registers\[23\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6476_ RF.registers\[17\]\[22\] _3139_ _3135_ VGND VGND VPWR VPWR _3140_ sky130_fd_sc_hd__mux2_1
X_8215_ RF.registers\[1\]\[19\] _3495_ _4072_ VGND VGND VPWR VPWR _4082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9195_ clknet_leaf_98_CLK _0355_ VGND VGND VPWR VPWR RF.registers\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_5427_ RF.registers\[20\]\[11\] RF.registers\[21\]\[11\] RF.registers\[22\]\[11\]
+ RF.registers\[23\]\[11\] _1675_ _1692_ VGND VGND VPWR VPWR _2183_ sky130_fd_sc_hd__mux4_1
XFILLER_0_100_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8146_ _4045_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__clkbuf_1
X_5358_ _2052_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__buf_4
X_8077_ RF.registers\[20\]\[18\] _3493_ _4000_ VGND VGND VPWR VPWR _4009_ sky130_fd_sc_hd__mux2_1
X_4309_ A2[0] VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__buf_4
X_7028_ RF.registers\[3\]\[21\] _3137_ _3435_ VGND VGND VPWR VPWR _3437_ sky130_fd_sc_hd__mux2_1
X_5289_ _2042_ _2043_ _2044_ VGND VGND VPWR VPWR _2045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_8979_ clknet_leaf_25_CLK _0139_ VGND VGND VPWR VPWR RF.registers\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4660_ _1399_ _1415_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4591_ _1341_ _1343_ _1346_ _1187_ _1215_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_12_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6330_ _3039_ RF.registers\[22\]\[8\] _3023_ VGND VGND VPWR VPWR _3040_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6261_ _2934_ _2940_ _2951_ _2932_ VGND VGND VPWR VPWR _2987_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5212_ _1966_ _1967_ _1745_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6192_ _2918_ _2920_ VGND VGND VPWR VPWR _2921_ sky130_fd_sc_hd__xor2_1
X_8000_ _3122_ RF.registers\[21\]\[14\] _3963_ VGND VGND VPWR VPWR _3968_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5143_ RF.registers\[4\]\[31\] RF.registers\[5\]\[31\] RF.registers\[6\]\[31\] RF.registers\[7\]\[31\]
+ _1896_ _1898_ VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__mux4_1
X_5074_ RF.registers\[12\]\[19\] RF.registers\[13\]\[19\] RF.registers\[14\]\[19\]
+ RF.registers\[15\]\[19\] _1689_ _1693_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8902_ clknet_leaf_62_CLK _0062_ VGND VGND VPWR VPWR RF.registers\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_8833_ clknet_leaf_72_CLK _1017_ VGND VGND VPWR VPWR RF.registers\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_121_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8764_ clknet_leaf_17_CLK _0948_ VGND VGND VPWR VPWR RF.registers\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_5976_ _2344_ _2342_ VGND VGND VPWR VPWR _2717_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8695_ clknet_leaf_47_CLK _0879_ VGND VGND VPWR VPWR RF.registers\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4927_ RF.registers\[16\]\[23\] RF.registers\[17\]\[23\] RF.registers\[18\]\[23\]
+ RF.registers\[19\]\[23\] _1676_ _1681_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__mux4_1
X_7715_ _3039_ RF.registers\[30\]\[8\] _3808_ VGND VGND VPWR VPWR _3817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4858_ RF.registers\[8\]\[19\] RF.registers\[9\]\[19\] RF.registers\[10\]\[19\] RF.registers\[11\]\[19\]
+ _1173_ _1175_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7646_ _3780_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_9316_ clknet_leaf_94_CLK _0476_ VGND VGND VPWR VPWR RF.registers\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_4789_ _1543_ _1544_ _1034_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__mux2_1
X_7577_ _3037_ RF.registers\[28\]\[7\] _3736_ VGND VGND VPWR VPWR _3744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_80_CLK sky130_fd_sc_hd__clkbuf_8
X_6528_ _3170_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_132_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6459_ net22 VGND VGND VPWR VPWR _3128_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9247_ clknet_leaf_64_CLK _0407_ VGND VGND VPWR VPWR RF.registers\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_9178_ clknet_leaf_35_CLK _0338_ VGND VGND VPWR VPWR RF.registers\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8129_ RF.registers\[24\]\[10\] _3476_ _4036_ VGND VGND VPWR VPWR _4037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_CLK clknet_3_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_71_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5830_ _2577_ _2498_ _1803_ VGND VGND VPWR VPWR _2578_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5761_ _2511_ _2512_ VGND VGND VPWR VPWR _2513_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8480_ _4222_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__clkbuf_1
X_7500_ _3703_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
X_4712_ RF.registers\[28\]\[13\] RF.registers\[29\]\[13\] RF.registers\[30\]\[13\]
+ RF.registers\[31\]\[13\] _1027_ _1029_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5692_ _1666_ _2445_ VGND VGND VPWR VPWR _2446_ sky130_fd_sc_hd__nor2_1
X_7431_ _3027_ RF.registers\[25\]\[2\] _3664_ VGND VGND VPWR VPWR _3667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4643_ _1025_ _1390_ _1398_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__o21ai_4
X_4574_ RF.registers\[4\]\[31\] RF.registers\[5\]\[31\] RF.registers\[6\]\[31\] RF.registers\[7\]\[31\]
+ _1324_ _1325_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__mux4_1
X_7362_ _3630_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_62_CLK clknet_3_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_62_CLK sky130_fd_sc_hd__clkbuf_8
X_9101_ clknet_leaf_4_CLK _0261_ VGND VGND VPWR VPWR RF.registers\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_6313_ _3028_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__clkbuf_1
X_7293_ _3593_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6244_ _2672_ _2674_ _1803_ VGND VGND VPWR VPWR _2970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_9032_ clknet_leaf_1_CLK _0192_ VGND VGND VPWR VPWR RF.registers\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_6175_ _2887_ _2890_ _2892_ VGND VGND VPWR VPWR _2905_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5126_ _1881_ VGND VGND VPWR VPWR _1882_ sky130_fd_sc_hd__buf_4
X_5057_ RF.registers\[12\]\[18\] RF.registers\[13\]\[18\] RF.registers\[14\]\[18\]
+ RF.registers\[15\]\[18\] _1689_ _1693_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8816_ clknet_leaf_58_CLK _1000_ VGND VGND VPWR VPWR RF.registers\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5959_ _2335_ _2701_ VGND VGND VPWR VPWR _2702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8747_ clknet_leaf_89_CLK _0931_ VGND VGND VPWR VPWR RF.registers\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8678_ clknet_leaf_63_CLK _0862_ VGND VGND VPWR VPWR RF.registers\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7629_ _3005_ _3153_ VGND VGND VPWR VPWR _3771_ sky130_fd_sc_hd__nor2_4
XFILLER_0_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_53_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_CLK clknet_3_6__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_44_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _1700_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4290_ _1040_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_60_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7980_ _3957_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6931_ RF.registers\[4\]\[8\] _3109_ _3376_ VGND VGND VPWR VPWR _3385_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6862_ _3348_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_8601_ clknet_leaf_27_CLK _0785_ VGND VGND VPWR VPWR RF.registers\[22\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_5813_ _2271_ _2538_ VGND VGND VPWR VPWR _2562_ sky130_fd_sc_hd__or2_1
X_9581_ clknet_leaf_11_CLK _0741_ VGND VGND VPWR VPWR RF.registers\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6793_ RF.registers\[6\]\[7\] _3107_ _3304_ VGND VGND VPWR VPWR _3312_ sky130_fd_sc_hd__mux2_1
X_8532_ _4249_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__clkbuf_1
X_5744_ _2495_ VGND VGND VPWR VPWR _2496_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5675_ _1800_ _2247_ VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__nor2_1
X_8463_ _4213_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__clkbuf_1
X_4626_ _1380_ _1381_ _1190_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_CLK clknet_3_7__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_35_CLK sky130_fd_sc_hd__clkbuf_8
X_7414_ _3657_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_8394_ RF.registers\[12\]\[7\] _3470_ _4169_ VGND VGND VPWR VPWR _4177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7345_ _3620_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4557_ _1311_ _1312_ _1199_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_7276_ _3077_ RF.registers\[29\]\[26\] _3577_ VGND VGND VPWR VPWR _3584_ sky130_fd_sc_hd__mux2_1
X_4488_ RF.registers\[24\]\[20\] RF.registers\[25\]\[20\] RF.registers\[26\]\[20\]
+ RF.registers\[27\]\[20\] _1207_ _1208_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__mux4_1
X_9015_ clknet_leaf_31_CLK _0175_ VGND VGND VPWR VPWR RF.registers\[31\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6227_ _2934_ _2940_ _2932_ VGND VGND VPWR VPWR _2954_ sky130_fd_sc_hd__a21oi_1
X_6158_ _1370_ _2888_ VGND VGND VPWR VPWR _2889_ sky130_fd_sc_hd__xor2_1
X_5109_ _1861_ _1862_ _1863_ _1864_ _1713_ _1717_ VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__mux4_1
X_6089_ _2756_ _2751_ _2426_ VGND VGND VPWR VPWR _2824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_26_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput52 net52 VGND VGND VPWR VPWR ALU_result[12] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_56_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput63 net63 VGND VGND VPWR VPWR ALU_result[22] sky130_fd_sc_hd__buf_1
Xoutput74 net74 VGND VGND VPWR VPWR ALU_result[3] sky130_fd_sc_hd__buf_1
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_CLK clknet_3_5__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_17_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5460_ _2214_ _2215_ _1685_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4411_ _1166_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5391_ _2145_ _2146_ _1684_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__mux2_1
X_7130_ RF.registers\[19\]\[23\] _3504_ _3498_ VGND VGND VPWR VPWR _3505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4342_ _1038_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4273_ _1028_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__buf_4
X_7061_ net25 VGND VGND VPWR VPWR _3458_ sky130_fd_sc_hd__buf_2
X_6012_ _2649_ _2697_ _2327_ VGND VGND VPWR VPWR _2751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

