VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO project1
  CLASS BLOCK ;
  FOREIGN project1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 60.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 49.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 49.200 ;
    END
  END VPWR
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END in[0]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END in[1]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END in[2]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END in[3]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END in[4]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END in[5]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END in[6]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END in[7]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END out[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 34.230 49.045 ;
      LAYER li1 ;
        RECT 5.520 10.795 34.040 49.045 ;
      LAYER met1 ;
        RECT 4.210 10.640 34.040 49.200 ;
      LAYER met2 ;
        RECT 4.230 3.555 32.560 54.925 ;
      LAYER met3 ;
        RECT 4.400 54.040 14.610 54.905 ;
        RECT 3.990 52.040 14.610 54.040 ;
        RECT 4.400 50.640 14.610 52.040 ;
        RECT 3.990 48.640 14.610 50.640 ;
        RECT 4.400 47.240 14.610 48.640 ;
        RECT 3.990 45.240 14.610 47.240 ;
        RECT 4.400 43.840 14.610 45.240 ;
        RECT 3.990 41.840 14.610 43.840 ;
        RECT 4.400 40.440 14.610 41.840 ;
        RECT 3.990 38.440 14.610 40.440 ;
        RECT 4.400 37.040 14.610 38.440 ;
        RECT 3.990 35.040 14.610 37.040 ;
        RECT 4.400 33.640 14.610 35.040 ;
        RECT 3.990 31.640 14.610 33.640 ;
        RECT 4.400 30.240 14.610 31.640 ;
        RECT 3.990 28.240 14.610 30.240 ;
        RECT 4.400 26.840 14.610 28.240 ;
        RECT 3.990 24.840 14.610 26.840 ;
        RECT 4.400 23.440 14.610 24.840 ;
        RECT 3.990 21.440 14.610 23.440 ;
        RECT 4.400 20.040 14.610 21.440 ;
        RECT 3.990 18.040 14.610 20.040 ;
        RECT 4.400 16.640 14.610 18.040 ;
        RECT 3.990 14.640 14.610 16.640 ;
        RECT 4.400 13.240 14.610 14.640 ;
        RECT 3.990 11.240 14.610 13.240 ;
        RECT 4.400 9.840 14.610 11.240 ;
        RECT 3.990 7.840 14.610 9.840 ;
        RECT 4.400 6.440 14.610 7.840 ;
        RECT 3.990 4.440 14.610 6.440 ;
        RECT 4.400 3.575 14.610 4.440 ;
  END
END project1
END LIBRARY

