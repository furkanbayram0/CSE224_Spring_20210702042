magic
tech sky130A
magscale 1 2
timestamp 1746400034
<< checkpaint >>
rect -3932 -3932 23932 23932
<< viali >>
rect 10517 17833 10551 17867
rect 12541 17833 12575 17867
rect 11897 17765 11931 17799
rect 9229 17629 9263 17663
rect 9965 17629 9999 17663
rect 10701 17629 10735 17663
rect 11253 17629 11287 17663
rect 11713 17629 11747 17663
rect 12725 17629 12759 17663
rect 9413 17561 9447 17595
rect 10057 17493 10091 17527
rect 11161 17493 11195 17527
rect 10701 14433 10735 14467
rect 10609 14365 10643 14399
rect 10977 14229 11011 14263
rect 10701 14025 10735 14059
rect 11529 14025 11563 14059
rect 13093 13957 13127 13991
rect 8585 13889 8619 13923
rect 9781 13889 9815 13923
rect 9965 13889 9999 13923
rect 10241 13889 10275 13923
rect 10425 13889 10459 13923
rect 11345 13889 11379 13923
rect 11437 13889 11471 13923
rect 12817 13889 12851 13923
rect 13277 13889 13311 13923
rect 8677 13821 8711 13855
rect 10057 13821 10091 13855
rect 10885 13821 10919 13855
rect 10977 13821 11011 13855
rect 11069 13821 11103 13855
rect 11161 13821 11195 13855
rect 11805 13821 11839 13855
rect 12449 13821 12483 13855
rect 12909 13821 12943 13855
rect 13461 13821 13495 13855
rect 8953 13753 8987 13787
rect 9873 13685 9907 13719
rect 8493 13481 8527 13515
rect 8861 13481 8895 13515
rect 10977 13481 11011 13515
rect 13001 13481 13035 13515
rect 13369 13481 13403 13515
rect 11069 13413 11103 13447
rect 13553 13345 13587 13379
rect 13737 13345 13771 13379
rect 8953 13277 8987 13311
rect 9229 13277 9263 13311
rect 9505 13277 9539 13311
rect 10425 13277 10459 13311
rect 10609 13277 10643 13311
rect 10701 13277 10735 13311
rect 10793 13277 10827 13311
rect 11069 13277 11103 13311
rect 11253 13277 11287 13311
rect 13277 13277 13311 13311
rect 13369 13277 13403 13311
rect 13461 13277 13495 13311
rect 9045 13209 9079 13243
rect 9413 13209 9447 13243
rect 10517 13209 10551 13243
rect 10977 13209 11011 13243
rect 13737 13141 13771 13175
rect 8953 12937 8987 12971
rect 9045 12937 9079 12971
rect 13461 12937 13495 12971
rect 13645 12937 13679 12971
rect 8769 12869 8803 12903
rect 2605 12801 2639 12835
rect 6745 12801 6779 12835
rect 8585 12801 8619 12835
rect 9229 12801 9263 12835
rect 9413 12801 9447 12835
rect 13185 12801 13219 12835
rect 13277 12801 13311 12835
rect 13553 12801 13587 12835
rect 13737 12801 13771 12835
rect 16865 12801 16899 12835
rect 6837 12733 6871 12767
rect 16313 12733 16347 12767
rect 16589 12733 16623 12767
rect 7113 12665 7147 12699
rect 2421 12597 2455 12631
rect 6929 12393 6963 12427
rect 7297 12393 7331 12427
rect 7389 12393 7423 12427
rect 8769 12393 8803 12427
rect 10149 12393 10183 12427
rect 12081 12393 12115 12427
rect 12541 12393 12575 12427
rect 8953 12325 8987 12359
rect 6653 12257 6687 12291
rect 7481 12257 7515 12291
rect 8585 12257 8619 12291
rect 9413 12257 9447 12291
rect 10517 12257 10551 12291
rect 6561 12189 6595 12223
rect 7205 12189 7239 12223
rect 8493 12189 8527 12223
rect 9137 12189 9171 12223
rect 9321 12189 9355 12223
rect 10425 12189 10459 12223
rect 11989 12189 12023 12223
rect 12265 12189 12299 12223
rect 12357 12189 12391 12223
rect 9781 11849 9815 11883
rect 11805 11849 11839 11883
rect 12449 11849 12483 11883
rect 13185 11849 13219 11883
rect 13829 11849 13863 11883
rect 11161 11781 11195 11815
rect 2605 11713 2639 11747
rect 9965 11713 9999 11747
rect 10149 11713 10183 11747
rect 10241 11713 10275 11747
rect 10609 11713 10643 11747
rect 10885 11713 10919 11747
rect 10977 11713 11011 11747
rect 11253 11713 11287 11747
rect 11345 11713 11379 11747
rect 11529 11713 11563 11747
rect 11621 11713 11655 11747
rect 12633 11713 12667 11747
rect 12725 11713 12759 11747
rect 12817 11713 12851 11747
rect 13001 11713 13035 11747
rect 13093 11713 13127 11747
rect 13369 11713 13403 11747
rect 13461 11713 13495 11747
rect 13737 11713 13771 11747
rect 14013 11713 14047 11747
rect 14289 11713 14323 11747
rect 17325 11713 17359 11747
rect 10701 11645 10735 11679
rect 2421 11577 2455 11611
rect 13645 11577 13679 11611
rect 14105 11577 14139 11611
rect 14197 11577 14231 11611
rect 17141 11577 17175 11611
rect 7665 11305 7699 11339
rect 8677 11305 8711 11339
rect 9137 11305 9171 11339
rect 10977 11305 11011 11339
rect 12541 11305 12575 11339
rect 13553 11305 13587 11339
rect 14289 11305 14323 11339
rect 17417 11305 17451 11339
rect 2513 11237 2547 11271
rect 14841 11237 14875 11271
rect 2329 11101 2363 11135
rect 7021 11101 7055 11135
rect 7205 11101 7239 11135
rect 7297 11101 7331 11135
rect 7389 11101 7423 11135
rect 8861 11101 8895 11135
rect 8953 11101 8987 11135
rect 9229 11101 9263 11135
rect 10701 11101 10735 11135
rect 12817 11101 12851 11135
rect 13737 11101 13771 11135
rect 13921 11101 13955 11135
rect 14013 11101 14047 11135
rect 14565 11101 14599 11135
rect 14657 11101 14691 11135
rect 14841 11101 14875 11135
rect 10977 11033 11011 11067
rect 12541 11033 12575 11067
rect 14105 11033 14139 11067
rect 14305 11033 14339 11067
rect 17509 11033 17543 11067
rect 10793 10965 10827 10999
rect 12725 10965 12759 10999
rect 14473 10965 14507 10999
rect 6377 10761 6411 10795
rect 7113 10761 7147 10795
rect 9597 10761 9631 10795
rect 10977 10761 11011 10795
rect 11897 10761 11931 10795
rect 7665 10693 7699 10727
rect 9045 10693 9079 10727
rect 9137 10693 9171 10727
rect 9965 10693 9999 10727
rect 10701 10693 10735 10727
rect 11621 10693 11655 10727
rect 2605 10625 2639 10659
rect 6009 10625 6043 10659
rect 6469 10625 6503 10659
rect 6653 10625 6687 10659
rect 6929 10625 6963 10659
rect 7297 10625 7331 10659
rect 7481 10625 7515 10659
rect 7573 10625 7607 10659
rect 7783 10625 7817 10659
rect 7941 10625 7975 10659
rect 8125 10625 8159 10659
rect 8341 10625 8375 10659
rect 8493 10625 8527 10659
rect 8953 10625 8987 10659
rect 9321 10625 9355 10659
rect 9413 10625 9447 10659
rect 9505 10625 9539 10659
rect 9781 10625 9815 10659
rect 9873 10625 9907 10659
rect 10057 10625 10091 10659
rect 10333 10625 10367 10659
rect 10481 10625 10515 10659
rect 10609 10625 10643 10659
rect 10839 10625 10873 10659
rect 11253 10625 11287 10659
rect 11346 10625 11380 10659
rect 11529 10625 11563 10659
rect 11718 10625 11752 10659
rect 14565 10625 14599 10659
rect 14841 10625 14875 10659
rect 15117 10625 15151 10659
rect 17417 10625 17451 10659
rect 2329 10557 2363 10591
rect 5917 10557 5951 10591
rect 8217 10557 8251 10591
rect 14657 10557 14691 10591
rect 15393 10557 15427 10591
rect 9781 10489 9815 10523
rect 15209 10489 15243 10523
rect 17233 10489 17267 10523
rect 8677 10421 8711 10455
rect 8769 10421 8803 10455
rect 15025 10421 15059 10455
rect 15117 10421 15151 10455
rect 6929 10217 6963 10251
rect 7021 10217 7055 10251
rect 9229 10217 9263 10251
rect 10241 10217 10275 10251
rect 11069 10217 11103 10251
rect 15393 10149 15427 10183
rect 7113 10081 7147 10115
rect 10425 10081 10459 10115
rect 11989 10081 12023 10115
rect 13369 10081 13403 10115
rect 15301 10081 15335 10115
rect 6837 10013 6871 10047
rect 8585 10013 8619 10047
rect 8733 10013 8767 10047
rect 8861 10013 8895 10047
rect 8953 10013 8987 10047
rect 9091 10013 9125 10047
rect 10517 10013 10551 10047
rect 10609 10013 10643 10047
rect 10701 10013 10735 10047
rect 10885 10013 10919 10047
rect 11069 10013 11103 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 11437 10013 11471 10047
rect 11529 10013 11563 10047
rect 11713 10013 11747 10047
rect 11805 10013 11839 10047
rect 12357 10013 12391 10047
rect 12449 10013 12483 10047
rect 12541 10013 12575 10047
rect 12817 10013 12851 10047
rect 13093 10013 13127 10047
rect 13185 10013 13219 10047
rect 13461 10013 13495 10047
rect 13553 10013 13587 10047
rect 13737 10013 13771 10047
rect 13829 10013 13863 10047
rect 14657 10013 14691 10047
rect 14841 10013 14875 10047
rect 15025 10013 15059 10047
rect 15209 10013 15243 10047
rect 15485 10013 15519 10047
rect 17325 10013 17359 10047
rect 11253 9945 11287 9979
rect 12173 9945 12207 9979
rect 12679 9945 12713 9979
rect 12909 9877 12943 9911
rect 13651 9877 13685 9911
rect 14749 9877 14783 9911
rect 15669 9877 15703 9911
rect 17509 9877 17543 9911
rect 10609 9673 10643 9707
rect 9045 9605 9079 9639
rect 13185 9605 13219 9639
rect 8677 9537 8711 9571
rect 8861 9537 8895 9571
rect 9137 9537 9171 9571
rect 10517 9537 10551 9571
rect 10701 9537 10735 9571
rect 12633 9537 12667 9571
rect 12725 9537 12759 9571
rect 12909 9537 12943 9571
rect 13001 9537 13035 9571
rect 14657 9537 14691 9571
rect 15209 9537 15243 9571
rect 14197 9469 14231 9503
rect 14381 9469 14415 9503
rect 14473 9469 14507 9503
rect 14565 9469 14599 9503
rect 15301 9469 15335 9503
rect 9321 9401 9355 9435
rect 14841 9333 14875 9367
rect 7389 9129 7423 9163
rect 8677 9129 8711 9163
rect 8861 9129 8895 9163
rect 9137 9129 9171 9163
rect 15485 9129 15519 9163
rect 7113 9061 7147 9095
rect 7573 9061 7607 9095
rect 8585 8993 8619 9027
rect 6929 8925 6963 8959
rect 7757 8925 7791 8959
rect 8309 8925 8343 8959
rect 9413 8925 9447 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 10517 8925 10551 8959
rect 15025 8925 15059 8959
rect 15301 8925 15335 8959
rect 2421 8857 2455 8891
rect 2605 8857 2639 8891
rect 7205 8857 7239 8891
rect 7941 8857 7975 8891
rect 8125 8857 8159 8891
rect 8962 8857 8996 8891
rect 9137 8857 9171 8891
rect 10425 8857 10459 8891
rect 17325 8857 17359 8891
rect 17509 8857 17543 8891
rect 7389 8789 7423 8823
rect 10701 8789 10735 8823
rect 15117 8789 15151 8823
rect 8217 8585 8251 8619
rect 8861 8585 8895 8619
rect 7389 8517 7423 8551
rect 7573 8517 7607 8551
rect 8401 8517 8435 8551
rect 9413 8517 9447 8551
rect 12725 8517 12759 8551
rect 12817 8517 12851 8551
rect 6929 8449 6963 8483
rect 7021 8449 7055 8483
rect 8769 8449 8803 8483
rect 9229 8449 9263 8483
rect 9321 8449 9355 8483
rect 9597 8449 9631 8483
rect 10057 8449 10091 8483
rect 10241 8449 10275 8483
rect 10425 8449 10459 8483
rect 10517 8449 10551 8483
rect 10977 8449 11011 8483
rect 11253 8449 11287 8483
rect 11529 8449 11563 8483
rect 11713 8449 11747 8483
rect 12449 8449 12483 8483
rect 12542 8449 12576 8483
rect 12955 8449 12989 8483
rect 13185 8449 13219 8483
rect 13645 8449 13679 8483
rect 14841 8449 14875 8483
rect 17141 8449 17175 8483
rect 10609 8381 10643 8415
rect 10701 8381 10735 8415
rect 10885 8381 10919 8415
rect 11069 8381 11103 8415
rect 11621 8381 11655 8415
rect 13369 8381 13403 8415
rect 13461 8381 13495 8415
rect 14473 8381 14507 8415
rect 14749 8381 14783 8415
rect 9045 8313 9079 8347
rect 10241 8313 10275 8347
rect 11437 8313 11471 8347
rect 13093 8313 13127 8347
rect 13553 8313 13587 8347
rect 13829 8313 13863 8347
rect 17325 8313 17359 8347
rect 7573 8245 7607 8279
rect 7757 8245 7791 8279
rect 8033 8245 8067 8279
rect 8217 8245 8251 8279
rect 11253 8245 11287 8279
rect 7573 8041 7607 8075
rect 11253 8041 11287 8075
rect 13185 8041 13219 8075
rect 13829 8041 13863 8075
rect 15025 8041 15059 8075
rect 11345 7973 11379 8007
rect 12265 7973 12299 8007
rect 10149 7905 10183 7939
rect 10793 7905 10827 7939
rect 12725 7905 12759 7939
rect 12817 7905 12851 7939
rect 12909 7905 12943 7939
rect 13001 7905 13035 7939
rect 13369 7905 13403 7939
rect 10241 7837 10275 7871
rect 10425 7837 10459 7871
rect 10701 7837 10735 7871
rect 10977 7837 11011 7871
rect 11069 7837 11103 7871
rect 11621 7837 11655 7871
rect 12541 7837 12575 7871
rect 13277 7837 13311 7871
rect 13553 7837 13587 7871
rect 13645 7837 13679 7871
rect 13921 7837 13955 7871
rect 15025 7837 15059 7871
rect 15209 7837 15243 7871
rect 17325 7837 17359 7871
rect 17601 7837 17635 7871
rect 7665 7769 7699 7803
rect 11345 7769 11379 7803
rect 12265 7769 12299 7803
rect 10609 7701 10643 7735
rect 11529 7701 11563 7735
rect 12449 7701 12483 7735
rect 14013 7701 14047 7735
rect 7757 7497 7791 7531
rect 13369 7497 13403 7531
rect 14749 7497 14783 7531
rect 7021 7429 7055 7463
rect 14381 7429 14415 7463
rect 14581 7429 14615 7463
rect 15117 7429 15151 7463
rect 7113 7361 7147 7395
rect 7297 7361 7331 7395
rect 8125 7361 8159 7395
rect 8861 7361 8895 7395
rect 8953 7361 8987 7395
rect 9137 7361 9171 7395
rect 13001 7361 13035 7395
rect 14841 7361 14875 7395
rect 14933 7361 14967 7395
rect 7389 7293 7423 7327
rect 8033 7293 8067 7327
rect 13093 7293 13127 7327
rect 8585 7225 8619 7259
rect 15117 7225 15151 7259
rect 7481 7157 7515 7191
rect 7665 7157 7699 7191
rect 7941 7157 7975 7191
rect 8401 7157 8435 7191
rect 8953 7157 8987 7191
rect 13001 7157 13035 7191
rect 14565 7157 14599 7191
rect 7573 6953 7607 6987
rect 8953 6953 8987 6987
rect 11621 6953 11655 6987
rect 14105 6953 14139 6987
rect 14473 6953 14507 6987
rect 8217 6885 8251 6919
rect 9045 6817 9079 6851
rect 7665 6749 7699 6783
rect 7849 6749 7883 6783
rect 8125 6749 8159 6783
rect 8493 6749 8527 6783
rect 8585 6749 8619 6783
rect 8953 6749 8987 6783
rect 9229 6749 9263 6783
rect 9689 6749 9723 6783
rect 10057 6749 10091 6783
rect 10241 6749 10275 6783
rect 12265 6749 12299 6783
rect 12357 6749 12391 6783
rect 13093 6749 13127 6783
rect 13461 6749 13495 6783
rect 13645 6749 13679 6783
rect 13921 6749 13955 6783
rect 14473 6749 14507 6783
rect 8861 6681 8895 6715
rect 9873 6681 9907 6715
rect 11805 6681 11839 6715
rect 12081 6681 12115 6715
rect 13277 6681 13311 6715
rect 14197 6681 14231 6715
rect 14381 6681 14415 6715
rect 7941 6613 7975 6647
rect 8401 6613 8435 6647
rect 9413 6613 9447 6647
rect 9505 6613 9539 6647
rect 11437 6613 11471 6647
rect 11605 6613 11639 6647
rect 12179 6613 12213 6647
rect 13737 6613 13771 6647
rect 8769 6409 8803 6443
rect 10425 6409 10459 6443
rect 11805 6341 11839 6375
rect 11897 6341 11931 6375
rect 12265 6341 12299 6375
rect 8033 6273 8067 6307
rect 8217 6273 8251 6307
rect 8309 6273 8343 6307
rect 8585 6273 8619 6307
rect 10057 6273 10091 6307
rect 10517 6273 10551 6307
rect 10701 6273 10735 6307
rect 10793 6273 10827 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 11253 6273 11287 6307
rect 11529 6273 11563 6307
rect 11989 6273 12023 6307
rect 8401 6205 8435 6239
rect 10149 6205 10183 6239
rect 10609 6205 10643 6239
rect 11345 6205 11379 6239
rect 12265 6205 12299 6239
rect 12081 6069 12115 6103
rect 11529 5865 11563 5899
rect 11437 5797 11471 5831
rect 11345 5661 11379 5695
rect 11621 5593 11655 5627
rect 10701 3009 10735 3043
rect 10517 2805 10551 2839
rect 8769 2601 8803 2635
rect 11253 2601 11287 2635
rect 11989 2533 12023 2567
rect 8125 2465 8159 2499
rect 9873 2465 9907 2499
rect 10149 2465 10183 2499
rect 12725 2465 12759 2499
rect 7849 2397 7883 2431
rect 8953 2397 8987 2431
rect 9413 2397 9447 2431
rect 11069 2397 11103 2431
rect 12449 2397 12483 2431
rect 11805 2329 11839 2363
rect 9597 2261 9631 2295
<< metal1 >>
rect 2024 17978 17940 18000
rect 2024 17926 3859 17978
rect 3911 17926 3923 17978
rect 3975 17926 3987 17978
rect 4039 17926 4051 17978
rect 4103 17926 4115 17978
rect 4167 17926 7838 17978
rect 7890 17926 7902 17978
rect 7954 17926 7966 17978
rect 8018 17926 8030 17978
rect 8082 17926 8094 17978
rect 8146 17926 11817 17978
rect 11869 17926 11881 17978
rect 11933 17926 11945 17978
rect 11997 17926 12009 17978
rect 12061 17926 12073 17978
rect 12125 17926 15796 17978
rect 15848 17926 15860 17978
rect 15912 17926 15924 17978
rect 15976 17926 15988 17978
rect 16040 17926 16052 17978
rect 16104 17926 17940 17978
rect 2024 17904 17940 17926
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 10505 17867 10563 17873
rect 10505 17864 10517 17867
rect 10376 17836 10517 17864
rect 10376 17824 10382 17836
rect 10505 17833 10517 17836
rect 10551 17833 10563 17867
rect 10505 17827 10563 17833
rect 12250 17824 12256 17876
rect 12308 17864 12314 17876
rect 12529 17867 12587 17873
rect 12529 17864 12541 17867
rect 12308 17836 12541 17864
rect 12308 17824 12314 17836
rect 12529 17833 12541 17836
rect 12575 17833 12587 17867
rect 12529 17827 12587 17833
rect 10594 17756 10600 17808
rect 10652 17796 10658 17808
rect 11885 17799 11943 17805
rect 11885 17796 11897 17799
rect 10652 17768 11897 17796
rect 10652 17756 10658 17768
rect 11885 17765 11897 17768
rect 11931 17765 11943 17799
rect 11885 17759 11943 17765
rect 9030 17620 9036 17672
rect 9088 17660 9094 17672
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 9088 17632 9229 17660
rect 9088 17620 9094 17632
rect 9217 17629 9229 17632
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 9953 17663 10011 17669
rect 9953 17660 9965 17663
rect 9732 17632 9965 17660
rect 9732 17620 9738 17632
rect 9953 17629 9965 17632
rect 9999 17629 10011 17663
rect 9953 17623 10011 17629
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17629 10747 17663
rect 10689 17623 10747 17629
rect 9398 17552 9404 17604
rect 9456 17552 9462 17604
rect 10704 17592 10732 17623
rect 10962 17620 10968 17672
rect 11020 17660 11026 17672
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 11020 17632 11253 17660
rect 11020 17620 11026 17632
rect 11241 17629 11253 17632
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11664 17632 11713 17660
rect 11664 17620 11670 17632
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17660 12771 17663
rect 12802 17660 12808 17672
rect 12759 17632 12808 17660
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 11422 17592 11428 17604
rect 10704 17564 11428 17592
rect 11422 17552 11428 17564
rect 11480 17552 11486 17604
rect 10042 17484 10048 17536
rect 10100 17484 10106 17536
rect 11149 17527 11207 17533
rect 11149 17493 11161 17527
rect 11195 17524 11207 17527
rect 11330 17524 11336 17536
rect 11195 17496 11336 17524
rect 11195 17493 11207 17496
rect 11149 17487 11207 17493
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 2024 17434 17940 17456
rect 2024 17382 4519 17434
rect 4571 17382 4583 17434
rect 4635 17382 4647 17434
rect 4699 17382 4711 17434
rect 4763 17382 4775 17434
rect 4827 17382 8498 17434
rect 8550 17382 8562 17434
rect 8614 17382 8626 17434
rect 8678 17382 8690 17434
rect 8742 17382 8754 17434
rect 8806 17382 12477 17434
rect 12529 17382 12541 17434
rect 12593 17382 12605 17434
rect 12657 17382 12669 17434
rect 12721 17382 12733 17434
rect 12785 17382 16456 17434
rect 16508 17382 16520 17434
rect 16572 17382 16584 17434
rect 16636 17382 16648 17434
rect 16700 17382 16712 17434
rect 16764 17382 17940 17434
rect 2024 17360 17940 17382
rect 2024 16890 17940 16912
rect 2024 16838 3859 16890
rect 3911 16838 3923 16890
rect 3975 16838 3987 16890
rect 4039 16838 4051 16890
rect 4103 16838 4115 16890
rect 4167 16838 7838 16890
rect 7890 16838 7902 16890
rect 7954 16838 7966 16890
rect 8018 16838 8030 16890
rect 8082 16838 8094 16890
rect 8146 16838 11817 16890
rect 11869 16838 11881 16890
rect 11933 16838 11945 16890
rect 11997 16838 12009 16890
rect 12061 16838 12073 16890
rect 12125 16838 15796 16890
rect 15848 16838 15860 16890
rect 15912 16838 15924 16890
rect 15976 16838 15988 16890
rect 16040 16838 16052 16890
rect 16104 16838 17940 16890
rect 2024 16816 17940 16838
rect 2024 16346 17940 16368
rect 2024 16294 4519 16346
rect 4571 16294 4583 16346
rect 4635 16294 4647 16346
rect 4699 16294 4711 16346
rect 4763 16294 4775 16346
rect 4827 16294 8498 16346
rect 8550 16294 8562 16346
rect 8614 16294 8626 16346
rect 8678 16294 8690 16346
rect 8742 16294 8754 16346
rect 8806 16294 12477 16346
rect 12529 16294 12541 16346
rect 12593 16294 12605 16346
rect 12657 16294 12669 16346
rect 12721 16294 12733 16346
rect 12785 16294 16456 16346
rect 16508 16294 16520 16346
rect 16572 16294 16584 16346
rect 16636 16294 16648 16346
rect 16700 16294 16712 16346
rect 16764 16294 17940 16346
rect 2024 16272 17940 16294
rect 2024 15802 17940 15824
rect 2024 15750 3859 15802
rect 3911 15750 3923 15802
rect 3975 15750 3987 15802
rect 4039 15750 4051 15802
rect 4103 15750 4115 15802
rect 4167 15750 7838 15802
rect 7890 15750 7902 15802
rect 7954 15750 7966 15802
rect 8018 15750 8030 15802
rect 8082 15750 8094 15802
rect 8146 15750 11817 15802
rect 11869 15750 11881 15802
rect 11933 15750 11945 15802
rect 11997 15750 12009 15802
rect 12061 15750 12073 15802
rect 12125 15750 15796 15802
rect 15848 15750 15860 15802
rect 15912 15750 15924 15802
rect 15976 15750 15988 15802
rect 16040 15750 16052 15802
rect 16104 15750 17940 15802
rect 2024 15728 17940 15750
rect 2024 15258 17940 15280
rect 2024 15206 4519 15258
rect 4571 15206 4583 15258
rect 4635 15206 4647 15258
rect 4699 15206 4711 15258
rect 4763 15206 4775 15258
rect 4827 15206 8498 15258
rect 8550 15206 8562 15258
rect 8614 15206 8626 15258
rect 8678 15206 8690 15258
rect 8742 15206 8754 15258
rect 8806 15206 12477 15258
rect 12529 15206 12541 15258
rect 12593 15206 12605 15258
rect 12657 15206 12669 15258
rect 12721 15206 12733 15258
rect 12785 15206 16456 15258
rect 16508 15206 16520 15258
rect 16572 15206 16584 15258
rect 16636 15206 16648 15258
rect 16700 15206 16712 15258
rect 16764 15206 17940 15258
rect 2024 15184 17940 15206
rect 2024 14714 17940 14736
rect 2024 14662 3859 14714
rect 3911 14662 3923 14714
rect 3975 14662 3987 14714
rect 4039 14662 4051 14714
rect 4103 14662 4115 14714
rect 4167 14662 7838 14714
rect 7890 14662 7902 14714
rect 7954 14662 7966 14714
rect 8018 14662 8030 14714
rect 8082 14662 8094 14714
rect 8146 14662 11817 14714
rect 11869 14662 11881 14714
rect 11933 14662 11945 14714
rect 11997 14662 12009 14714
rect 12061 14662 12073 14714
rect 12125 14662 15796 14714
rect 15848 14662 15860 14714
rect 15912 14662 15924 14714
rect 15976 14662 15988 14714
rect 16040 14662 16052 14714
rect 16104 14662 17940 14714
rect 2024 14640 17940 14662
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 11514 14464 11520 14476
rect 10735 14436 11520 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 11054 14396 11060 14408
rect 10643 14368 11060 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 10965 14263 11023 14269
rect 10965 14229 10977 14263
rect 11011 14260 11023 14263
rect 11606 14260 11612 14272
rect 11011 14232 11612 14260
rect 11011 14229 11023 14232
rect 10965 14223 11023 14229
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 2024 14170 17940 14192
rect 2024 14118 4519 14170
rect 4571 14118 4583 14170
rect 4635 14118 4647 14170
rect 4699 14118 4711 14170
rect 4763 14118 4775 14170
rect 4827 14118 8498 14170
rect 8550 14118 8562 14170
rect 8614 14118 8626 14170
rect 8678 14118 8690 14170
rect 8742 14118 8754 14170
rect 8806 14118 12477 14170
rect 12529 14118 12541 14170
rect 12593 14118 12605 14170
rect 12657 14118 12669 14170
rect 12721 14118 12733 14170
rect 12785 14118 16456 14170
rect 16508 14118 16520 14170
rect 16572 14118 16584 14170
rect 16636 14118 16648 14170
rect 16700 14118 16712 14170
rect 16764 14118 17940 14170
rect 2024 14096 17940 14118
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 10689 14059 10747 14065
rect 10689 14056 10701 14059
rect 9548 14028 10701 14056
rect 9548 14016 9554 14028
rect 10689 14025 10701 14028
rect 10735 14025 10747 14059
rect 11238 14056 11244 14068
rect 10689 14019 10747 14025
rect 10888 14028 11244 14056
rect 10888 13988 10916 14028
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11514 14016 11520 14068
rect 11572 14016 11578 14068
rect 11608 14028 13400 14056
rect 11608 13988 11636 14028
rect 13081 13991 13139 13997
rect 13081 13988 13093 13991
rect 10428 13960 10916 13988
rect 10980 13960 11636 13988
rect 12406 13960 13093 13988
rect 8570 13880 8576 13932
rect 8628 13880 8634 13932
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 10134 13920 10140 13932
rect 9999 13892 10140 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13852 8723 13855
rect 9490 13852 9496 13864
rect 8711 13824 9496 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 9490 13812 9496 13824
rect 9548 13812 9554 13864
rect 9784 13852 9812 13883
rect 10134 13880 10140 13892
rect 10192 13920 10198 13932
rect 10428 13929 10456 13960
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 10192 13892 10241 13920
rect 10192 13880 10198 13892
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 10229 13883 10287 13889
rect 10413 13923 10471 13929
rect 10413 13889 10425 13923
rect 10459 13889 10471 13923
rect 10413 13883 10471 13889
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 9784 13824 10057 13852
rect 10045 13821 10057 13824
rect 10091 13852 10103 13855
rect 10594 13852 10600 13864
rect 10091 13824 10600 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 10980 13861 11008 13960
rect 11348 13929 11376 13960
rect 11333 13923 11391 13929
rect 11333 13889 11345 13923
rect 11379 13889 11391 13923
rect 11333 13883 11391 13889
rect 11425 13923 11483 13929
rect 11425 13889 11437 13923
rect 11471 13920 11483 13923
rect 12406 13920 12434 13960
rect 12820 13929 12848 13960
rect 13081 13957 13093 13960
rect 13127 13957 13139 13991
rect 13081 13951 13139 13957
rect 11471 13892 12434 13920
rect 12805 13923 12863 13929
rect 11471 13889 11483 13892
rect 11425 13883 11483 13889
rect 12805 13889 12817 13923
rect 12851 13889 12863 13923
rect 12805 13883 12863 13889
rect 10873 13855 10931 13861
rect 10873 13821 10885 13855
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 8941 13787 8999 13793
rect 8941 13753 8953 13787
rect 8987 13784 8999 13787
rect 9122 13784 9128 13796
rect 8987 13756 9128 13784
rect 8987 13753 8999 13756
rect 8941 13747 8999 13753
rect 9122 13744 9128 13756
rect 9180 13744 9186 13796
rect 9858 13676 9864 13728
rect 9916 13676 9922 13728
rect 10888 13716 10916 13815
rect 11072 13784 11100 13815
rect 11146 13812 11152 13864
rect 11204 13812 11210 13864
rect 11440 13852 11468 13883
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13265 13923 13323 13929
rect 13265 13920 13277 13923
rect 13044 13892 13277 13920
rect 13044 13880 13050 13892
rect 13265 13889 13277 13892
rect 13311 13889 13323 13923
rect 13265 13883 13323 13889
rect 13372 13920 13400 14028
rect 13998 13920 14004 13932
rect 13372 13892 14004 13920
rect 11256 13824 11468 13852
rect 11256 13784 11284 13824
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11756 13824 11805 13852
rect 11756 13812 11762 13824
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 11072 13756 11284 13784
rect 11808 13784 11836 13815
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12216 13824 12449 13852
rect 12216 13812 12222 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13372 13852 13400 13892
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 12943 13824 13400 13852
rect 13449 13855 13507 13861
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13449 13821 13461 13855
rect 13495 13821 13507 13855
rect 13449 13815 13507 13821
rect 13464 13784 13492 13815
rect 13722 13784 13728 13796
rect 11808 13756 13728 13784
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 11054 13716 11060 13728
rect 10888 13688 11060 13716
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 2024 13626 17940 13648
rect 2024 13574 3859 13626
rect 3911 13574 3923 13626
rect 3975 13574 3987 13626
rect 4039 13574 4051 13626
rect 4103 13574 4115 13626
rect 4167 13574 7838 13626
rect 7890 13574 7902 13626
rect 7954 13574 7966 13626
rect 8018 13574 8030 13626
rect 8082 13574 8094 13626
rect 8146 13574 11817 13626
rect 11869 13574 11881 13626
rect 11933 13574 11945 13626
rect 11997 13574 12009 13626
rect 12061 13574 12073 13626
rect 12125 13574 15796 13626
rect 15848 13574 15860 13626
rect 15912 13574 15924 13626
rect 15976 13574 15988 13626
rect 16040 13574 16052 13626
rect 16104 13574 17940 13626
rect 2024 13552 17940 13574
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8570 13512 8576 13524
rect 8527 13484 8576 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 8849 13515 8907 13521
rect 8849 13481 8861 13515
rect 8895 13481 8907 13515
rect 8849 13475 8907 13481
rect 10965 13515 11023 13521
rect 10965 13481 10977 13515
rect 11011 13512 11023 13515
rect 11146 13512 11152 13524
rect 11011 13484 11152 13512
rect 11011 13481 11023 13484
rect 10965 13475 11023 13481
rect 8864 13376 8892 13475
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 12986 13472 12992 13524
rect 13044 13472 13050 13524
rect 13357 13515 13415 13521
rect 13357 13481 13369 13515
rect 13403 13512 13415 13515
rect 13403 13484 13676 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 11054 13404 11060 13456
rect 11112 13404 11118 13456
rect 9030 13376 9036 13388
rect 8864 13348 9036 13376
rect 9030 13336 9036 13348
rect 9088 13376 9094 13388
rect 9088 13348 9260 13376
rect 9088 13336 9094 13348
rect 8938 13268 8944 13320
rect 8996 13308 9002 13320
rect 9232 13317 9260 13348
rect 9858 13336 9864 13388
rect 9916 13376 9922 13388
rect 11698 13376 11704 13388
rect 9916 13348 10732 13376
rect 9916 13336 9922 13348
rect 9217 13311 9275 13317
rect 8996 13280 9168 13308
rect 8996 13268 9002 13280
rect 9033 13243 9091 13249
rect 9033 13240 9045 13243
rect 6886 13212 9045 13240
rect 6730 13132 6736 13184
rect 6788 13172 6794 13184
rect 6886 13172 6914 13212
rect 9033 13209 9045 13212
rect 9079 13209 9091 13243
rect 9140 13240 9168 13280
rect 9217 13277 9229 13311
rect 9263 13277 9275 13311
rect 9217 13271 9275 13277
rect 9490 13268 9496 13320
rect 9548 13268 9554 13320
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 10192 13280 10425 13308
rect 10192 13268 10198 13280
rect 10413 13277 10425 13280
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 10594 13268 10600 13320
rect 10652 13268 10658 13320
rect 10704 13317 10732 13348
rect 10796 13348 11704 13376
rect 10796 13317 10824 13348
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 13372 13348 13553 13376
rect 13372 13320 13400 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 13648 13320 13676 13484
rect 13725 13379 13783 13385
rect 13725 13345 13737 13379
rect 13771 13345 13783 13379
rect 13725 13339 13783 13345
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13277 10839 13311
rect 11057 13311 11115 13317
rect 11057 13308 11069 13311
rect 10781 13271 10839 13277
rect 10980 13280 11069 13308
rect 10980 13249 11008 13280
rect 11057 13277 11069 13280
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 11238 13268 11244 13320
rect 11296 13268 11302 13320
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 13354 13268 13360 13320
rect 13412 13268 13418 13320
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13308 13507 13311
rect 13630 13308 13636 13320
rect 13495 13280 13636 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9140 13212 9413 13240
rect 9033 13203 9091 13209
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9401 13203 9459 13209
rect 10505 13243 10563 13249
rect 10505 13209 10517 13243
rect 10551 13240 10563 13243
rect 10965 13243 11023 13249
rect 10965 13240 10977 13243
rect 10551 13212 10977 13240
rect 10551 13209 10563 13212
rect 10505 13203 10563 13209
rect 10965 13209 10977 13212
rect 11011 13209 11023 13243
rect 13280 13240 13308 13268
rect 13740 13240 13768 13339
rect 13280 13212 13768 13240
rect 10965 13203 11023 13209
rect 6788 13144 6914 13172
rect 6788 13132 6794 13144
rect 13722 13132 13728 13184
rect 13780 13132 13786 13184
rect 2024 13082 17940 13104
rect 2024 13030 4519 13082
rect 4571 13030 4583 13082
rect 4635 13030 4647 13082
rect 4699 13030 4711 13082
rect 4763 13030 4775 13082
rect 4827 13030 8498 13082
rect 8550 13030 8562 13082
rect 8614 13030 8626 13082
rect 8678 13030 8690 13082
rect 8742 13030 8754 13082
rect 8806 13030 12477 13082
rect 12529 13030 12541 13082
rect 12593 13030 12605 13082
rect 12657 13030 12669 13082
rect 12721 13030 12733 13082
rect 12785 13030 16456 13082
rect 16508 13030 16520 13082
rect 16572 13030 16584 13082
rect 16636 13030 16648 13082
rect 16700 13030 16712 13082
rect 16764 13030 17940 13082
rect 2024 13008 17940 13030
rect 8938 12928 8944 12980
rect 8996 12928 9002 12980
rect 9030 12928 9036 12980
rect 9088 12928 9094 12980
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 13449 12971 13507 12977
rect 13449 12968 13461 12971
rect 13412 12940 13461 12968
rect 13412 12928 13418 12940
rect 13449 12937 13461 12940
rect 13495 12937 13507 12971
rect 13449 12931 13507 12937
rect 13630 12928 13636 12980
rect 13688 12928 13694 12980
rect 7374 12900 7380 12912
rect 2608 12872 7380 12900
rect 2608 12841 2636 12872
rect 7374 12860 7380 12872
rect 7432 12860 7438 12912
rect 8757 12903 8815 12909
rect 8757 12869 8769 12903
rect 8803 12900 8815 12903
rect 8803 12872 9444 12900
rect 8803 12869 8815 12872
rect 8757 12863 8815 12869
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 8570 12792 8576 12844
rect 8628 12792 8634 12844
rect 9416 12841 9444 12872
rect 13188 12872 16896 12900
rect 9217 12835 9275 12841
rect 9217 12801 9229 12835
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 10042 12832 10048 12844
rect 9447 12804 10048 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 6914 12764 6920 12776
rect 6871 12736 6920 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 8588 12764 8616 12792
rect 9232 12764 9260 12795
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 13188 12841 13216 12872
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 13538 12832 13544 12844
rect 13311 12804 13544 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 13722 12832 13728 12844
rect 13683 12804 13728 12832
rect 13722 12792 13728 12804
rect 13780 12832 13786 12844
rect 13832 12832 13860 12872
rect 16868 12841 16896 12872
rect 13780 12804 13860 12832
rect 16853 12835 16911 12841
rect 13780 12792 13786 12804
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 8588 12736 9260 12764
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16482 12764 16488 12776
rect 16347 12736 16488 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16482 12724 16488 12736
rect 16540 12764 16546 12776
rect 16577 12767 16635 12773
rect 16577 12764 16589 12767
rect 16540 12736 16589 12764
rect 16540 12724 16546 12736
rect 16577 12733 16589 12736
rect 16623 12733 16635 12767
rect 16577 12727 16635 12733
rect 7098 12656 7104 12708
rect 7156 12656 7162 12708
rect 2406 12588 2412 12640
rect 2464 12588 2470 12640
rect 2024 12538 17940 12560
rect 2024 12486 3859 12538
rect 3911 12486 3923 12538
rect 3975 12486 3987 12538
rect 4039 12486 4051 12538
rect 4103 12486 4115 12538
rect 4167 12486 7838 12538
rect 7890 12486 7902 12538
rect 7954 12486 7966 12538
rect 8018 12486 8030 12538
rect 8082 12486 8094 12538
rect 8146 12486 11817 12538
rect 11869 12486 11881 12538
rect 11933 12486 11945 12538
rect 11997 12486 12009 12538
rect 12061 12486 12073 12538
rect 12125 12486 15796 12538
rect 15848 12486 15860 12538
rect 15912 12486 15924 12538
rect 15976 12486 15988 12538
rect 16040 12486 16052 12538
rect 16104 12486 17940 12538
rect 2024 12464 17940 12486
rect 6914 12384 6920 12436
rect 6972 12384 6978 12436
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 7156 12396 7297 12424
rect 7156 12384 7162 12396
rect 7285 12393 7297 12396
rect 7331 12393 7343 12427
rect 7285 12387 7343 12393
rect 7374 12384 7380 12436
rect 7432 12384 7438 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 8757 12427 8815 12433
rect 8757 12424 8769 12427
rect 8628 12396 8769 12424
rect 8628 12384 8634 12396
rect 8757 12393 8769 12396
rect 8803 12393 8815 12427
rect 8757 12387 8815 12393
rect 10134 12384 10140 12436
rect 10192 12384 10198 12436
rect 12069 12427 12127 12433
rect 12069 12393 12081 12427
rect 12115 12424 12127 12427
rect 12158 12424 12164 12436
rect 12115 12396 12164 12424
rect 12115 12393 12127 12396
rect 12069 12387 12127 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12424 12587 12427
rect 12802 12424 12808 12436
rect 12575 12396 12808 12424
rect 12575 12393 12587 12396
rect 12529 12387 12587 12393
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 8941 12359 8999 12365
rect 8941 12356 8953 12359
rect 6656 12328 8953 12356
rect 6656 12297 6684 12328
rect 8941 12325 8953 12328
rect 8987 12325 8999 12359
rect 8941 12319 8999 12325
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12288 7527 12291
rect 7650 12288 7656 12300
rect 7515 12260 7656 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 8619 12260 9352 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 9324 12232 9352 12260
rect 9398 12248 9404 12300
rect 9456 12248 9462 12300
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 10008 12260 10517 12288
rect 10008 12248 10014 12260
rect 10505 12257 10517 12260
rect 10551 12288 10563 12291
rect 13814 12288 13820 12300
rect 10551 12260 13820 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 6362 12180 6368 12232
rect 6420 12220 6426 12232
rect 6549 12223 6607 12229
rect 6549 12220 6561 12223
rect 6420 12192 6561 12220
rect 6420 12180 6426 12192
rect 6549 12189 6561 12192
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 8202 12220 8208 12232
rect 7239 12192 8208 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 9214 12220 9220 12232
rect 9171 12192 9220 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 8496 12152 8524 12183
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 9306 12180 9312 12232
rect 9364 12180 9370 12232
rect 9030 12152 9036 12164
rect 8496 12124 9036 12152
rect 9030 12112 9036 12124
rect 9088 12152 9094 12164
rect 9416 12152 9444 12248
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12220 10471 12223
rect 10686 12220 10692 12232
rect 10459 12192 10692 12220
rect 10459 12189 10471 12192
rect 10413 12183 10471 12189
rect 10686 12180 10692 12192
rect 10744 12220 10750 12232
rect 11330 12220 11336 12232
rect 10744 12192 11336 12220
rect 10744 12180 10750 12192
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 9088 12124 9444 12152
rect 9088 12112 9094 12124
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 11992 12084 12020 12183
rect 12250 12180 12256 12232
rect 12308 12180 12314 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 13170 12220 13176 12232
rect 12391 12192 13176 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 8260 12056 12020 12084
rect 8260 12044 8266 12056
rect 2024 11994 17940 12016
rect 2024 11942 4519 11994
rect 4571 11942 4583 11994
rect 4635 11942 4647 11994
rect 4699 11942 4711 11994
rect 4763 11942 4775 11994
rect 4827 11942 8498 11994
rect 8550 11942 8562 11994
rect 8614 11942 8626 11994
rect 8678 11942 8690 11994
rect 8742 11942 8754 11994
rect 8806 11942 12477 11994
rect 12529 11942 12541 11994
rect 12593 11942 12605 11994
rect 12657 11942 12669 11994
rect 12721 11942 12733 11994
rect 12785 11942 16456 11994
rect 16508 11942 16520 11994
rect 16572 11942 16584 11994
rect 16636 11942 16648 11994
rect 16700 11942 16712 11994
rect 16764 11942 17940 11994
rect 2024 11920 17940 11942
rect 9306 11840 9312 11892
rect 9364 11880 9370 11892
rect 9769 11883 9827 11889
rect 9769 11880 9781 11883
rect 9364 11852 9781 11880
rect 9364 11840 9370 11852
rect 9769 11849 9781 11852
rect 9815 11849 9827 11883
rect 9769 11843 9827 11849
rect 11422 11840 11428 11892
rect 11480 11880 11486 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11480 11852 11805 11880
rect 11480 11840 11486 11852
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 12250 11840 12256 11892
rect 12308 11880 12314 11892
rect 12437 11883 12495 11889
rect 12437 11880 12449 11883
rect 12308 11852 12449 11880
rect 12308 11840 12314 11852
rect 12437 11849 12449 11852
rect 12483 11849 12495 11883
rect 12437 11843 12495 11849
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 12860 11852 13124 11880
rect 12860 11840 12866 11852
rect 9214 11772 9220 11824
rect 9272 11812 9278 11824
rect 11054 11812 11060 11824
rect 9272 11784 11060 11812
rect 9272 11772 9278 11784
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11744 2651 11747
rect 8662 11744 8668 11756
rect 2639 11716 8668 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9950 11704 9956 11756
rect 10008 11704 10014 11756
rect 10244 11753 10272 11784
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 11149 11815 11207 11821
rect 11149 11781 11161 11815
rect 11195 11812 11207 11815
rect 13096 11812 13124 11852
rect 13170 11840 13176 11892
rect 13228 11840 13234 11892
rect 13814 11840 13820 11892
rect 13872 11840 13878 11892
rect 13262 11812 13268 11824
rect 11195 11784 11376 11812
rect 11195 11781 11207 11784
rect 11149 11775 11207 11781
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 10152 11676 10180 11707
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 10594 11744 10600 11756
rect 10376 11716 10600 11744
rect 10376 11704 10382 11716
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 10870 11704 10876 11756
rect 10928 11704 10934 11756
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 10686 11676 10692 11688
rect 10152 11648 10692 11676
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 1210 11568 1216 11620
rect 1268 11608 1274 11620
rect 2409 11611 2467 11617
rect 2409 11608 2421 11611
rect 1268 11580 2421 11608
rect 1268 11568 1274 11580
rect 2409 11577 2421 11580
rect 2455 11577 2467 11611
rect 10980 11608 11008 11707
rect 11238 11704 11244 11756
rect 11296 11704 11302 11756
rect 11348 11753 11376 11784
rect 11532 11784 13032 11812
rect 13096 11784 13268 11812
rect 11532 11753 11560 11784
rect 13004 11756 13032 11784
rect 13262 11772 13268 11784
rect 13320 11812 13326 11824
rect 17402 11812 17408 11824
rect 13320 11784 17408 11812
rect 13320 11772 13326 11784
rect 11333 11747 11391 11753
rect 11333 11713 11345 11747
rect 11379 11713 11391 11747
rect 11333 11707 11391 11713
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 12621 11747 12679 11753
rect 12621 11744 12633 11747
rect 12492 11716 12633 11744
rect 12492 11704 12498 11716
rect 12621 11713 12633 11716
rect 12667 11713 12679 11747
rect 12621 11707 12679 11713
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11713 12771 11747
rect 12713 11707 12771 11713
rect 12728 11676 12756 11707
rect 12802 11704 12808 11756
rect 12860 11704 12866 11756
rect 12986 11704 12992 11756
rect 13044 11704 13050 11756
rect 13078 11704 13084 11756
rect 13136 11704 13142 11756
rect 13170 11704 13176 11756
rect 13228 11744 13234 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 13228 11716 13369 11744
rect 13228 11704 13234 11716
rect 13357 11713 13369 11716
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 13446 11704 13452 11756
rect 13504 11704 13510 11756
rect 13740 11753 13768 11784
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11713 13783 11747
rect 13725 11707 13783 11713
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 12894 11676 12900 11688
rect 12728 11648 12900 11676
rect 12894 11636 12900 11648
rect 12952 11676 12958 11688
rect 14016 11676 14044 11707
rect 14274 11704 14280 11756
rect 14332 11704 14338 11756
rect 17310 11704 17316 11756
rect 17368 11704 17374 11756
rect 12952 11648 13676 11676
rect 14016 11648 14872 11676
rect 12952 11636 12958 11648
rect 13170 11608 13176 11620
rect 10980 11580 13176 11608
rect 2409 11571 2467 11577
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 13648 11617 13676 11648
rect 14844 11620 14872 11648
rect 13633 11611 13691 11617
rect 13633 11577 13645 11611
rect 13679 11608 13691 11611
rect 13722 11608 13728 11620
rect 13679 11580 13728 11608
rect 13679 11577 13691 11580
rect 13633 11571 13691 11577
rect 13722 11568 13728 11580
rect 13780 11608 13786 11620
rect 14093 11611 14151 11617
rect 14093 11608 14105 11611
rect 13780 11580 14105 11608
rect 13780 11568 13786 11580
rect 14093 11577 14105 11580
rect 14139 11577 14151 11611
rect 14093 11571 14151 11577
rect 14182 11568 14188 11620
rect 14240 11568 14246 11620
rect 14826 11568 14832 11620
rect 14884 11608 14890 11620
rect 17129 11611 17187 11617
rect 17129 11608 17141 11611
rect 14884 11580 17141 11608
rect 14884 11568 14890 11580
rect 17129 11577 17141 11580
rect 17175 11577 17187 11611
rect 17129 11571 17187 11577
rect 2024 11450 17940 11472
rect 2024 11398 3859 11450
rect 3911 11398 3923 11450
rect 3975 11398 3987 11450
rect 4039 11398 4051 11450
rect 4103 11398 4115 11450
rect 4167 11398 7838 11450
rect 7890 11398 7902 11450
rect 7954 11398 7966 11450
rect 8018 11398 8030 11450
rect 8082 11398 8094 11450
rect 8146 11398 11817 11450
rect 11869 11398 11881 11450
rect 11933 11398 11945 11450
rect 11997 11398 12009 11450
rect 12061 11398 12073 11450
rect 12125 11398 15796 11450
rect 15848 11398 15860 11450
rect 15912 11398 15924 11450
rect 15976 11398 15988 11450
rect 16040 11398 16052 11450
rect 16104 11398 17940 11450
rect 2024 11376 17940 11398
rect 7650 11296 7656 11348
rect 7708 11296 7714 11348
rect 8662 11296 8668 11348
rect 8720 11296 8726 11348
rect 9122 11296 9128 11348
rect 9180 11296 9186 11348
rect 10870 11296 10876 11348
rect 10928 11336 10934 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10928 11308 10977 11336
rect 10928 11296 10934 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 12529 11339 12587 11345
rect 12529 11305 12541 11339
rect 12575 11336 12587 11339
rect 13446 11336 13452 11348
rect 12575 11308 13452 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13538 11296 13544 11348
rect 13596 11296 13602 11348
rect 14274 11336 14280 11348
rect 13740 11308 14280 11336
rect 2501 11271 2559 11277
rect 2501 11237 2513 11271
rect 2547 11268 2559 11271
rect 5902 11268 5908 11280
rect 2547 11240 5908 11268
rect 2547 11237 2559 11240
rect 2501 11231 2559 11237
rect 5902 11228 5908 11240
rect 5960 11228 5966 11280
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 8202 11200 8208 11212
rect 7156 11172 8208 11200
rect 7156 11160 7162 11172
rect 8202 11160 8208 11172
rect 8260 11200 8266 11212
rect 8260 11172 9260 11200
rect 8260 11160 8266 11172
rect 2314 11092 2320 11144
rect 2372 11092 2378 11144
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 6362 11024 6368 11076
rect 6420 11064 6426 11076
rect 7300 11064 7328 11095
rect 7374 11092 7380 11144
rect 7432 11092 7438 11144
rect 8846 11092 8852 11144
rect 8904 11092 8910 11144
rect 8938 11092 8944 11144
rect 8996 11092 9002 11144
rect 9232 11141 9260 11172
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 12158 11200 12164 11212
rect 11112 11172 12164 11200
rect 11112 11160 11118 11172
rect 12158 11160 12164 11172
rect 12216 11200 12222 11212
rect 13740 11200 13768 11308
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 17402 11296 17408 11348
rect 17460 11296 17466 11348
rect 14182 11200 14188 11212
rect 12216 11172 13768 11200
rect 12216 11160 12222 11172
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 10686 11092 10692 11144
rect 10744 11092 10750 11144
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11132 12863 11135
rect 12894 11132 12900 11144
rect 12851 11104 12900 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13740 11141 13768 11172
rect 13924 11172 14188 11200
rect 13924 11144 13952 11172
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 14292 11200 14320 11296
rect 14829 11271 14887 11277
rect 14829 11237 14841 11271
rect 14875 11268 14887 11271
rect 14918 11268 14924 11280
rect 14875 11240 14924 11268
rect 14875 11237 14887 11240
rect 14829 11231 14887 11237
rect 14918 11228 14924 11240
rect 14976 11228 14982 11280
rect 14292 11172 14688 11200
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11101 13783 11135
rect 13725 11095 13783 11101
rect 13906 11092 13912 11144
rect 13964 11092 13970 11144
rect 14001 11135 14059 11141
rect 14001 11101 14013 11135
rect 14047 11132 14059 11135
rect 14200 11132 14228 11160
rect 14660 11141 14688 11172
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 14047 11104 14136 11132
rect 14200 11104 14565 11132
rect 14047 11101 14059 11104
rect 14001 11095 14059 11101
rect 6420 11036 7328 11064
rect 7392 11064 7420 11092
rect 9766 11064 9772 11076
rect 7392 11036 9772 11064
rect 6420 11024 6426 11036
rect 9766 11024 9772 11036
rect 9824 11064 9830 11076
rect 10965 11067 11023 11073
rect 10965 11064 10977 11067
rect 9824 11036 10977 11064
rect 9824 11024 9830 11036
rect 10965 11033 10977 11036
rect 11011 11064 11023 11067
rect 12529 11067 12587 11073
rect 12529 11064 12541 11067
rect 11011 11036 12541 11064
rect 11011 11033 11023 11036
rect 10965 11027 11023 11033
rect 12529 11033 12541 11036
rect 12575 11064 12587 11067
rect 13538 11064 13544 11076
rect 12575 11036 13544 11064
rect 12575 11033 12587 11036
rect 12529 11027 12587 11033
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 14108 11073 14136 11104
rect 14292 11073 14320 11104
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 14553 11095 14611 11101
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 14093 11067 14151 11073
rect 14093 11033 14105 11067
rect 14139 11033 14151 11067
rect 14292 11067 14351 11073
rect 14292 11036 14305 11067
rect 14093 11027 14151 11033
rect 14293 11033 14305 11036
rect 14339 11033 14351 11067
rect 14844 11064 14872 11092
rect 14293 11027 14351 11033
rect 14384 11036 14872 11064
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 9858 10996 9864 11008
rect 6696 10968 9864 10996
rect 6696 10956 6702 10968
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 10778 10996 10784 11008
rect 10376 10968 10784 10996
rect 10376 10956 10382 10968
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 12713 10999 12771 11005
rect 12713 10965 12725 10999
rect 12759 10996 12771 10999
rect 12802 10996 12808 11008
rect 12759 10968 12808 10996
rect 12759 10965 12771 10968
rect 12713 10959 12771 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14108 10996 14136 11027
rect 14384 10996 14412 11036
rect 17494 11024 17500 11076
rect 17552 11024 17558 11076
rect 13872 10968 14412 10996
rect 13872 10956 13878 10968
rect 14458 10956 14464 11008
rect 14516 10956 14522 11008
rect 2024 10906 17940 10928
rect 2024 10854 4519 10906
rect 4571 10854 4583 10906
rect 4635 10854 4647 10906
rect 4699 10854 4711 10906
rect 4763 10854 4775 10906
rect 4827 10854 8498 10906
rect 8550 10854 8562 10906
rect 8614 10854 8626 10906
rect 8678 10854 8690 10906
rect 8742 10854 8754 10906
rect 8806 10854 12477 10906
rect 12529 10854 12541 10906
rect 12593 10854 12605 10906
rect 12657 10854 12669 10906
rect 12721 10854 12733 10906
rect 12785 10854 16456 10906
rect 16508 10854 16520 10906
rect 16572 10854 16584 10906
rect 16636 10854 16648 10906
rect 16700 10854 16712 10906
rect 16764 10854 17940 10906
rect 2024 10832 17940 10854
rect 6362 10752 6368 10804
rect 6420 10752 6426 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 7064 10764 7113 10792
rect 7064 10752 7070 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 7101 10755 7159 10761
rect 8128 10764 9597 10792
rect 7653 10727 7711 10733
rect 7653 10724 7665 10727
rect 6472 10696 7665 10724
rect 6472 10668 6500 10696
rect 7653 10693 7665 10696
rect 7699 10693 7711 10727
rect 7653 10687 7711 10693
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 2639 10628 6009 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 5997 10625 6009 10628
rect 6043 10656 6055 10659
rect 6454 10656 6460 10668
rect 6043 10628 6460 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 6963 10628 7297 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7466 10616 7472 10668
rect 7524 10616 7530 10668
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 1118 10548 1124 10600
rect 1176 10588 1182 10600
rect 2317 10591 2375 10597
rect 2317 10588 2329 10591
rect 1176 10560 2329 10588
rect 1176 10548 1182 10560
rect 2317 10557 2329 10560
rect 2363 10557 2375 10591
rect 2317 10551 2375 10557
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 7576 10588 7604 10619
rect 7742 10616 7748 10668
rect 7800 10665 7806 10668
rect 8128 10665 8156 10764
rect 9030 10724 9036 10736
rect 8220 10696 9036 10724
rect 7800 10659 7829 10665
rect 7817 10625 7829 10659
rect 7800 10619 7829 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8113 10659 8171 10665
rect 8113 10656 8125 10659
rect 7975 10628 8125 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8113 10625 8125 10628
rect 8159 10625 8171 10659
rect 8113 10619 8171 10625
rect 7800 10616 7806 10619
rect 8220 10597 8248 10696
rect 9030 10684 9036 10696
rect 9088 10684 9094 10736
rect 9140 10733 9168 10764
rect 9585 10761 9597 10764
rect 9631 10792 9643 10795
rect 10042 10792 10048 10804
rect 9631 10764 10048 10792
rect 9631 10761 9643 10764
rect 9585 10755 9643 10761
rect 10042 10752 10048 10764
rect 10100 10792 10106 10804
rect 10100 10764 10732 10792
rect 10100 10752 10106 10764
rect 10704 10733 10732 10764
rect 10778 10752 10784 10804
rect 10836 10752 10842 10804
rect 10965 10795 11023 10801
rect 10965 10761 10977 10795
rect 11011 10792 11023 10795
rect 11238 10792 11244 10804
rect 11011 10764 11244 10792
rect 11011 10761 11023 10764
rect 10965 10755 11023 10761
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 13078 10792 13084 10804
rect 11931 10764 13084 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10693 9183 10727
rect 9953 10727 10011 10733
rect 9953 10724 9965 10727
rect 9125 10687 9183 10693
rect 9416 10696 9965 10724
rect 8329 10659 8387 10665
rect 8329 10656 8341 10659
rect 8312 10625 8341 10656
rect 8375 10625 8387 10659
rect 8312 10619 8387 10625
rect 5960 10560 7604 10588
rect 8205 10591 8263 10597
rect 5960 10548 5966 10560
rect 8205 10557 8217 10591
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8312 10520 8340 10619
rect 8478 10616 8484 10668
rect 8536 10616 8542 10668
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8628 10628 8953 10656
rect 8628 10616 8634 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9048 10588 9076 10684
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9416 10665 9444 10696
rect 9953 10693 9965 10696
rect 9999 10693 10011 10727
rect 9953 10687 10011 10693
rect 10689 10727 10747 10733
rect 10689 10693 10701 10727
rect 10735 10693 10747 10727
rect 10796 10724 10824 10752
rect 11609 10727 11667 10733
rect 11609 10724 11621 10727
rect 10796 10696 11621 10724
rect 10689 10687 10747 10693
rect 11609 10693 11621 10696
rect 11655 10693 11667 10727
rect 11609 10687 11667 10693
rect 13722 10684 13728 10736
rect 13780 10724 13786 10736
rect 13780 10696 15424 10724
rect 13780 10684 13786 10696
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9508 10588 9536 10619
rect 9766 10616 9772 10668
rect 9824 10616 9830 10668
rect 9858 10616 9864 10668
rect 9916 10616 9922 10668
rect 10042 10616 10048 10668
rect 10100 10616 10106 10668
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10502 10665 10508 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10284 10628 10333 10656
rect 10284 10616 10290 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10469 10659 10508 10665
rect 10469 10625 10481 10659
rect 10469 10619 10508 10625
rect 10502 10616 10508 10619
rect 10560 10616 10566 10668
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10656 10655 10659
rect 10827 10659 10885 10665
rect 10643 10628 10732 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 9048 10560 9536 10588
rect 9769 10523 9827 10529
rect 9769 10520 9781 10523
rect 8312 10492 9781 10520
rect 9769 10489 9781 10492
rect 9815 10489 9827 10523
rect 9769 10483 9827 10489
rect 10704 10520 10732 10628
rect 10827 10625 10839 10659
rect 10873 10656 10885 10659
rect 10873 10628 11008 10656
rect 10873 10625 10885 10628
rect 10827 10619 10885 10625
rect 10980 10588 11008 10628
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11241 10659 11299 10665
rect 11241 10656 11253 10659
rect 11112 10628 11253 10656
rect 11112 10616 11118 10628
rect 11241 10625 11253 10628
rect 11287 10625 11299 10659
rect 11241 10619 11299 10625
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11388 10628 11433 10656
rect 11388 10616 11394 10628
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 11706 10659 11764 10665
rect 11706 10625 11718 10659
rect 11752 10656 11764 10659
rect 12618 10656 12624 10668
rect 11752 10628 12624 10656
rect 11752 10625 11764 10628
rect 11706 10619 11764 10625
rect 11716 10588 11744 10619
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 14458 10616 14464 10668
rect 14516 10656 14522 10668
rect 14844 10665 14872 10696
rect 14553 10659 14611 10665
rect 14553 10656 14565 10659
rect 14516 10628 14565 10656
rect 14516 10616 14522 10628
rect 14553 10625 14565 10628
rect 14599 10625 14611 10659
rect 14553 10619 14611 10625
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10625 14887 10659
rect 14829 10619 14887 10625
rect 10980 10560 11744 10588
rect 11606 10520 11612 10532
rect 10704 10492 11612 10520
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 8478 10452 8484 10464
rect 7708 10424 8484 10452
rect 7708 10412 7714 10424
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 8570 10412 8576 10464
rect 8628 10452 8634 10464
rect 8665 10455 8723 10461
rect 8665 10452 8677 10455
rect 8628 10424 8677 10452
rect 8628 10412 8634 10424
rect 8665 10421 8677 10424
rect 8711 10421 8723 10455
rect 8665 10415 8723 10421
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 10704 10452 10732 10492
rect 11606 10480 11612 10492
rect 11664 10480 11670 10532
rect 14568 10520 14596 10619
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14976 10628 15117 10656
rect 14976 10616 14982 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 14936 10588 14964 10616
rect 15396 10597 15424 10696
rect 17402 10616 17408 10668
rect 17460 10616 17466 10668
rect 14691 10560 14964 10588
rect 15381 10591 15439 10597
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 15381 10557 15393 10591
rect 15427 10557 15439 10591
rect 15381 10551 15439 10557
rect 14826 10520 14832 10532
rect 14568 10492 14832 10520
rect 14826 10480 14832 10492
rect 14884 10520 14890 10532
rect 15197 10523 15255 10529
rect 15197 10520 15209 10523
rect 14884 10492 15209 10520
rect 14884 10480 14890 10492
rect 15197 10489 15209 10492
rect 15243 10489 15255 10523
rect 15396 10520 15424 10551
rect 15470 10520 15476 10532
rect 15396 10492 15476 10520
rect 15197 10483 15255 10489
rect 15470 10480 15476 10492
rect 15528 10520 15534 10532
rect 17221 10523 17279 10529
rect 17221 10520 17233 10523
rect 15528 10492 17233 10520
rect 15528 10480 15534 10492
rect 17221 10489 17233 10492
rect 17267 10489 17279 10523
rect 17221 10483 17279 10489
rect 8904 10424 10732 10452
rect 8904 10412 8910 10424
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12802 10452 12808 10464
rect 12492 10424 12808 10452
rect 12492 10412 12498 10424
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 15010 10412 15016 10464
rect 15068 10412 15074 10464
rect 15102 10412 15108 10464
rect 15160 10412 15166 10464
rect 2024 10362 17940 10384
rect 2024 10310 3859 10362
rect 3911 10310 3923 10362
rect 3975 10310 3987 10362
rect 4039 10310 4051 10362
rect 4103 10310 4115 10362
rect 4167 10310 7838 10362
rect 7890 10310 7902 10362
rect 7954 10310 7966 10362
rect 8018 10310 8030 10362
rect 8082 10310 8094 10362
rect 8146 10310 11817 10362
rect 11869 10310 11881 10362
rect 11933 10310 11945 10362
rect 11997 10310 12009 10362
rect 12061 10310 12073 10362
rect 12125 10310 15796 10362
rect 15848 10310 15860 10362
rect 15912 10310 15924 10362
rect 15976 10310 15988 10362
rect 16040 10310 16052 10362
rect 16104 10310 17940 10362
rect 2024 10288 17940 10310
rect 5902 10208 5908 10260
rect 5960 10248 5966 10260
rect 6917 10251 6975 10257
rect 6917 10248 6929 10251
rect 5960 10220 6929 10248
rect 5960 10208 5966 10220
rect 6917 10217 6929 10220
rect 6963 10217 6975 10251
rect 6917 10211 6975 10217
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7190 10248 7196 10260
rect 7055 10220 7196 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 8938 10208 8944 10260
rect 8996 10248 9002 10260
rect 9217 10251 9275 10257
rect 9217 10248 9229 10251
rect 8996 10220 9229 10248
rect 8996 10208 9002 10220
rect 9217 10217 9229 10220
rect 9263 10217 9275 10251
rect 9217 10211 9275 10217
rect 10226 10208 10232 10260
rect 10284 10208 10290 10260
rect 11054 10208 11060 10260
rect 11112 10208 11118 10260
rect 12434 10248 12440 10260
rect 11164 10220 12440 10248
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 8536 10152 10456 10180
rect 8536 10140 8542 10152
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 8386 10112 8392 10124
rect 7147 10084 8392 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 10428 10121 10456 10152
rect 10502 10140 10508 10192
rect 10560 10180 10566 10192
rect 10560 10152 10916 10180
rect 10560 10140 10566 10152
rect 10413 10115 10471 10121
rect 8496 10084 8984 10112
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6512 10016 6837 10044
rect 6512 10004 6518 10016
rect 6825 10013 6837 10016
rect 6871 10044 6883 10047
rect 8496 10044 8524 10084
rect 6871 10016 8524 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 8721 10047 8779 10053
rect 8721 10013 8733 10047
rect 8767 10044 8779 10047
rect 8767 10013 8800 10044
rect 8721 10007 8800 10013
rect 8772 9976 8800 10007
rect 8846 10004 8852 10056
rect 8904 10004 8910 10056
rect 8956 10053 8984 10084
rect 10413 10081 10425 10115
rect 10459 10112 10471 10115
rect 10778 10112 10784 10124
rect 10459 10084 10784 10112
rect 10459 10081 10471 10084
rect 10413 10075 10471 10081
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 10888 10112 10916 10152
rect 11164 10112 11192 10220
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14884 10220 15424 10248
rect 14884 10208 14890 10220
rect 11330 10140 11336 10192
rect 11388 10180 11394 10192
rect 12526 10180 12532 10192
rect 11388 10152 12532 10180
rect 11388 10140 11394 10152
rect 12526 10140 12532 10152
rect 12584 10180 12590 10192
rect 13722 10180 13728 10192
rect 12584 10152 13728 10180
rect 12584 10140 12590 10152
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 14918 10140 14924 10192
rect 14976 10180 14982 10192
rect 15396 10189 15424 10220
rect 15381 10183 15439 10189
rect 14976 10152 15332 10180
rect 14976 10140 14982 10152
rect 10888 10084 11192 10112
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9079 10047 9137 10053
rect 9079 10013 9091 10047
rect 9125 10044 9137 10047
rect 9398 10044 9404 10056
rect 9125 10016 9404 10044
rect 9125 10013 9137 10016
rect 9079 10007 9137 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 10597 10047 10655 10053
rect 10597 10013 10609 10047
rect 10643 10013 10655 10047
rect 10597 10007 10655 10013
rect 10318 9976 10324 9988
rect 8772 9948 10324 9976
rect 10318 9936 10324 9948
rect 10376 9976 10382 9988
rect 10612 9976 10640 10007
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 10888 10053 10916 10084
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10013 10931 10047
rect 10873 10007 10931 10013
rect 10962 10004 10968 10056
rect 11020 10044 11026 10056
rect 11348 10053 11376 10140
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 11664 10084 11836 10112
rect 11664 10072 11670 10084
rect 11057 10047 11115 10053
rect 11057 10044 11069 10047
rect 11020 10016 11069 10044
rect 11020 10004 11026 10016
rect 11057 10013 11069 10016
rect 11103 10044 11115 10047
rect 11149 10047 11207 10053
rect 11149 10044 11161 10047
rect 11103 10016 11161 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 11149 10013 11161 10016
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 10376 9948 10640 9976
rect 11241 9979 11299 9985
rect 10376 9936 10382 9948
rect 10520 9920 10548 9948
rect 11241 9945 11253 9979
rect 11287 9976 11299 9979
rect 11440 9976 11468 10007
rect 11287 9948 11468 9976
rect 11532 9976 11560 10007
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 11808 10053 11836 10084
rect 11974 10072 11980 10124
rect 12032 10072 12038 10124
rect 13357 10115 13415 10121
rect 13357 10112 13369 10115
rect 12452 10084 13369 10112
rect 11793 10047 11851 10053
rect 11793 10013 11805 10047
rect 11839 10044 11851 10047
rect 12250 10044 12256 10056
rect 11839 10016 12256 10044
rect 11839 10013 11851 10016
rect 11793 10007 11851 10013
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 12452 10053 12480 10084
rect 13357 10081 13369 10084
rect 13403 10112 13415 10115
rect 15102 10112 15108 10124
rect 13403 10084 13860 10112
rect 13403 10081 13415 10084
rect 13357 10075 13415 10081
rect 13832 10056 13860 10084
rect 14844 10084 15108 10112
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 12161 9979 12219 9985
rect 12161 9976 12173 9979
rect 11532 9948 12173 9976
rect 11287 9945 11299 9948
rect 11241 9939 11299 9945
rect 12161 9945 12173 9948
rect 12207 9945 12219 9979
rect 12161 9939 12219 9945
rect 12360 9920 12388 10007
rect 12526 10004 12532 10056
rect 12584 10004 12590 10056
rect 12802 10004 12808 10056
rect 12860 10004 12866 10056
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10013 13231 10047
rect 13449 10047 13507 10053
rect 13449 10044 13461 10047
rect 13173 10007 13231 10013
rect 13372 10016 13461 10044
rect 12618 9936 12624 9988
rect 12676 9985 12682 9988
rect 12676 9979 12725 9985
rect 12676 9945 12679 9979
rect 12713 9976 12725 9979
rect 12713 9948 13124 9976
rect 12713 9945 12725 9948
rect 12676 9939 12725 9945
rect 12676 9936 12682 9939
rect 13096 9920 13124 9948
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7742 9908 7748 9920
rect 7616 9880 7748 9908
rect 7616 9868 7622 9880
rect 7742 9868 7748 9880
rect 7800 9908 7806 9920
rect 8846 9908 8852 9920
rect 7800 9880 8852 9908
rect 7800 9868 7806 9880
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 10502 9868 10508 9920
rect 10560 9868 10566 9920
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 12342 9908 12348 9920
rect 10836 9880 12348 9908
rect 10836 9868 10842 9880
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 12897 9911 12955 9917
rect 12897 9908 12909 9911
rect 12860 9880 12909 9908
rect 12860 9868 12866 9880
rect 12897 9877 12909 9880
rect 12943 9877 12955 9911
rect 12897 9871 12955 9877
rect 13078 9868 13084 9920
rect 13136 9868 13142 9920
rect 13188 9908 13216 10007
rect 13262 9936 13268 9988
rect 13320 9976 13326 9988
rect 13372 9976 13400 10016
rect 13449 10013 13461 10016
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 13722 10004 13728 10056
rect 13780 10004 13786 10056
rect 13814 10004 13820 10056
rect 13872 10004 13878 10056
rect 14844 10053 14872 10084
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15304 10121 15332 10152
rect 15381 10149 15393 10183
rect 15427 10149 15439 10183
rect 15381 10143 15439 10149
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 13740 9976 13768 10004
rect 13320 9948 13768 9976
rect 14660 9976 14688 10007
rect 15010 10004 15016 10056
rect 15068 10004 15074 10056
rect 15194 10004 15200 10056
rect 15252 10004 15258 10056
rect 15470 10004 15476 10056
rect 15528 10004 15534 10056
rect 17310 10004 17316 10056
rect 17368 10004 17374 10056
rect 15028 9976 15056 10004
rect 14660 9948 15056 9976
rect 13320 9936 13326 9948
rect 13639 9911 13697 9917
rect 13639 9908 13651 9911
rect 13188 9880 13651 9908
rect 13639 9877 13651 9880
rect 13685 9877 13697 9911
rect 13639 9871 13697 9877
rect 14734 9868 14740 9920
rect 14792 9868 14798 9920
rect 15654 9868 15660 9920
rect 15712 9868 15718 9920
rect 17494 9868 17500 9920
rect 17552 9868 17558 9920
rect 2024 9818 17940 9840
rect 2024 9766 4519 9818
rect 4571 9766 4583 9818
rect 4635 9766 4647 9818
rect 4699 9766 4711 9818
rect 4763 9766 4775 9818
rect 4827 9766 8498 9818
rect 8550 9766 8562 9818
rect 8614 9766 8626 9818
rect 8678 9766 8690 9818
rect 8742 9766 8754 9818
rect 8806 9766 12477 9818
rect 12529 9766 12541 9818
rect 12593 9766 12605 9818
rect 12657 9766 12669 9818
rect 12721 9766 12733 9818
rect 12785 9766 16456 9818
rect 16508 9766 16520 9818
rect 16572 9766 16584 9818
rect 16636 9766 16648 9818
rect 16700 9766 16712 9818
rect 16764 9766 17940 9818
rect 2024 9744 17940 9766
rect 10597 9707 10655 9713
rect 10597 9673 10609 9707
rect 10643 9704 10655 9707
rect 10686 9704 10692 9716
rect 10643 9676 10692 9704
rect 10643 9673 10655 9676
rect 10597 9667 10655 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11974 9664 11980 9716
rect 12032 9704 12038 9716
rect 12032 9676 12664 9704
rect 12032 9664 12038 9676
rect 9033 9639 9091 9645
rect 9033 9605 9045 9639
rect 9079 9636 9091 9639
rect 9306 9636 9312 9648
rect 9079 9608 9312 9636
rect 9079 9605 9091 9608
rect 9033 9599 9091 9605
rect 9306 9596 9312 9608
rect 9364 9636 9370 9648
rect 9582 9636 9588 9648
rect 9364 9608 9588 9636
rect 9364 9596 9370 9608
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 10226 9636 10232 9648
rect 9916 9608 10232 9636
rect 9916 9596 9922 9608
rect 10226 9596 10232 9608
rect 10284 9636 10290 9648
rect 10962 9636 10968 9648
rect 10284 9608 10968 9636
rect 10284 9596 10290 9608
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 8849 9571 8907 9577
rect 8849 9537 8861 9571
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 8864 9500 8892 9531
rect 8938 9528 8944 9580
rect 8996 9568 9002 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8996 9540 9137 9568
rect 8996 9528 9002 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 10704 9577 10732 9608
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 12636 9577 12664 9676
rect 14568 9676 15792 9704
rect 13173 9639 13231 9645
rect 13173 9605 13185 9639
rect 13219 9636 13231 9639
rect 14568 9636 14596 9676
rect 15654 9636 15660 9648
rect 13219 9608 14596 9636
rect 14660 9608 15660 9636
rect 13219 9605 13231 9608
rect 13173 9599 13231 9605
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 12621 9571 12679 9577
rect 12621 9537 12633 9571
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 12713 9571 12771 9577
rect 12713 9537 12725 9571
rect 12759 9568 12771 9571
rect 12802 9568 12808 9580
rect 12759 9540 12808 9568
rect 12759 9537 12771 9540
rect 12713 9531 12771 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 12894 9528 12900 9580
rect 12952 9528 12958 9580
rect 14660 9577 14688 9608
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 15764 9636 15792 9676
rect 17310 9636 17316 9648
rect 15764 9608 17316 9636
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 9030 9500 9036 9512
rect 8864 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 12912 9500 12940 9528
rect 12492 9472 12940 9500
rect 12492 9460 12498 9472
rect 9214 9392 9220 9444
rect 9272 9432 9278 9444
rect 9309 9435 9367 9441
rect 9309 9432 9321 9435
rect 9272 9404 9321 9432
rect 9272 9392 9278 9404
rect 9309 9401 9321 9404
rect 9355 9401 9367 9435
rect 13004 9432 13032 9531
rect 14734 9528 14740 9580
rect 14792 9568 14798 9580
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 14792 9540 15209 9568
rect 14792 9528 14798 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 13998 9460 14004 9512
rect 14056 9500 14062 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 14056 9472 14197 9500
rect 14056 9460 14062 9472
rect 14185 9469 14197 9472
rect 14231 9469 14243 9503
rect 14185 9463 14243 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 14384 9432 14412 9463
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 14550 9460 14556 9512
rect 14608 9460 14614 9512
rect 14752 9432 14780 9528
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9500 15347 9503
rect 15470 9500 15476 9512
rect 15335 9472 15476 9500
rect 15335 9469 15347 9472
rect 15289 9463 15347 9469
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 13004 9404 13952 9432
rect 14384 9404 14780 9432
rect 9309 9395 9367 9401
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 10134 9364 10140 9376
rect 7156 9336 10140 9364
rect 7156 9324 7162 9336
rect 10134 9324 10140 9336
rect 10192 9364 10198 9376
rect 10778 9364 10784 9376
rect 10192 9336 10784 9364
rect 10192 9324 10198 9336
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 13924 9364 13952 9404
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 13924 9336 14841 9364
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 2024 9274 17940 9296
rect 2024 9222 3859 9274
rect 3911 9222 3923 9274
rect 3975 9222 3987 9274
rect 4039 9222 4051 9274
rect 4103 9222 4115 9274
rect 4167 9222 7838 9274
rect 7890 9222 7902 9274
rect 7954 9222 7966 9274
rect 8018 9222 8030 9274
rect 8082 9222 8094 9274
rect 8146 9222 11817 9274
rect 11869 9222 11881 9274
rect 11933 9222 11945 9274
rect 11997 9222 12009 9274
rect 12061 9222 12073 9274
rect 12125 9222 15796 9274
rect 15848 9222 15860 9274
rect 15912 9222 15924 9274
rect 15976 9222 15988 9274
rect 16040 9222 16052 9274
rect 16104 9222 17940 9274
rect 2024 9200 17940 9222
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 8202 9160 8208 9172
rect 7423 9132 8208 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8665 9163 8723 9169
rect 8665 9129 8677 9163
rect 8711 9129 8723 9163
rect 8665 9123 8723 9129
rect 8849 9163 8907 9169
rect 8849 9129 8861 9163
rect 8895 9160 8907 9163
rect 8938 9160 8944 9172
rect 8895 9132 8944 9160
rect 8895 9129 8907 9132
rect 8849 9123 8907 9129
rect 7098 9052 7104 9104
rect 7156 9052 7162 9104
rect 7558 9052 7564 9104
rect 7616 9052 7622 9104
rect 8680 9092 8708 9123
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9030 9120 9036 9172
rect 9088 9160 9094 9172
rect 9125 9163 9183 9169
rect 9125 9160 9137 9163
rect 9088 9132 9137 9160
rect 9088 9120 9094 9132
rect 9125 9129 9137 9132
rect 9171 9129 9183 9163
rect 9125 9123 9183 9129
rect 15470 9120 15476 9172
rect 15528 9120 15534 9172
rect 10318 9092 10324 9104
rect 8680 9064 9168 9092
rect 9140 9036 9168 9064
rect 9646 9064 10324 9092
rect 8573 9027 8631 9033
rect 8573 9024 8585 9027
rect 7944 8996 8585 9024
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 6963 8928 7757 8956
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 7745 8925 7757 8928
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 2409 8891 2467 8897
rect 2409 8888 2421 8891
rect 1268 8860 2421 8888
rect 1268 8848 1274 8860
rect 2409 8857 2421 8860
rect 2455 8857 2467 8891
rect 2409 8851 2467 8857
rect 2593 8891 2651 8897
rect 2593 8857 2605 8891
rect 2639 8888 2651 8891
rect 6822 8888 6828 8900
rect 2639 8860 6828 8888
rect 2639 8857 2651 8860
rect 2593 8851 2651 8857
rect 6822 8848 6828 8860
rect 6880 8888 6886 8900
rect 7944 8897 7972 8996
rect 8573 8993 8585 8996
rect 8619 9024 8631 9027
rect 8662 9024 8668 9036
rect 8619 8996 8668 9024
rect 8619 8993 8631 8996
rect 8573 8987 8631 8993
rect 8662 8984 8668 8996
rect 8720 9024 8726 9036
rect 8938 9024 8944 9036
rect 8720 8996 8944 9024
rect 8720 8984 8726 8996
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9122 8984 9128 9036
rect 9180 8984 9186 9036
rect 9646 9024 9674 9064
rect 10318 9052 10324 9064
rect 10376 9052 10382 9104
rect 12250 9024 12256 9036
rect 9416 8996 9674 9024
rect 10244 8996 12256 9024
rect 9416 8968 9444 8996
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 8076 8928 8309 8956
rect 8076 8916 8082 8928
rect 8297 8925 8309 8928
rect 8343 8956 8355 8959
rect 8343 8928 9168 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 7193 8891 7251 8897
rect 7193 8888 7205 8891
rect 6880 8860 7205 8888
rect 6880 8848 6886 8860
rect 7193 8857 7205 8860
rect 7239 8888 7251 8891
rect 7929 8891 7987 8897
rect 7929 8888 7941 8891
rect 7239 8860 7941 8888
rect 7239 8857 7251 8860
rect 7193 8851 7251 8857
rect 7929 8857 7941 8860
rect 7975 8857 7987 8891
rect 7929 8851 7987 8857
rect 8113 8891 8171 8897
rect 8113 8857 8125 8891
rect 8159 8857 8171 8891
rect 8113 8851 8171 8857
rect 7377 8823 7435 8829
rect 7377 8789 7389 8823
rect 7423 8820 7435 8823
rect 7466 8820 7472 8832
rect 7423 8792 7472 8820
rect 7423 8789 7435 8792
rect 7377 8783 7435 8789
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 8128 8820 8156 8851
rect 8938 8848 8944 8900
rect 8996 8897 9002 8900
rect 9140 8897 9168 8928
rect 9398 8916 9404 8968
rect 9456 8916 9462 8968
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10244 8956 10272 8996
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 10244 8928 10333 8956
rect 10137 8919 10195 8925
rect 10321 8925 10333 8928
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 8996 8888 9008 8897
rect 9125 8891 9183 8897
rect 8996 8860 9041 8888
rect 8996 8851 9008 8860
rect 9125 8857 9137 8891
rect 9171 8857 9183 8891
rect 9125 8851 9183 8857
rect 8996 8848 9002 8851
rect 9306 8848 9312 8900
rect 9364 8888 9370 8900
rect 10152 8888 10180 8919
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 13078 8956 13084 8968
rect 10560 8928 13084 8956
rect 10560 8916 10566 8928
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 14458 8916 14464 8968
rect 14516 8956 14522 8968
rect 14734 8956 14740 8968
rect 14516 8928 14740 8956
rect 14516 8916 14522 8928
rect 14734 8916 14740 8928
rect 14792 8956 14798 8968
rect 15013 8959 15071 8965
rect 15013 8956 15025 8959
rect 14792 8928 15025 8956
rect 14792 8916 14798 8928
rect 15013 8925 15025 8928
rect 15059 8925 15071 8959
rect 15013 8919 15071 8925
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15252 8928 15301 8956
rect 15252 8916 15258 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 9364 8860 10180 8888
rect 10413 8891 10471 8897
rect 9364 8848 9370 8860
rect 10413 8857 10425 8891
rect 10459 8888 10471 8891
rect 11698 8888 11704 8900
rect 10459 8860 11704 8888
rect 10459 8857 10471 8860
rect 10413 8851 10471 8857
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 13998 8848 14004 8900
rect 14056 8888 14062 8900
rect 17313 8891 17371 8897
rect 17313 8888 17325 8891
rect 14056 8860 17325 8888
rect 14056 8848 14062 8860
rect 17313 8857 17325 8860
rect 17359 8857 17371 8891
rect 17313 8851 17371 8857
rect 17494 8848 17500 8900
rect 17552 8848 17558 8900
rect 8202 8820 8208 8832
rect 8128 8792 8208 8820
rect 8202 8780 8208 8792
rect 8260 8820 8266 8832
rect 9030 8820 9036 8832
rect 8260 8792 9036 8820
rect 8260 8780 8266 8792
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 10594 8780 10600 8832
rect 10652 8820 10658 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 10652 8792 10701 8820
rect 10652 8780 10658 8792
rect 10689 8789 10701 8792
rect 10735 8789 10747 8823
rect 10689 8783 10747 8789
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 13354 8820 13360 8832
rect 10836 8792 13360 8820
rect 10836 8780 10842 8792
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 14642 8780 14648 8832
rect 14700 8820 14706 8832
rect 15105 8823 15163 8829
rect 15105 8820 15117 8823
rect 14700 8792 15117 8820
rect 14700 8780 14706 8792
rect 15105 8789 15117 8792
rect 15151 8789 15163 8823
rect 15105 8783 15163 8789
rect 2024 8730 17940 8752
rect 2024 8678 4519 8730
rect 4571 8678 4583 8730
rect 4635 8678 4647 8730
rect 4699 8678 4711 8730
rect 4763 8678 4775 8730
rect 4827 8678 8498 8730
rect 8550 8678 8562 8730
rect 8614 8678 8626 8730
rect 8678 8678 8690 8730
rect 8742 8678 8754 8730
rect 8806 8678 12477 8730
rect 12529 8678 12541 8730
rect 12593 8678 12605 8730
rect 12657 8678 12669 8730
rect 12721 8678 12733 8730
rect 12785 8678 16456 8730
rect 16508 8678 16520 8730
rect 16572 8678 16584 8730
rect 16636 8678 16648 8730
rect 16700 8678 16712 8730
rect 16764 8678 17940 8730
rect 2024 8656 17940 8678
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 8018 8616 8024 8628
rect 7340 8588 8024 8616
rect 7340 8576 7346 8588
rect 8018 8576 8024 8588
rect 8076 8616 8082 8628
rect 8205 8619 8263 8625
rect 8205 8616 8217 8619
rect 8076 8588 8217 8616
rect 8076 8576 8082 8588
rect 8205 8585 8217 8588
rect 8251 8585 8263 8619
rect 8205 8579 8263 8585
rect 8849 8619 8907 8625
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 9030 8616 9036 8628
rect 8895 8588 9036 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 12342 8616 12348 8628
rect 9640 8588 12348 8616
rect 9640 8576 9646 8588
rect 7377 8551 7435 8557
rect 7377 8517 7389 8551
rect 7423 8517 7435 8551
rect 7377 8511 7435 8517
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6880 8452 6929 8480
rect 6880 8440 6886 8452
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8480 7067 8483
rect 7392 8480 7420 8511
rect 7558 8508 7564 8560
rect 7616 8508 7622 8560
rect 8386 8508 8392 8560
rect 8444 8508 8450 8560
rect 9398 8508 9404 8560
rect 9456 8508 9462 8560
rect 10594 8548 10600 8560
rect 10428 8520 10600 8548
rect 8404 8480 8432 8508
rect 7055 8452 8432 8480
rect 8757 8483 8815 8489
rect 7055 8449 7067 8452
rect 7009 8443 7067 8449
rect 8757 8449 8769 8483
rect 8803 8480 8815 8483
rect 9122 8480 9128 8492
rect 8803 8452 9128 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 9232 8412 9260 8443
rect 9306 8440 9312 8492
rect 9364 8440 9370 8492
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9631 8452 10057 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 10060 8412 10088 8443
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 10428 8489 10456 8520
rect 10594 8508 10600 8520
rect 10652 8508 10658 8560
rect 11054 8508 11060 8560
rect 11112 8508 11118 8560
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8480 10563 8483
rect 10778 8480 10784 8492
rect 10551 8452 10784 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 10520 8412 10548 8443
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 11072 8480 11100 8508
rect 11256 8489 11284 8588
rect 12342 8576 12348 8588
rect 12400 8616 12406 8628
rect 12618 8616 12624 8628
rect 12400 8588 12624 8616
rect 12400 8576 12406 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12250 8508 12256 8560
rect 12308 8548 12314 8560
rect 12713 8551 12771 8557
rect 12713 8548 12725 8551
rect 12308 8520 12725 8548
rect 12308 8508 12314 8520
rect 12713 8517 12725 8520
rect 12759 8517 12771 8551
rect 12713 8511 12771 8517
rect 12805 8551 12863 8557
rect 12805 8517 12817 8551
rect 12851 8548 12863 8551
rect 13262 8548 13268 8560
rect 12851 8520 13268 8548
rect 12851 8517 12863 8520
rect 12805 8511 12863 8517
rect 13262 8508 13268 8520
rect 13320 8508 13326 8560
rect 11241 8483 11299 8489
rect 11072 8452 11192 8480
rect 10965 8443 11023 8449
rect 8956 8384 9628 8412
rect 10060 8384 10548 8412
rect 7926 8344 7932 8356
rect 7576 8316 7932 8344
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 7576 8285 7604 8316
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8294 8344 8300 8356
rect 8036 8316 8300 8344
rect 7561 8279 7619 8285
rect 7561 8276 7573 8279
rect 7524 8248 7573 8276
rect 7524 8236 7530 8248
rect 7561 8245 7573 8248
rect 7607 8245 7619 8279
rect 7561 8239 7619 8245
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 8036 8285 8064 8316
rect 8294 8304 8300 8316
rect 8352 8344 8358 8356
rect 8956 8344 8984 8384
rect 8352 8316 8984 8344
rect 8352 8304 8358 8316
rect 9030 8304 9036 8356
rect 9088 8304 9094 8356
rect 7745 8279 7803 8285
rect 7745 8276 7757 8279
rect 7708 8248 7757 8276
rect 7708 8236 7714 8248
rect 7745 8245 7757 8248
rect 7791 8245 7803 8279
rect 7745 8239 7803 8245
rect 8021 8279 8079 8285
rect 8021 8245 8033 8279
rect 8067 8245 8079 8279
rect 8021 8239 8079 8245
rect 8202 8236 8208 8288
rect 8260 8236 8266 8288
rect 9600 8276 9628 8384
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 10686 8372 10692 8424
rect 10744 8372 10750 8424
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8412 10931 8415
rect 10980 8412 11008 8443
rect 10919 8384 11008 8412
rect 11057 8415 11115 8421
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 11057 8381 11069 8415
rect 11103 8381 11115 8415
rect 11164 8412 11192 8452
rect 11241 8449 11253 8483
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11532 8412 11560 8443
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12530 8483 12588 8489
rect 12530 8449 12542 8483
rect 12576 8449 12588 8483
rect 12530 8443 12588 8449
rect 12943 8483 13001 8489
rect 12943 8449 12955 8483
rect 12989 8480 13001 8483
rect 13078 8480 13084 8492
rect 12989 8452 13084 8480
rect 12989 8449 13001 8452
rect 12943 8443 13001 8449
rect 11164 8384 11560 8412
rect 11609 8415 11667 8421
rect 11057 8375 11115 8381
rect 11609 8381 11621 8415
rect 11655 8412 11667 8415
rect 12452 8412 12480 8443
rect 11655 8384 12480 8412
rect 11655 8381 11667 8384
rect 11609 8375 11667 8381
rect 10229 8347 10287 8353
rect 10229 8313 10241 8347
rect 10275 8344 10287 8347
rect 11072 8344 11100 8375
rect 10275 8316 11100 8344
rect 10275 8313 10287 8316
rect 10229 8307 10287 8313
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11425 8347 11483 8353
rect 11425 8344 11437 8347
rect 11204 8316 11437 8344
rect 11204 8304 11210 8316
rect 11425 8313 11437 8316
rect 11471 8313 11483 8347
rect 11425 8307 11483 8313
rect 11514 8304 11520 8356
rect 11572 8344 11578 8356
rect 12544 8344 12572 8443
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13633 8483 13691 8489
rect 13219 8452 13584 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13354 8372 13360 8424
rect 13412 8372 13418 8424
rect 13449 8415 13507 8421
rect 13449 8381 13461 8415
rect 13495 8381 13507 8415
rect 13556 8412 13584 8452
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 13814 8480 13820 8492
rect 13679 8452 13820 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14829 8483 14887 8489
rect 14829 8480 14841 8483
rect 14700 8452 14841 8480
rect 14700 8440 14706 8452
rect 14829 8449 14841 8452
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 13556 8384 14473 8412
rect 13449 8375 13507 8381
rect 14461 8381 14473 8384
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 11572 8316 12572 8344
rect 13081 8347 13139 8353
rect 11572 8304 11578 8316
rect 13081 8313 13093 8347
rect 13127 8344 13139 8347
rect 13464 8344 13492 8375
rect 14734 8372 14740 8424
rect 14792 8372 14798 8424
rect 13127 8316 13492 8344
rect 13127 8313 13139 8316
rect 13081 8307 13139 8313
rect 13538 8304 13544 8356
rect 13596 8304 13602 8356
rect 13817 8347 13875 8353
rect 13817 8313 13829 8347
rect 13863 8344 13875 8347
rect 17144 8344 17172 8443
rect 13863 8316 17172 8344
rect 13863 8313 13875 8316
rect 13817 8307 13875 8313
rect 17310 8304 17316 8356
rect 17368 8304 17374 8356
rect 11054 8276 11060 8288
rect 9600 8248 11060 8276
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 11238 8236 11244 8288
rect 11296 8236 11302 8288
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 13170 8276 13176 8288
rect 11388 8248 13176 8276
rect 11388 8236 11394 8248
rect 13170 8236 13176 8248
rect 13228 8276 13234 8288
rect 13630 8276 13636 8288
rect 13228 8248 13636 8276
rect 13228 8236 13234 8248
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 2024 8186 17940 8208
rect 2024 8134 3859 8186
rect 3911 8134 3923 8186
rect 3975 8134 3987 8186
rect 4039 8134 4051 8186
rect 4103 8134 4115 8186
rect 4167 8134 7838 8186
rect 7890 8134 7902 8186
rect 7954 8134 7966 8186
rect 8018 8134 8030 8186
rect 8082 8134 8094 8186
rect 8146 8134 11817 8186
rect 11869 8134 11881 8186
rect 11933 8134 11945 8186
rect 11997 8134 12009 8186
rect 12061 8134 12073 8186
rect 12125 8134 15796 8186
rect 15848 8134 15860 8186
rect 15912 8134 15924 8186
rect 15976 8134 15988 8186
rect 16040 8134 16052 8186
rect 16104 8134 17940 8186
rect 2024 8112 17940 8134
rect 7561 8075 7619 8081
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 9674 8072 9680 8084
rect 7607 8044 9680 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 9674 8032 9680 8044
rect 9732 8072 9738 8084
rect 10226 8072 10232 8084
rect 9732 8044 10232 8072
rect 9732 8032 9738 8044
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 11238 8032 11244 8084
rect 11296 8032 11302 8084
rect 13173 8075 13231 8081
rect 13173 8041 13185 8075
rect 13219 8072 13231 8075
rect 13538 8072 13544 8084
rect 13219 8044 13544 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 13814 8032 13820 8084
rect 13872 8032 13878 8084
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14792 8044 15025 8072
rect 14792 8032 14798 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 11146 8004 11152 8016
rect 10428 7976 11152 8004
rect 10134 7896 10140 7948
rect 10192 7896 10198 7948
rect 10226 7828 10232 7880
rect 10284 7828 10290 7880
rect 10428 7877 10456 7976
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 11333 8007 11391 8013
rect 11333 7973 11345 8007
rect 11379 7973 11391 8007
rect 11333 7967 11391 7973
rect 12253 8007 12311 8013
rect 12253 7973 12265 8007
rect 12299 8004 12311 8007
rect 12299 7976 13492 8004
rect 12299 7973 12311 7976
rect 12253 7967 12311 7973
rect 10594 7896 10600 7948
rect 10652 7936 10658 7948
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 10652 7908 10793 7936
rect 10652 7896 10658 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 11348 7936 11376 7967
rect 10781 7899 10839 7905
rect 10980 7908 11376 7936
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10686 7828 10692 7880
rect 10744 7828 10750 7880
rect 7653 7803 7711 7809
rect 7653 7769 7665 7803
rect 7699 7800 7711 7803
rect 7742 7800 7748 7812
rect 7699 7772 7748 7800
rect 7699 7769 7711 7772
rect 7653 7763 7711 7769
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 10796 7800 10824 7899
rect 10980 7877 11008 7908
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 12713 7939 12771 7945
rect 12713 7936 12725 7939
rect 12676 7908 12725 7936
rect 12676 7896 12682 7908
rect 12713 7905 12725 7908
rect 12759 7905 12771 7939
rect 12713 7899 12771 7905
rect 12802 7896 12808 7948
rect 12860 7896 12866 7948
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7905 12955 7939
rect 12897 7899 12955 7905
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11164 7840 11621 7868
rect 11164 7800 11192 7840
rect 11609 7837 11621 7840
rect 11655 7868 11667 7871
rect 12158 7868 12164 7880
rect 11655 7840 12164 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 12529 7871 12587 7877
rect 12529 7837 12541 7871
rect 12575 7868 12587 7871
rect 12575 7862 12756 7868
rect 12912 7862 12940 7899
rect 12986 7896 12992 7948
rect 13044 7896 13050 7948
rect 13354 7936 13360 7948
rect 13188 7908 13360 7936
rect 13188 7868 13216 7908
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 13004 7862 13216 7868
rect 12575 7840 13216 7862
rect 13265 7871 13323 7877
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 12728 7834 13032 7840
rect 13265 7837 13277 7871
rect 13311 7837 13323 7871
rect 13464 7868 13492 7976
rect 13630 7964 13636 8016
rect 13688 7964 13694 8016
rect 13654 7877 13682 7964
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13464 7840 13553 7868
rect 13265 7831 13323 7837
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 13633 7871 13691 7877
rect 13633 7837 13645 7871
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7868 13967 7871
rect 13998 7868 14004 7880
rect 13955 7840 14004 7868
rect 13955 7837 13967 7840
rect 13909 7831 13967 7837
rect 10796 7772 11192 7800
rect 11330 7760 11336 7812
rect 11388 7800 11394 7812
rect 12253 7803 12311 7809
rect 12253 7800 12265 7803
rect 11388 7772 12265 7800
rect 11388 7760 11394 7772
rect 12253 7769 12265 7772
rect 12299 7769 12311 7803
rect 12253 7763 12311 7769
rect 13280 7800 13308 7831
rect 13924 7800 13952 7831
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 15013 7871 15071 7877
rect 15013 7868 15025 7871
rect 14792 7840 15025 7868
rect 14792 7828 14798 7840
rect 15013 7837 15025 7840
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 15194 7828 15200 7880
rect 15252 7828 15258 7880
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 17586 7828 17592 7880
rect 17644 7828 17650 7880
rect 13280 7772 13952 7800
rect 10597 7735 10655 7741
rect 10597 7701 10609 7735
rect 10643 7732 10655 7735
rect 10686 7732 10692 7744
rect 10643 7704 10692 7732
rect 10643 7701 10655 7704
rect 10597 7695 10655 7701
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 11514 7732 11520 7744
rect 11020 7704 11520 7732
rect 11020 7692 11026 7704
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 12437 7735 12495 7741
rect 12437 7732 12449 7735
rect 11756 7704 12449 7732
rect 11756 7692 11762 7704
rect 12437 7701 12449 7704
rect 12483 7732 12495 7735
rect 12710 7732 12716 7744
rect 12483 7704 12716 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12710 7692 12716 7704
rect 12768 7732 12774 7744
rect 13280 7732 13308 7772
rect 12768 7704 13308 7732
rect 14001 7735 14059 7741
rect 12768 7692 12774 7704
rect 14001 7701 14013 7735
rect 14047 7732 14059 7735
rect 14366 7732 14372 7744
rect 14047 7704 14372 7732
rect 14047 7701 14059 7704
rect 14001 7695 14059 7701
rect 14366 7692 14372 7704
rect 14424 7692 14430 7744
rect 2024 7642 17940 7664
rect 2024 7590 4519 7642
rect 4571 7590 4583 7642
rect 4635 7590 4647 7642
rect 4699 7590 4711 7642
rect 4763 7590 4775 7642
rect 4827 7590 8498 7642
rect 8550 7590 8562 7642
rect 8614 7590 8626 7642
rect 8678 7590 8690 7642
rect 8742 7590 8754 7642
rect 8806 7590 12477 7642
rect 12529 7590 12541 7642
rect 12593 7590 12605 7642
rect 12657 7590 12669 7642
rect 12721 7590 12733 7642
rect 12785 7590 16456 7642
rect 16508 7590 16520 7642
rect 16572 7590 16584 7642
rect 16636 7590 16648 7642
rect 16700 7590 16712 7642
rect 16764 7590 17940 7642
rect 2024 7568 17940 7590
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 11330 7528 11336 7540
rect 7892 7500 11336 7528
rect 7892 7488 7898 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 13357 7531 13415 7537
rect 13357 7497 13369 7531
rect 13403 7528 13415 7531
rect 13906 7528 13912 7540
rect 13403 7500 13912 7528
rect 13403 7497 13415 7500
rect 13357 7491 13415 7497
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 14734 7488 14740 7540
rect 14792 7488 14798 7540
rect 7009 7463 7067 7469
rect 7009 7429 7021 7463
rect 7055 7460 7067 7463
rect 7558 7460 7564 7472
rect 7055 7432 7564 7460
rect 7055 7429 7067 7432
rect 7009 7423 7067 7429
rect 7558 7420 7564 7432
rect 7616 7460 7622 7472
rect 9674 7460 9680 7472
rect 7616 7432 8156 7460
rect 7616 7420 7622 7432
rect 7101 7395 7159 7401
rect 7101 7361 7113 7395
rect 7147 7392 7159 7395
rect 7282 7392 7288 7404
rect 7147 7364 7288 7392
rect 7147 7361 7159 7364
rect 7101 7355 7159 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 8128 7401 8156 7432
rect 8956 7432 9680 7460
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8202 7392 8208 7404
rect 8159 7364 8208 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 8956 7401 8984 7432
rect 9674 7420 9680 7432
rect 9732 7420 9738 7472
rect 14366 7420 14372 7472
rect 14424 7420 14430 7472
rect 14550 7420 14556 7472
rect 14608 7469 14614 7472
rect 14608 7463 14627 7469
rect 14615 7429 14627 7463
rect 15105 7463 15163 7469
rect 15105 7460 15117 7463
rect 14608 7423 14627 7429
rect 14660 7432 15117 7460
rect 14608 7420 14614 7423
rect 8849 7395 8907 7401
rect 8849 7392 8861 7395
rect 8536 7364 8861 7392
rect 8536 7352 8542 7364
rect 8849 7361 8861 7364
rect 8895 7361 8907 7395
rect 8849 7355 8907 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 9306 7392 9312 7404
rect 9171 7364 9312 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 7423 7296 8033 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 8021 7293 8033 7296
rect 8067 7324 8079 7327
rect 8386 7324 8392 7336
rect 8067 7296 8392 7324
rect 8067 7293 8079 7296
rect 8021 7287 8079 7293
rect 8386 7284 8392 7296
rect 8444 7284 8450 7336
rect 8573 7259 8631 7265
rect 7484 7228 7972 7256
rect 7484 7200 7512 7228
rect 7466 7148 7472 7200
rect 7524 7148 7530 7200
rect 7650 7148 7656 7200
rect 7708 7148 7714 7200
rect 7944 7197 7972 7228
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 8662 7256 8668 7268
rect 8619 7228 8668 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 8662 7216 8668 7228
rect 8720 7256 8726 7268
rect 9140 7256 9168 7355
rect 9306 7352 9312 7364
rect 9364 7392 9370 7404
rect 9582 7392 9588 7404
rect 9364 7364 9588 7392
rect 9364 7352 9370 7364
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7392 13047 7395
rect 13354 7392 13360 7404
rect 13035 7364 13360 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 14384 7392 14412 7420
rect 14660 7392 14688 7432
rect 15105 7429 15117 7432
rect 15151 7429 15163 7463
rect 15105 7423 15163 7429
rect 14384 7364 14688 7392
rect 14826 7352 14832 7404
rect 14884 7352 14890 7404
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 13081 7327 13139 7333
rect 13081 7324 13093 7327
rect 12860 7296 13093 7324
rect 12860 7284 12866 7296
rect 13081 7293 13093 7296
rect 13127 7293 13139 7327
rect 14936 7324 14964 7355
rect 13081 7287 13139 7293
rect 14568 7296 14964 7324
rect 8720 7228 9168 7256
rect 8720 7216 8726 7228
rect 7929 7191 7987 7197
rect 7929 7157 7941 7191
rect 7975 7157 7987 7191
rect 7929 7151 7987 7157
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 8352 7160 8401 7188
rect 8352 7148 8358 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 8389 7151 8447 7157
rect 8938 7148 8944 7200
rect 8996 7148 9002 7200
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 12989 7191 13047 7197
rect 12989 7188 13001 7191
rect 12216 7160 13001 7188
rect 12216 7148 12222 7160
rect 12989 7157 13001 7160
rect 13035 7157 13047 7191
rect 12989 7151 13047 7157
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 14568 7197 14596 7296
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7256 15163 7259
rect 15194 7256 15200 7268
rect 15151 7228 15200 7256
rect 15151 7225 15163 7228
rect 15105 7219 15163 7225
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 14553 7191 14611 7197
rect 14553 7188 14565 7191
rect 14148 7160 14565 7188
rect 14148 7148 14154 7160
rect 14553 7157 14565 7160
rect 14599 7157 14611 7191
rect 14553 7151 14611 7157
rect 2024 7098 17940 7120
rect 2024 7046 3859 7098
rect 3911 7046 3923 7098
rect 3975 7046 3987 7098
rect 4039 7046 4051 7098
rect 4103 7046 4115 7098
rect 4167 7046 7838 7098
rect 7890 7046 7902 7098
rect 7954 7046 7966 7098
rect 8018 7046 8030 7098
rect 8082 7046 8094 7098
rect 8146 7046 11817 7098
rect 11869 7046 11881 7098
rect 11933 7046 11945 7098
rect 11997 7046 12009 7098
rect 12061 7046 12073 7098
rect 12125 7046 15796 7098
rect 15848 7046 15860 7098
rect 15912 7046 15924 7098
rect 15976 7046 15988 7098
rect 16040 7046 16052 7098
rect 16104 7046 17940 7098
rect 2024 7024 17940 7046
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 7432 6956 7573 6984
rect 7432 6944 7438 6956
rect 7561 6953 7573 6956
rect 7607 6984 7619 6987
rect 7742 6984 7748 6996
rect 7607 6956 7748 6984
rect 7607 6953 7619 6956
rect 7561 6947 7619 6953
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 8846 6944 8852 6996
rect 8904 6984 8910 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8904 6956 8953 6984
rect 8904 6944 8910 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 11609 6987 11667 6993
rect 11609 6953 11621 6987
rect 11655 6984 11667 6987
rect 12158 6984 12164 6996
rect 11655 6956 12164 6984
rect 11655 6953 11667 6956
rect 11609 6947 11667 6953
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 14090 6944 14096 6996
rect 14148 6944 14154 6996
rect 14461 6987 14519 6993
rect 14461 6953 14473 6987
rect 14507 6984 14519 6987
rect 14550 6984 14556 6996
rect 14507 6956 14556 6984
rect 14507 6953 14519 6956
rect 14461 6947 14519 6953
rect 14550 6944 14556 6956
rect 14608 6984 14614 6996
rect 14826 6984 14832 6996
rect 14608 6956 14832 6984
rect 14608 6944 14614 6956
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 7834 6916 7840 6928
rect 7340 6888 7840 6916
rect 7340 6876 7346 6888
rect 7834 6876 7840 6888
rect 7892 6916 7898 6928
rect 8205 6919 8263 6925
rect 8205 6916 8217 6919
rect 7892 6888 8217 6916
rect 7892 6876 7898 6888
rect 8205 6885 8217 6888
rect 8251 6885 8263 6919
rect 8205 6879 8263 6885
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 12342 6916 12348 6928
rect 8536 6888 9628 6916
rect 8536 6876 8542 6888
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7524 6820 8616 6848
rect 7524 6808 7530 6820
rect 7650 6740 7656 6792
rect 7708 6740 7714 6792
rect 7852 6789 7880 6820
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 8128 6712 8156 6743
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 8588 6789 8616 6820
rect 9030 6808 9036 6860
rect 9088 6808 9094 6860
rect 9600 6848 9628 6888
rect 12084 6888 12348 6916
rect 9600 6820 10272 6848
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 8938 6740 8944 6792
rect 8996 6740 9002 6792
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9217 6743 9275 6749
rect 9416 6752 9689 6780
rect 8662 6712 8668 6724
rect 8128 6684 8668 6712
rect 8662 6672 8668 6684
rect 8720 6672 8726 6724
rect 8849 6715 8907 6721
rect 8849 6681 8861 6715
rect 8895 6712 8907 6715
rect 9232 6712 9260 6743
rect 8895 6684 9260 6712
rect 8895 6681 8907 6684
rect 8849 6675 8907 6681
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6644 7987 6647
rect 8018 6644 8024 6656
rect 7975 6616 8024 6644
rect 7975 6613 7987 6616
rect 7929 6607 7987 6613
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 9416 6653 9444 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 10045 6783 10103 6789
rect 10045 6780 10057 6783
rect 9677 6743 9735 6749
rect 9784 6752 10057 6780
rect 9582 6672 9588 6724
rect 9640 6712 9646 6724
rect 9784 6712 9812 6752
rect 10045 6749 10057 6752
rect 10091 6780 10103 6783
rect 10134 6780 10140 6792
rect 10091 6752 10140 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10244 6789 10272 6820
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 12084 6848 12112 6888
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 11664 6820 12112 6848
rect 11664 6808 11670 6820
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12216 6820 13124 6848
rect 12216 6808 12222 6820
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 10229 6743 10287 6749
rect 11808 6752 12265 6780
rect 9640 6684 9812 6712
rect 9640 6672 9646 6684
rect 9858 6672 9864 6724
rect 9916 6672 9922 6724
rect 10244 6712 10272 6743
rect 11808 6721 11836 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 11793 6715 11851 6721
rect 11793 6712 11805 6715
rect 10244 6684 11805 6712
rect 11793 6681 11805 6684
rect 11839 6681 11851 6715
rect 11793 6675 11851 6681
rect 12066 6672 12072 6724
rect 12124 6672 12130 6724
rect 12268 6712 12296 6743
rect 12342 6740 12348 6792
rect 12400 6740 12406 6792
rect 13096 6789 13124 6820
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 13412 6820 13952 6848
rect 13412 6808 13418 6820
rect 13924 6789 13952 6820
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13633 6783 13691 6789
rect 13633 6780 13645 6783
rect 13495 6752 13645 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13633 6749 13645 6752
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 14461 6783 14519 6789
rect 14461 6780 14473 6783
rect 13955 6752 14473 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 14461 6749 14473 6752
rect 14507 6780 14519 6783
rect 17310 6780 17316 6792
rect 14507 6752 17316 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 12802 6712 12808 6724
rect 12268 6684 12808 6712
rect 12802 6672 12808 6684
rect 12860 6712 12866 6724
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 12860 6684 13277 6712
rect 12860 6672 12866 6684
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13648 6712 13676 6743
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 14185 6715 14243 6721
rect 14185 6712 14197 6715
rect 13648 6684 14197 6712
rect 13265 6675 13323 6681
rect 14185 6681 14197 6684
rect 14231 6681 14243 6715
rect 14185 6675 14243 6681
rect 14369 6715 14427 6721
rect 14369 6681 14381 6715
rect 14415 6681 14427 6715
rect 14369 6675 14427 6681
rect 9401 6647 9459 6653
rect 9401 6613 9413 6647
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 9490 6604 9496 6656
rect 9548 6604 9554 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 11606 6653 11612 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 11204 6616 11437 6644
rect 11204 6604 11210 6616
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 11593 6647 11612 6653
rect 11593 6613 11605 6647
rect 11593 6607 11612 6613
rect 11606 6604 11612 6607
rect 11664 6604 11670 6656
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 12167 6647 12225 6653
rect 12167 6644 12179 6647
rect 12032 6616 12179 6644
rect 12032 6604 12038 6616
rect 12167 6613 12179 6616
rect 12213 6613 12225 6647
rect 12167 6607 12225 6613
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 12400 6616 13737 6644
rect 12400 6604 12406 6616
rect 13725 6613 13737 6616
rect 13771 6644 13783 6647
rect 14384 6644 14412 6675
rect 13771 6616 14412 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 2024 6554 17940 6576
rect 2024 6502 4519 6554
rect 4571 6502 4583 6554
rect 4635 6502 4647 6554
rect 4699 6502 4711 6554
rect 4763 6502 4775 6554
rect 4827 6502 8498 6554
rect 8550 6502 8562 6554
rect 8614 6502 8626 6554
rect 8678 6502 8690 6554
rect 8742 6502 8754 6554
rect 8806 6502 12477 6554
rect 12529 6502 12541 6554
rect 12593 6502 12605 6554
rect 12657 6502 12669 6554
rect 12721 6502 12733 6554
rect 12785 6502 16456 6554
rect 16508 6502 16520 6554
rect 16572 6502 16584 6554
rect 16636 6502 16648 6554
rect 16700 6502 16712 6554
rect 16764 6502 17940 6554
rect 2024 6480 17940 6502
rect 8757 6443 8815 6449
rect 8757 6409 8769 6443
rect 8803 6440 8815 6443
rect 8846 6440 8852 6452
rect 8803 6412 8852 6440
rect 8803 6409 8815 6412
rect 8757 6403 8815 6409
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10284 6412 10425 6440
rect 10284 6400 10290 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 14642 6440 14648 6452
rect 10413 6403 10471 6409
rect 10520 6412 11560 6440
rect 8220 6344 9904 6372
rect 8018 6264 8024 6316
rect 8076 6264 8082 6316
rect 8220 6313 8248 6344
rect 9876 6316 9904 6344
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8536 6276 8585 6304
rect 8536 6264 8542 6276
rect 8573 6273 8585 6276
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 10520 6313 10548 6412
rect 11532 6316 11560 6412
rect 11808 6412 14648 6440
rect 11808 6381 11836 6412
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 11793 6375 11851 6381
rect 11793 6341 11805 6375
rect 11839 6341 11851 6375
rect 11793 6335 11851 6341
rect 11885 6375 11943 6381
rect 11885 6341 11897 6375
rect 11931 6372 11943 6375
rect 12253 6375 12311 6381
rect 12253 6372 12265 6375
rect 11931 6344 12265 6372
rect 11931 6341 11943 6344
rect 11885 6335 11943 6341
rect 12253 6341 12265 6344
rect 12299 6341 12311 6375
rect 12253 6335 12311 6341
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9916 6276 10057 6304
rect 9916 6264 9922 6276
rect 10045 6273 10057 6276
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10735 6276 10793 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6205 8447 6239
rect 8389 6199 8447 6205
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 8404 6168 8432 6199
rect 8260 6140 8432 6168
rect 10060 6168 10088 6267
rect 10962 6264 10968 6316
rect 11020 6264 11026 6316
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 11287 6276 11468 6304
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 11440 6248 11468 6276
rect 11514 6264 11520 6316
rect 11572 6264 11578 6316
rect 11974 6264 11980 6316
rect 12032 6264 12038 6316
rect 10137 6239 10195 6245
rect 10137 6205 10149 6239
rect 10183 6236 10195 6239
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 10183 6208 10609 6236
rect 10183 6205 10195 6208
rect 10137 6199 10195 6205
rect 10597 6205 10609 6208
rect 10643 6205 10655 6239
rect 11333 6239 11391 6245
rect 11333 6228 11345 6239
rect 10597 6199 10655 6205
rect 11164 6205 11345 6228
rect 11379 6205 11391 6239
rect 11164 6200 11391 6205
rect 11164 6168 11192 6200
rect 11333 6199 11391 6200
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 11992 6236 12020 6264
rect 11480 6208 12020 6236
rect 11480 6196 11486 6208
rect 12250 6196 12256 6248
rect 12308 6196 12314 6248
rect 10060 6140 11192 6168
rect 8260 6128 8266 6140
rect 11146 6060 11152 6112
rect 11204 6100 11210 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11204 6072 12081 6100
rect 11204 6060 11210 6072
rect 12069 6069 12081 6072
rect 12115 6069 12127 6103
rect 12069 6063 12127 6069
rect 2024 6010 17940 6032
rect 2024 5958 3859 6010
rect 3911 5958 3923 6010
rect 3975 5958 3987 6010
rect 4039 5958 4051 6010
rect 4103 5958 4115 6010
rect 4167 5958 7838 6010
rect 7890 5958 7902 6010
rect 7954 5958 7966 6010
rect 8018 5958 8030 6010
rect 8082 5958 8094 6010
rect 8146 5958 11817 6010
rect 11869 5958 11881 6010
rect 11933 5958 11945 6010
rect 11997 5958 12009 6010
rect 12061 5958 12073 6010
rect 12125 5958 15796 6010
rect 15848 5958 15860 6010
rect 15912 5958 15924 6010
rect 15976 5958 15988 6010
rect 16040 5958 16052 6010
rect 16104 5958 17940 6010
rect 2024 5936 17940 5958
rect 11514 5856 11520 5908
rect 11572 5856 11578 5908
rect 11422 5788 11428 5840
rect 11480 5788 11486 5840
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 11333 5695 11391 5701
rect 11333 5692 11345 5695
rect 11204 5664 11345 5692
rect 11204 5652 11210 5664
rect 11333 5661 11345 5664
rect 11379 5661 11391 5695
rect 11333 5655 11391 5661
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 11238 5624 11244 5636
rect 11020 5596 11244 5624
rect 11020 5584 11026 5596
rect 11238 5584 11244 5596
rect 11296 5624 11302 5636
rect 11609 5627 11667 5633
rect 11609 5624 11621 5627
rect 11296 5596 11621 5624
rect 11296 5584 11302 5596
rect 11609 5593 11621 5596
rect 11655 5624 11667 5627
rect 12250 5624 12256 5636
rect 11655 5596 12256 5624
rect 11655 5593 11667 5596
rect 11609 5587 11667 5593
rect 12250 5584 12256 5596
rect 12308 5584 12314 5636
rect 2024 5466 17940 5488
rect 2024 5414 4519 5466
rect 4571 5414 4583 5466
rect 4635 5414 4647 5466
rect 4699 5414 4711 5466
rect 4763 5414 4775 5466
rect 4827 5414 8498 5466
rect 8550 5414 8562 5466
rect 8614 5414 8626 5466
rect 8678 5414 8690 5466
rect 8742 5414 8754 5466
rect 8806 5414 12477 5466
rect 12529 5414 12541 5466
rect 12593 5414 12605 5466
rect 12657 5414 12669 5466
rect 12721 5414 12733 5466
rect 12785 5414 16456 5466
rect 16508 5414 16520 5466
rect 16572 5414 16584 5466
rect 16636 5414 16648 5466
rect 16700 5414 16712 5466
rect 16764 5414 17940 5466
rect 2024 5392 17940 5414
rect 2024 4922 17940 4944
rect 2024 4870 3859 4922
rect 3911 4870 3923 4922
rect 3975 4870 3987 4922
rect 4039 4870 4051 4922
rect 4103 4870 4115 4922
rect 4167 4870 7838 4922
rect 7890 4870 7902 4922
rect 7954 4870 7966 4922
rect 8018 4870 8030 4922
rect 8082 4870 8094 4922
rect 8146 4870 11817 4922
rect 11869 4870 11881 4922
rect 11933 4870 11945 4922
rect 11997 4870 12009 4922
rect 12061 4870 12073 4922
rect 12125 4870 15796 4922
rect 15848 4870 15860 4922
rect 15912 4870 15924 4922
rect 15976 4870 15988 4922
rect 16040 4870 16052 4922
rect 16104 4870 17940 4922
rect 2024 4848 17940 4870
rect 2024 4378 17940 4400
rect 2024 4326 4519 4378
rect 4571 4326 4583 4378
rect 4635 4326 4647 4378
rect 4699 4326 4711 4378
rect 4763 4326 4775 4378
rect 4827 4326 8498 4378
rect 8550 4326 8562 4378
rect 8614 4326 8626 4378
rect 8678 4326 8690 4378
rect 8742 4326 8754 4378
rect 8806 4326 12477 4378
rect 12529 4326 12541 4378
rect 12593 4326 12605 4378
rect 12657 4326 12669 4378
rect 12721 4326 12733 4378
rect 12785 4326 16456 4378
rect 16508 4326 16520 4378
rect 16572 4326 16584 4378
rect 16636 4326 16648 4378
rect 16700 4326 16712 4378
rect 16764 4326 17940 4378
rect 2024 4304 17940 4326
rect 2024 3834 17940 3856
rect 2024 3782 3859 3834
rect 3911 3782 3923 3834
rect 3975 3782 3987 3834
rect 4039 3782 4051 3834
rect 4103 3782 4115 3834
rect 4167 3782 7838 3834
rect 7890 3782 7902 3834
rect 7954 3782 7966 3834
rect 8018 3782 8030 3834
rect 8082 3782 8094 3834
rect 8146 3782 11817 3834
rect 11869 3782 11881 3834
rect 11933 3782 11945 3834
rect 11997 3782 12009 3834
rect 12061 3782 12073 3834
rect 12125 3782 15796 3834
rect 15848 3782 15860 3834
rect 15912 3782 15924 3834
rect 15976 3782 15988 3834
rect 16040 3782 16052 3834
rect 16104 3782 17940 3834
rect 2024 3760 17940 3782
rect 2024 3290 17940 3312
rect 2024 3238 4519 3290
rect 4571 3238 4583 3290
rect 4635 3238 4647 3290
rect 4699 3238 4711 3290
rect 4763 3238 4775 3290
rect 4827 3238 8498 3290
rect 8550 3238 8562 3290
rect 8614 3238 8626 3290
rect 8678 3238 8690 3290
rect 8742 3238 8754 3290
rect 8806 3238 12477 3290
rect 12529 3238 12541 3290
rect 12593 3238 12605 3290
rect 12657 3238 12669 3290
rect 12721 3238 12733 3290
rect 12785 3238 16456 3290
rect 16508 3238 16520 3290
rect 16572 3238 16584 3290
rect 16636 3238 16648 3290
rect 16700 3238 16712 3290
rect 16764 3238 17940 3290
rect 2024 3216 17940 3238
rect 10686 3000 10692 3052
rect 10744 3000 10750 3052
rect 10318 2796 10324 2848
rect 10376 2836 10382 2848
rect 10505 2839 10563 2845
rect 10505 2836 10517 2839
rect 10376 2808 10517 2836
rect 10376 2796 10382 2808
rect 10505 2805 10517 2808
rect 10551 2805 10563 2839
rect 10505 2799 10563 2805
rect 2024 2746 17940 2768
rect 2024 2694 3859 2746
rect 3911 2694 3923 2746
rect 3975 2694 3987 2746
rect 4039 2694 4051 2746
rect 4103 2694 4115 2746
rect 4167 2694 7838 2746
rect 7890 2694 7902 2746
rect 7954 2694 7966 2746
rect 8018 2694 8030 2746
rect 8082 2694 8094 2746
rect 8146 2694 11817 2746
rect 11869 2694 11881 2746
rect 11933 2694 11945 2746
rect 11997 2694 12009 2746
rect 12061 2694 12073 2746
rect 12125 2694 15796 2746
rect 15848 2694 15860 2746
rect 15912 2694 15924 2746
rect 15976 2694 15988 2746
rect 16040 2694 16052 2746
rect 16104 2694 17940 2746
rect 2024 2672 17940 2694
rect 8757 2635 8815 2641
rect 8757 2601 8769 2635
rect 8803 2632 8815 2635
rect 9122 2632 9128 2644
rect 8803 2604 9128 2632
rect 8803 2601 8815 2604
rect 8757 2595 8815 2601
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 7742 2524 7748 2576
rect 7800 2564 7806 2576
rect 11977 2567 12035 2573
rect 7800 2536 8156 2564
rect 7800 2524 7806 2536
rect 8128 2505 8156 2536
rect 11977 2533 11989 2567
rect 12023 2564 12035 2567
rect 12158 2564 12164 2576
rect 12023 2536 12164 2564
rect 12023 2533 12035 2536
rect 11977 2527 12035 2533
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2465 8171 2499
rect 8113 2459 8171 2465
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9861 2499 9919 2505
rect 9861 2496 9873 2499
rect 9088 2468 9873 2496
rect 9088 2456 9094 2468
rect 9861 2465 9873 2468
rect 9907 2465 9919 2499
rect 9861 2459 9919 2465
rect 10134 2456 10140 2508
rect 10192 2456 10198 2508
rect 12713 2499 12771 2505
rect 12713 2465 12725 2499
rect 12759 2496 12771 2499
rect 12802 2496 12808 2508
rect 12759 2468 12808 2496
rect 12759 2465 12771 2468
rect 12713 2459 12771 2465
rect 12802 2456 12808 2468
rect 12860 2456 12866 2508
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7800 2400 7849 2428
rect 7800 2388 7806 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8444 2400 8953 2428
rect 8444 2388 8450 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2428 9459 2431
rect 9490 2428 9496 2440
rect 9447 2400 9496 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 11020 2400 11069 2428
rect 11020 2388 11026 2400
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12437 2431 12495 2437
rect 12437 2428 12449 2431
rect 12308 2400 12449 2428
rect 12308 2388 12314 2400
rect 12437 2397 12449 2400
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11664 2332 11805 2360
rect 11664 2320 11670 2332
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 9585 2295 9643 2301
rect 9585 2261 9597 2295
rect 9631 2292 9643 2295
rect 9674 2292 9680 2304
rect 9631 2264 9680 2292
rect 9631 2261 9643 2264
rect 9585 2255 9643 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 2024 2202 17940 2224
rect 2024 2150 4519 2202
rect 4571 2150 4583 2202
rect 4635 2150 4647 2202
rect 4699 2150 4711 2202
rect 4763 2150 4775 2202
rect 4827 2150 8498 2202
rect 8550 2150 8562 2202
rect 8614 2150 8626 2202
rect 8678 2150 8690 2202
rect 8742 2150 8754 2202
rect 8806 2150 12477 2202
rect 12529 2150 12541 2202
rect 12593 2150 12605 2202
rect 12657 2150 12669 2202
rect 12721 2150 12733 2202
rect 12785 2150 16456 2202
rect 16508 2150 16520 2202
rect 16572 2150 16584 2202
rect 16636 2150 16648 2202
rect 16700 2150 16712 2202
rect 16764 2150 17940 2202
rect 2024 2128 17940 2150
<< via1 >>
rect 3859 17926 3911 17978
rect 3923 17926 3975 17978
rect 3987 17926 4039 17978
rect 4051 17926 4103 17978
rect 4115 17926 4167 17978
rect 7838 17926 7890 17978
rect 7902 17926 7954 17978
rect 7966 17926 8018 17978
rect 8030 17926 8082 17978
rect 8094 17926 8146 17978
rect 11817 17926 11869 17978
rect 11881 17926 11933 17978
rect 11945 17926 11997 17978
rect 12009 17926 12061 17978
rect 12073 17926 12125 17978
rect 15796 17926 15848 17978
rect 15860 17926 15912 17978
rect 15924 17926 15976 17978
rect 15988 17926 16040 17978
rect 16052 17926 16104 17978
rect 10324 17824 10376 17876
rect 12256 17824 12308 17876
rect 10600 17756 10652 17808
rect 9036 17620 9088 17672
rect 9680 17620 9732 17672
rect 9404 17595 9456 17604
rect 9404 17561 9413 17595
rect 9413 17561 9447 17595
rect 9447 17561 9456 17595
rect 9404 17552 9456 17561
rect 10968 17620 11020 17672
rect 11612 17620 11664 17672
rect 12808 17620 12860 17672
rect 11428 17552 11480 17604
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 11336 17484 11388 17536
rect 4519 17382 4571 17434
rect 4583 17382 4635 17434
rect 4647 17382 4699 17434
rect 4711 17382 4763 17434
rect 4775 17382 4827 17434
rect 8498 17382 8550 17434
rect 8562 17382 8614 17434
rect 8626 17382 8678 17434
rect 8690 17382 8742 17434
rect 8754 17382 8806 17434
rect 12477 17382 12529 17434
rect 12541 17382 12593 17434
rect 12605 17382 12657 17434
rect 12669 17382 12721 17434
rect 12733 17382 12785 17434
rect 16456 17382 16508 17434
rect 16520 17382 16572 17434
rect 16584 17382 16636 17434
rect 16648 17382 16700 17434
rect 16712 17382 16764 17434
rect 3859 16838 3911 16890
rect 3923 16838 3975 16890
rect 3987 16838 4039 16890
rect 4051 16838 4103 16890
rect 4115 16838 4167 16890
rect 7838 16838 7890 16890
rect 7902 16838 7954 16890
rect 7966 16838 8018 16890
rect 8030 16838 8082 16890
rect 8094 16838 8146 16890
rect 11817 16838 11869 16890
rect 11881 16838 11933 16890
rect 11945 16838 11997 16890
rect 12009 16838 12061 16890
rect 12073 16838 12125 16890
rect 15796 16838 15848 16890
rect 15860 16838 15912 16890
rect 15924 16838 15976 16890
rect 15988 16838 16040 16890
rect 16052 16838 16104 16890
rect 4519 16294 4571 16346
rect 4583 16294 4635 16346
rect 4647 16294 4699 16346
rect 4711 16294 4763 16346
rect 4775 16294 4827 16346
rect 8498 16294 8550 16346
rect 8562 16294 8614 16346
rect 8626 16294 8678 16346
rect 8690 16294 8742 16346
rect 8754 16294 8806 16346
rect 12477 16294 12529 16346
rect 12541 16294 12593 16346
rect 12605 16294 12657 16346
rect 12669 16294 12721 16346
rect 12733 16294 12785 16346
rect 16456 16294 16508 16346
rect 16520 16294 16572 16346
rect 16584 16294 16636 16346
rect 16648 16294 16700 16346
rect 16712 16294 16764 16346
rect 3859 15750 3911 15802
rect 3923 15750 3975 15802
rect 3987 15750 4039 15802
rect 4051 15750 4103 15802
rect 4115 15750 4167 15802
rect 7838 15750 7890 15802
rect 7902 15750 7954 15802
rect 7966 15750 8018 15802
rect 8030 15750 8082 15802
rect 8094 15750 8146 15802
rect 11817 15750 11869 15802
rect 11881 15750 11933 15802
rect 11945 15750 11997 15802
rect 12009 15750 12061 15802
rect 12073 15750 12125 15802
rect 15796 15750 15848 15802
rect 15860 15750 15912 15802
rect 15924 15750 15976 15802
rect 15988 15750 16040 15802
rect 16052 15750 16104 15802
rect 4519 15206 4571 15258
rect 4583 15206 4635 15258
rect 4647 15206 4699 15258
rect 4711 15206 4763 15258
rect 4775 15206 4827 15258
rect 8498 15206 8550 15258
rect 8562 15206 8614 15258
rect 8626 15206 8678 15258
rect 8690 15206 8742 15258
rect 8754 15206 8806 15258
rect 12477 15206 12529 15258
rect 12541 15206 12593 15258
rect 12605 15206 12657 15258
rect 12669 15206 12721 15258
rect 12733 15206 12785 15258
rect 16456 15206 16508 15258
rect 16520 15206 16572 15258
rect 16584 15206 16636 15258
rect 16648 15206 16700 15258
rect 16712 15206 16764 15258
rect 3859 14662 3911 14714
rect 3923 14662 3975 14714
rect 3987 14662 4039 14714
rect 4051 14662 4103 14714
rect 4115 14662 4167 14714
rect 7838 14662 7890 14714
rect 7902 14662 7954 14714
rect 7966 14662 8018 14714
rect 8030 14662 8082 14714
rect 8094 14662 8146 14714
rect 11817 14662 11869 14714
rect 11881 14662 11933 14714
rect 11945 14662 11997 14714
rect 12009 14662 12061 14714
rect 12073 14662 12125 14714
rect 15796 14662 15848 14714
rect 15860 14662 15912 14714
rect 15924 14662 15976 14714
rect 15988 14662 16040 14714
rect 16052 14662 16104 14714
rect 11520 14424 11572 14476
rect 11060 14356 11112 14408
rect 11612 14220 11664 14272
rect 4519 14118 4571 14170
rect 4583 14118 4635 14170
rect 4647 14118 4699 14170
rect 4711 14118 4763 14170
rect 4775 14118 4827 14170
rect 8498 14118 8550 14170
rect 8562 14118 8614 14170
rect 8626 14118 8678 14170
rect 8690 14118 8742 14170
rect 8754 14118 8806 14170
rect 12477 14118 12529 14170
rect 12541 14118 12593 14170
rect 12605 14118 12657 14170
rect 12669 14118 12721 14170
rect 12733 14118 12785 14170
rect 16456 14118 16508 14170
rect 16520 14118 16572 14170
rect 16584 14118 16636 14170
rect 16648 14118 16700 14170
rect 16712 14118 16764 14170
rect 9496 14016 9548 14068
rect 11244 14016 11296 14068
rect 11520 14059 11572 14068
rect 11520 14025 11529 14059
rect 11529 14025 11563 14059
rect 11563 14025 11572 14059
rect 11520 14016 11572 14025
rect 8576 13923 8628 13932
rect 8576 13889 8585 13923
rect 8585 13889 8619 13923
rect 8619 13889 8628 13923
rect 8576 13880 8628 13889
rect 9496 13812 9548 13864
rect 10140 13880 10192 13932
rect 10600 13812 10652 13864
rect 9128 13744 9180 13796
rect 9864 13719 9916 13728
rect 9864 13685 9873 13719
rect 9873 13685 9907 13719
rect 9907 13685 9916 13719
rect 9864 13676 9916 13685
rect 11152 13855 11204 13864
rect 11152 13821 11161 13855
rect 11161 13821 11195 13855
rect 11195 13821 11204 13855
rect 11152 13812 11204 13821
rect 12992 13880 13044 13932
rect 11704 13812 11756 13864
rect 12164 13812 12216 13864
rect 14004 13880 14056 13932
rect 13728 13744 13780 13796
rect 11060 13676 11112 13728
rect 3859 13574 3911 13626
rect 3923 13574 3975 13626
rect 3987 13574 4039 13626
rect 4051 13574 4103 13626
rect 4115 13574 4167 13626
rect 7838 13574 7890 13626
rect 7902 13574 7954 13626
rect 7966 13574 8018 13626
rect 8030 13574 8082 13626
rect 8094 13574 8146 13626
rect 11817 13574 11869 13626
rect 11881 13574 11933 13626
rect 11945 13574 11997 13626
rect 12009 13574 12061 13626
rect 12073 13574 12125 13626
rect 15796 13574 15848 13626
rect 15860 13574 15912 13626
rect 15924 13574 15976 13626
rect 15988 13574 16040 13626
rect 16052 13574 16104 13626
rect 8576 13472 8628 13524
rect 11152 13472 11204 13524
rect 12992 13515 13044 13524
rect 12992 13481 13001 13515
rect 13001 13481 13035 13515
rect 13035 13481 13044 13515
rect 12992 13472 13044 13481
rect 11060 13447 11112 13456
rect 11060 13413 11069 13447
rect 11069 13413 11103 13447
rect 11103 13413 11112 13447
rect 11060 13404 11112 13413
rect 9036 13336 9088 13388
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 9864 13336 9916 13388
rect 8944 13268 8996 13277
rect 6736 13132 6788 13184
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 10140 13268 10192 13320
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 11704 13336 11756 13388
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 13636 13268 13688 13320
rect 13728 13175 13780 13184
rect 13728 13141 13737 13175
rect 13737 13141 13771 13175
rect 13771 13141 13780 13175
rect 13728 13132 13780 13141
rect 4519 13030 4571 13082
rect 4583 13030 4635 13082
rect 4647 13030 4699 13082
rect 4711 13030 4763 13082
rect 4775 13030 4827 13082
rect 8498 13030 8550 13082
rect 8562 13030 8614 13082
rect 8626 13030 8678 13082
rect 8690 13030 8742 13082
rect 8754 13030 8806 13082
rect 12477 13030 12529 13082
rect 12541 13030 12593 13082
rect 12605 13030 12657 13082
rect 12669 13030 12721 13082
rect 12733 13030 12785 13082
rect 16456 13030 16508 13082
rect 16520 13030 16572 13082
rect 16584 13030 16636 13082
rect 16648 13030 16700 13082
rect 16712 13030 16764 13082
rect 8944 12971 8996 12980
rect 8944 12937 8953 12971
rect 8953 12937 8987 12971
rect 8987 12937 8996 12971
rect 8944 12928 8996 12937
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 13360 12928 13412 12980
rect 13636 12971 13688 12980
rect 13636 12937 13645 12971
rect 13645 12937 13679 12971
rect 13679 12937 13688 12971
rect 13636 12928 13688 12937
rect 7380 12860 7432 12912
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 8576 12835 8628 12844
rect 8576 12801 8585 12835
rect 8585 12801 8619 12835
rect 8619 12801 8628 12835
rect 8576 12792 8628 12801
rect 6920 12724 6972 12776
rect 10048 12792 10100 12844
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 16488 12724 16540 12776
rect 7104 12699 7156 12708
rect 7104 12665 7113 12699
rect 7113 12665 7147 12699
rect 7147 12665 7156 12699
rect 7104 12656 7156 12665
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 3859 12486 3911 12538
rect 3923 12486 3975 12538
rect 3987 12486 4039 12538
rect 4051 12486 4103 12538
rect 4115 12486 4167 12538
rect 7838 12486 7890 12538
rect 7902 12486 7954 12538
rect 7966 12486 8018 12538
rect 8030 12486 8082 12538
rect 8094 12486 8146 12538
rect 11817 12486 11869 12538
rect 11881 12486 11933 12538
rect 11945 12486 11997 12538
rect 12009 12486 12061 12538
rect 12073 12486 12125 12538
rect 15796 12486 15848 12538
rect 15860 12486 15912 12538
rect 15924 12486 15976 12538
rect 15988 12486 16040 12538
rect 16052 12486 16104 12538
rect 6920 12427 6972 12436
rect 6920 12393 6929 12427
rect 6929 12393 6963 12427
rect 6963 12393 6972 12427
rect 6920 12384 6972 12393
rect 7104 12384 7156 12436
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 8576 12384 8628 12436
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 12164 12384 12216 12436
rect 12808 12384 12860 12436
rect 7656 12248 7708 12300
rect 9404 12291 9456 12300
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 9404 12248 9456 12257
rect 9956 12248 10008 12300
rect 13820 12248 13872 12300
rect 6368 12180 6420 12232
rect 8208 12180 8260 12232
rect 9220 12180 9272 12232
rect 9312 12223 9364 12232
rect 9312 12189 9321 12223
rect 9321 12189 9355 12223
rect 9355 12189 9364 12223
rect 9312 12180 9364 12189
rect 9036 12112 9088 12164
rect 10692 12180 10744 12232
rect 11336 12180 11388 12232
rect 8208 12044 8260 12096
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 13176 12180 13228 12232
rect 4519 11942 4571 11994
rect 4583 11942 4635 11994
rect 4647 11942 4699 11994
rect 4711 11942 4763 11994
rect 4775 11942 4827 11994
rect 8498 11942 8550 11994
rect 8562 11942 8614 11994
rect 8626 11942 8678 11994
rect 8690 11942 8742 11994
rect 8754 11942 8806 11994
rect 12477 11942 12529 11994
rect 12541 11942 12593 11994
rect 12605 11942 12657 11994
rect 12669 11942 12721 11994
rect 12733 11942 12785 11994
rect 16456 11942 16508 11994
rect 16520 11942 16572 11994
rect 16584 11942 16636 11994
rect 16648 11942 16700 11994
rect 16712 11942 16764 11994
rect 9312 11840 9364 11892
rect 11428 11840 11480 11892
rect 12256 11840 12308 11892
rect 12808 11840 12860 11892
rect 9220 11772 9272 11824
rect 8668 11704 8720 11756
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 11060 11772 11112 11824
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 10324 11704 10376 11756
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 10876 11747 10928 11756
rect 10876 11713 10885 11747
rect 10885 11713 10919 11747
rect 10919 11713 10928 11747
rect 10876 11704 10928 11713
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 1216 11568 1268 11620
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 13268 11772 13320 11824
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 12440 11704 12492 11756
rect 12808 11747 12860 11756
rect 12808 11713 12817 11747
rect 12817 11713 12851 11747
rect 12851 11713 12860 11747
rect 12808 11704 12860 11713
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13084 11747 13136 11756
rect 13084 11713 13093 11747
rect 13093 11713 13127 11747
rect 13127 11713 13136 11747
rect 13084 11704 13136 11713
rect 13176 11704 13228 11756
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 17408 11772 17460 11824
rect 12900 11636 12952 11688
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 17316 11747 17368 11756
rect 17316 11713 17325 11747
rect 17325 11713 17359 11747
rect 17359 11713 17368 11747
rect 17316 11704 17368 11713
rect 13176 11568 13228 11620
rect 13728 11568 13780 11620
rect 14188 11611 14240 11620
rect 14188 11577 14197 11611
rect 14197 11577 14231 11611
rect 14231 11577 14240 11611
rect 14188 11568 14240 11577
rect 14832 11568 14884 11620
rect 3859 11398 3911 11450
rect 3923 11398 3975 11450
rect 3987 11398 4039 11450
rect 4051 11398 4103 11450
rect 4115 11398 4167 11450
rect 7838 11398 7890 11450
rect 7902 11398 7954 11450
rect 7966 11398 8018 11450
rect 8030 11398 8082 11450
rect 8094 11398 8146 11450
rect 11817 11398 11869 11450
rect 11881 11398 11933 11450
rect 11945 11398 11997 11450
rect 12009 11398 12061 11450
rect 12073 11398 12125 11450
rect 15796 11398 15848 11450
rect 15860 11398 15912 11450
rect 15924 11398 15976 11450
rect 15988 11398 16040 11450
rect 16052 11398 16104 11450
rect 7656 11339 7708 11348
rect 7656 11305 7665 11339
rect 7665 11305 7699 11339
rect 7699 11305 7708 11339
rect 7656 11296 7708 11305
rect 8668 11339 8720 11348
rect 8668 11305 8677 11339
rect 8677 11305 8711 11339
rect 8711 11305 8720 11339
rect 8668 11296 8720 11305
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 10876 11296 10928 11348
rect 13452 11296 13504 11348
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 14280 11339 14332 11348
rect 5908 11228 5960 11280
rect 7104 11160 7156 11212
rect 8208 11160 8260 11212
rect 2320 11135 2372 11144
rect 2320 11101 2329 11135
rect 2329 11101 2363 11135
rect 2363 11101 2372 11135
rect 2320 11092 2372 11101
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 6368 11024 6420 11076
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 8852 11135 8904 11144
rect 8852 11101 8861 11135
rect 8861 11101 8895 11135
rect 8895 11101 8904 11135
rect 8852 11092 8904 11101
rect 8944 11135 8996 11144
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 11060 11160 11112 11212
rect 12164 11160 12216 11212
rect 14280 11305 14289 11339
rect 14289 11305 14323 11339
rect 14323 11305 14332 11339
rect 14280 11296 14332 11305
rect 17408 11339 17460 11348
rect 17408 11305 17417 11339
rect 17417 11305 17451 11339
rect 17451 11305 17460 11339
rect 17408 11296 17460 11305
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 12900 11092 12952 11144
rect 14188 11160 14240 11212
rect 14924 11228 14976 11280
rect 13912 11135 13964 11144
rect 13912 11101 13921 11135
rect 13921 11101 13955 11135
rect 13955 11101 13964 11135
rect 13912 11092 13964 11101
rect 9772 11024 9824 11076
rect 13544 11024 13596 11076
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 6644 10956 6696 11008
rect 9864 10956 9916 11008
rect 10324 10956 10376 11008
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 12808 10956 12860 11008
rect 13820 10956 13872 11008
rect 17500 11067 17552 11076
rect 17500 11033 17509 11067
rect 17509 11033 17543 11067
rect 17543 11033 17552 11067
rect 17500 11024 17552 11033
rect 14464 10999 14516 11008
rect 14464 10965 14473 10999
rect 14473 10965 14507 10999
rect 14507 10965 14516 10999
rect 14464 10956 14516 10965
rect 4519 10854 4571 10906
rect 4583 10854 4635 10906
rect 4647 10854 4699 10906
rect 4711 10854 4763 10906
rect 4775 10854 4827 10906
rect 8498 10854 8550 10906
rect 8562 10854 8614 10906
rect 8626 10854 8678 10906
rect 8690 10854 8742 10906
rect 8754 10854 8806 10906
rect 12477 10854 12529 10906
rect 12541 10854 12593 10906
rect 12605 10854 12657 10906
rect 12669 10854 12721 10906
rect 12733 10854 12785 10906
rect 16456 10854 16508 10906
rect 16520 10854 16572 10906
rect 16584 10854 16636 10906
rect 16648 10854 16700 10906
rect 16712 10854 16764 10906
rect 6368 10795 6420 10804
rect 6368 10761 6377 10795
rect 6377 10761 6411 10795
rect 6411 10761 6420 10795
rect 6368 10752 6420 10761
rect 7012 10752 7064 10804
rect 6460 10659 6512 10668
rect 6460 10625 6469 10659
rect 6469 10625 6503 10659
rect 6503 10625 6512 10659
rect 6460 10616 6512 10625
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 7472 10659 7524 10668
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 1124 10548 1176 10600
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 7748 10659 7800 10668
rect 9036 10727 9088 10736
rect 7748 10625 7783 10659
rect 7783 10625 7800 10659
rect 7748 10616 7800 10625
rect 9036 10693 9045 10727
rect 9045 10693 9079 10727
rect 9079 10693 9088 10727
rect 9036 10684 9088 10693
rect 10048 10752 10100 10804
rect 10784 10752 10836 10804
rect 11244 10752 11296 10804
rect 13084 10752 13136 10804
rect 5908 10548 5960 10557
rect 8484 10659 8536 10668
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 8576 10616 8628 10668
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 13728 10684 13780 10736
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 10048 10659 10100 10668
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 10232 10616 10284 10668
rect 10508 10659 10560 10668
rect 10508 10625 10515 10659
rect 10515 10625 10560 10659
rect 10508 10616 10560 10625
rect 11060 10616 11112 10668
rect 11336 10659 11388 10668
rect 11336 10625 11346 10659
rect 11346 10625 11380 10659
rect 11380 10625 11388 10659
rect 11336 10616 11388 10625
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 12624 10616 12676 10668
rect 14464 10616 14516 10668
rect 7656 10412 7708 10464
rect 8484 10412 8536 10464
rect 8576 10412 8628 10464
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 8852 10412 8904 10464
rect 11612 10480 11664 10532
rect 14924 10616 14976 10668
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 14832 10480 14884 10532
rect 15476 10480 15528 10532
rect 12440 10412 12492 10464
rect 12808 10412 12860 10464
rect 15016 10455 15068 10464
rect 15016 10421 15025 10455
rect 15025 10421 15059 10455
rect 15059 10421 15068 10455
rect 15016 10412 15068 10421
rect 15108 10455 15160 10464
rect 15108 10421 15117 10455
rect 15117 10421 15151 10455
rect 15151 10421 15160 10455
rect 15108 10412 15160 10421
rect 3859 10310 3911 10362
rect 3923 10310 3975 10362
rect 3987 10310 4039 10362
rect 4051 10310 4103 10362
rect 4115 10310 4167 10362
rect 7838 10310 7890 10362
rect 7902 10310 7954 10362
rect 7966 10310 8018 10362
rect 8030 10310 8082 10362
rect 8094 10310 8146 10362
rect 11817 10310 11869 10362
rect 11881 10310 11933 10362
rect 11945 10310 11997 10362
rect 12009 10310 12061 10362
rect 12073 10310 12125 10362
rect 15796 10310 15848 10362
rect 15860 10310 15912 10362
rect 15924 10310 15976 10362
rect 15988 10310 16040 10362
rect 16052 10310 16104 10362
rect 5908 10208 5960 10260
rect 7196 10208 7248 10260
rect 8944 10208 8996 10260
rect 10232 10251 10284 10260
rect 10232 10217 10241 10251
rect 10241 10217 10275 10251
rect 10275 10217 10284 10251
rect 10232 10208 10284 10217
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 8484 10140 8536 10192
rect 8392 10072 8444 10124
rect 10508 10140 10560 10192
rect 6460 10004 6512 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 8852 10047 8904 10056
rect 8852 10013 8861 10047
rect 8861 10013 8895 10047
rect 8895 10013 8904 10047
rect 8852 10004 8904 10013
rect 10784 10072 10836 10124
rect 12440 10208 12492 10260
rect 14832 10208 14884 10260
rect 11336 10140 11388 10192
rect 12532 10140 12584 10192
rect 13728 10140 13780 10192
rect 14924 10140 14976 10192
rect 9404 10004 9456 10056
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 10324 9936 10376 9988
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 10968 10004 11020 10056
rect 11612 10072 11664 10124
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 12256 10004 12308 10056
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 12624 9936 12676 9988
rect 7564 9868 7616 9920
rect 7748 9868 7800 9920
rect 8852 9868 8904 9920
rect 10508 9868 10560 9920
rect 10784 9868 10836 9920
rect 12348 9868 12400 9920
rect 12808 9868 12860 9920
rect 13084 9868 13136 9920
rect 13268 9936 13320 9988
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 13820 10047 13872 10056
rect 13820 10013 13829 10047
rect 13829 10013 13863 10047
rect 13863 10013 13872 10047
rect 13820 10004 13872 10013
rect 15108 10072 15160 10124
rect 15016 10047 15068 10056
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 15200 10047 15252 10056
rect 15200 10013 15209 10047
rect 15209 10013 15243 10047
rect 15243 10013 15252 10047
rect 15200 10004 15252 10013
rect 15476 10047 15528 10056
rect 15476 10013 15485 10047
rect 15485 10013 15519 10047
rect 15519 10013 15528 10047
rect 15476 10004 15528 10013
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 14740 9911 14792 9920
rect 14740 9877 14749 9911
rect 14749 9877 14783 9911
rect 14783 9877 14792 9911
rect 14740 9868 14792 9877
rect 15660 9911 15712 9920
rect 15660 9877 15669 9911
rect 15669 9877 15703 9911
rect 15703 9877 15712 9911
rect 15660 9868 15712 9877
rect 17500 9911 17552 9920
rect 17500 9877 17509 9911
rect 17509 9877 17543 9911
rect 17543 9877 17552 9911
rect 17500 9868 17552 9877
rect 4519 9766 4571 9818
rect 4583 9766 4635 9818
rect 4647 9766 4699 9818
rect 4711 9766 4763 9818
rect 4775 9766 4827 9818
rect 8498 9766 8550 9818
rect 8562 9766 8614 9818
rect 8626 9766 8678 9818
rect 8690 9766 8742 9818
rect 8754 9766 8806 9818
rect 12477 9766 12529 9818
rect 12541 9766 12593 9818
rect 12605 9766 12657 9818
rect 12669 9766 12721 9818
rect 12733 9766 12785 9818
rect 16456 9766 16508 9818
rect 16520 9766 16572 9818
rect 16584 9766 16636 9818
rect 16648 9766 16700 9818
rect 16712 9766 16764 9818
rect 10692 9664 10744 9716
rect 11980 9664 12032 9716
rect 9312 9596 9364 9648
rect 9588 9596 9640 9648
rect 9864 9596 9916 9648
rect 10232 9596 10284 9648
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 8944 9528 8996 9580
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 10968 9596 11020 9648
rect 12808 9528 12860 9580
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 15660 9596 15712 9648
rect 17316 9596 17368 9648
rect 9036 9460 9088 9512
rect 12440 9460 12492 9512
rect 9220 9392 9272 9444
rect 14740 9528 14792 9580
rect 14004 9460 14056 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 14556 9503 14608 9512
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 15476 9460 15528 9512
rect 7104 9324 7156 9376
rect 10140 9324 10192 9376
rect 10784 9324 10836 9376
rect 3859 9222 3911 9274
rect 3923 9222 3975 9274
rect 3987 9222 4039 9274
rect 4051 9222 4103 9274
rect 4115 9222 4167 9274
rect 7838 9222 7890 9274
rect 7902 9222 7954 9274
rect 7966 9222 8018 9274
rect 8030 9222 8082 9274
rect 8094 9222 8146 9274
rect 11817 9222 11869 9274
rect 11881 9222 11933 9274
rect 11945 9222 11997 9274
rect 12009 9222 12061 9274
rect 12073 9222 12125 9274
rect 15796 9222 15848 9274
rect 15860 9222 15912 9274
rect 15924 9222 15976 9274
rect 15988 9222 16040 9274
rect 16052 9222 16104 9274
rect 8208 9120 8260 9172
rect 7104 9095 7156 9104
rect 7104 9061 7113 9095
rect 7113 9061 7147 9095
rect 7147 9061 7156 9095
rect 7104 9052 7156 9061
rect 7564 9095 7616 9104
rect 7564 9061 7573 9095
rect 7573 9061 7607 9095
rect 7607 9061 7616 9095
rect 7564 9052 7616 9061
rect 8944 9120 8996 9172
rect 9036 9120 9088 9172
rect 15476 9163 15528 9172
rect 15476 9129 15485 9163
rect 15485 9129 15519 9163
rect 15519 9129 15528 9163
rect 15476 9120 15528 9129
rect 1216 8848 1268 8900
rect 6828 8848 6880 8900
rect 8668 8984 8720 9036
rect 8944 8984 8996 9036
rect 9128 8984 9180 9036
rect 10324 9052 10376 9104
rect 8024 8916 8076 8968
rect 7472 8780 7524 8832
rect 8944 8891 8996 8900
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 12256 8984 12308 9036
rect 8944 8857 8962 8891
rect 8962 8857 8996 8891
rect 8944 8848 8996 8857
rect 9312 8848 9364 8900
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 13084 8916 13136 8968
rect 14464 8916 14516 8968
rect 14740 8916 14792 8968
rect 15200 8916 15252 8968
rect 11704 8848 11756 8900
rect 14004 8848 14056 8900
rect 17500 8891 17552 8900
rect 17500 8857 17509 8891
rect 17509 8857 17543 8891
rect 17543 8857 17552 8891
rect 17500 8848 17552 8857
rect 8208 8780 8260 8832
rect 9036 8780 9088 8832
rect 10600 8780 10652 8832
rect 10784 8780 10836 8832
rect 13360 8780 13412 8832
rect 14648 8780 14700 8832
rect 4519 8678 4571 8730
rect 4583 8678 4635 8730
rect 4647 8678 4699 8730
rect 4711 8678 4763 8730
rect 4775 8678 4827 8730
rect 8498 8678 8550 8730
rect 8562 8678 8614 8730
rect 8626 8678 8678 8730
rect 8690 8678 8742 8730
rect 8754 8678 8806 8730
rect 12477 8678 12529 8730
rect 12541 8678 12593 8730
rect 12605 8678 12657 8730
rect 12669 8678 12721 8730
rect 12733 8678 12785 8730
rect 16456 8678 16508 8730
rect 16520 8678 16572 8730
rect 16584 8678 16636 8730
rect 16648 8678 16700 8730
rect 16712 8678 16764 8730
rect 7288 8576 7340 8628
rect 8024 8576 8076 8628
rect 9036 8576 9088 8628
rect 9588 8576 9640 8628
rect 6828 8440 6880 8492
rect 7564 8551 7616 8560
rect 7564 8517 7573 8551
rect 7573 8517 7607 8551
rect 7607 8517 7616 8551
rect 7564 8508 7616 8517
rect 8392 8551 8444 8560
rect 8392 8517 8401 8551
rect 8401 8517 8435 8551
rect 8435 8517 8444 8551
rect 8392 8508 8444 8517
rect 9404 8551 9456 8560
rect 9404 8517 9413 8551
rect 9413 8517 9447 8551
rect 9447 8517 9456 8551
rect 9404 8508 9456 8517
rect 9128 8440 9180 8492
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 10600 8508 10652 8560
rect 11060 8508 11112 8560
rect 10784 8440 10836 8492
rect 12348 8576 12400 8628
rect 12624 8576 12676 8628
rect 12256 8508 12308 8560
rect 13268 8508 13320 8560
rect 7472 8236 7524 8288
rect 7932 8304 7984 8356
rect 7656 8236 7708 8288
rect 8300 8304 8352 8356
rect 9036 8347 9088 8356
rect 9036 8313 9045 8347
rect 9045 8313 9079 8347
rect 9079 8313 9088 8347
rect 9036 8304 9088 8313
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 8208 8236 8260 8245
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 10692 8415 10744 8424
rect 10692 8381 10701 8415
rect 10701 8381 10735 8415
rect 10735 8381 10744 8415
rect 10692 8372 10744 8381
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 11152 8304 11204 8356
rect 11520 8304 11572 8356
rect 13084 8440 13136 8492
rect 13360 8415 13412 8424
rect 13360 8381 13369 8415
rect 13369 8381 13403 8415
rect 13403 8381 13412 8415
rect 13360 8372 13412 8381
rect 13820 8440 13872 8492
rect 14648 8440 14700 8492
rect 14740 8415 14792 8424
rect 14740 8381 14749 8415
rect 14749 8381 14783 8415
rect 14783 8381 14792 8415
rect 14740 8372 14792 8381
rect 13544 8347 13596 8356
rect 13544 8313 13553 8347
rect 13553 8313 13587 8347
rect 13587 8313 13596 8347
rect 13544 8304 13596 8313
rect 17316 8347 17368 8356
rect 17316 8313 17325 8347
rect 17325 8313 17359 8347
rect 17359 8313 17368 8347
rect 17316 8304 17368 8313
rect 11060 8236 11112 8288
rect 11244 8279 11296 8288
rect 11244 8245 11253 8279
rect 11253 8245 11287 8279
rect 11287 8245 11296 8279
rect 11244 8236 11296 8245
rect 11336 8236 11388 8288
rect 13176 8236 13228 8288
rect 13636 8236 13688 8288
rect 3859 8134 3911 8186
rect 3923 8134 3975 8186
rect 3987 8134 4039 8186
rect 4051 8134 4103 8186
rect 4115 8134 4167 8186
rect 7838 8134 7890 8186
rect 7902 8134 7954 8186
rect 7966 8134 8018 8186
rect 8030 8134 8082 8186
rect 8094 8134 8146 8186
rect 11817 8134 11869 8186
rect 11881 8134 11933 8186
rect 11945 8134 11997 8186
rect 12009 8134 12061 8186
rect 12073 8134 12125 8186
rect 15796 8134 15848 8186
rect 15860 8134 15912 8186
rect 15924 8134 15976 8186
rect 15988 8134 16040 8186
rect 16052 8134 16104 8186
rect 9680 8032 9732 8084
rect 10232 8032 10284 8084
rect 11244 8075 11296 8084
rect 11244 8041 11253 8075
rect 11253 8041 11287 8075
rect 11287 8041 11296 8075
rect 11244 8032 11296 8041
rect 13544 8032 13596 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 14740 8032 14792 8084
rect 10140 7939 10192 7948
rect 10140 7905 10149 7939
rect 10149 7905 10183 7939
rect 10183 7905 10192 7939
rect 10140 7896 10192 7905
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 11152 7964 11204 8016
rect 10600 7896 10652 7948
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 7748 7760 7800 7812
rect 12624 7896 12676 7948
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 12164 7828 12216 7880
rect 12992 7939 13044 7948
rect 12992 7905 13001 7939
rect 13001 7905 13035 7939
rect 13035 7905 13044 7939
rect 12992 7896 13044 7905
rect 13360 7939 13412 7948
rect 13360 7905 13369 7939
rect 13369 7905 13403 7939
rect 13403 7905 13412 7939
rect 13360 7896 13412 7905
rect 13636 7964 13688 8016
rect 11336 7803 11388 7812
rect 11336 7769 11345 7803
rect 11345 7769 11379 7803
rect 11379 7769 11388 7803
rect 11336 7760 11388 7769
rect 14004 7828 14056 7880
rect 14740 7828 14792 7880
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 17316 7828 17368 7837
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 10692 7692 10744 7744
rect 10968 7692 11020 7744
rect 11520 7735 11572 7744
rect 11520 7701 11529 7735
rect 11529 7701 11563 7735
rect 11563 7701 11572 7735
rect 11520 7692 11572 7701
rect 11704 7692 11756 7744
rect 12716 7692 12768 7744
rect 14372 7692 14424 7744
rect 4519 7590 4571 7642
rect 4583 7590 4635 7642
rect 4647 7590 4699 7642
rect 4711 7590 4763 7642
rect 4775 7590 4827 7642
rect 8498 7590 8550 7642
rect 8562 7590 8614 7642
rect 8626 7590 8678 7642
rect 8690 7590 8742 7642
rect 8754 7590 8806 7642
rect 12477 7590 12529 7642
rect 12541 7590 12593 7642
rect 12605 7590 12657 7642
rect 12669 7590 12721 7642
rect 12733 7590 12785 7642
rect 16456 7590 16508 7642
rect 16520 7590 16572 7642
rect 16584 7590 16636 7642
rect 16648 7590 16700 7642
rect 16712 7590 16764 7642
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 7840 7488 7892 7540
rect 11336 7488 11388 7540
rect 13912 7488 13964 7540
rect 14740 7531 14792 7540
rect 14740 7497 14749 7531
rect 14749 7497 14783 7531
rect 14783 7497 14792 7531
rect 14740 7488 14792 7497
rect 7564 7420 7616 7472
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 8208 7352 8260 7404
rect 8484 7352 8536 7404
rect 9680 7420 9732 7472
rect 14372 7463 14424 7472
rect 14372 7429 14381 7463
rect 14381 7429 14415 7463
rect 14415 7429 14424 7463
rect 14372 7420 14424 7429
rect 14556 7463 14608 7472
rect 14556 7429 14581 7463
rect 14581 7429 14608 7463
rect 14556 7420 14608 7429
rect 8392 7284 8444 7336
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 7656 7191 7708 7200
rect 7656 7157 7665 7191
rect 7665 7157 7699 7191
rect 7699 7157 7708 7191
rect 7656 7148 7708 7157
rect 8668 7216 8720 7268
rect 9312 7352 9364 7404
rect 9588 7352 9640 7404
rect 13360 7352 13412 7404
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 12808 7284 12860 7336
rect 8300 7148 8352 7200
rect 8944 7191 8996 7200
rect 8944 7157 8953 7191
rect 8953 7157 8987 7191
rect 8987 7157 8996 7191
rect 8944 7148 8996 7157
rect 12164 7148 12216 7200
rect 14096 7148 14148 7200
rect 15200 7216 15252 7268
rect 3859 7046 3911 7098
rect 3923 7046 3975 7098
rect 3987 7046 4039 7098
rect 4051 7046 4103 7098
rect 4115 7046 4167 7098
rect 7838 7046 7890 7098
rect 7902 7046 7954 7098
rect 7966 7046 8018 7098
rect 8030 7046 8082 7098
rect 8094 7046 8146 7098
rect 11817 7046 11869 7098
rect 11881 7046 11933 7098
rect 11945 7046 11997 7098
rect 12009 7046 12061 7098
rect 12073 7046 12125 7098
rect 15796 7046 15848 7098
rect 15860 7046 15912 7098
rect 15924 7046 15976 7098
rect 15988 7046 16040 7098
rect 16052 7046 16104 7098
rect 7380 6944 7432 6996
rect 7748 6944 7800 6996
rect 8852 6944 8904 6996
rect 12164 6944 12216 6996
rect 14096 6987 14148 6996
rect 14096 6953 14105 6987
rect 14105 6953 14139 6987
rect 14139 6953 14148 6987
rect 14096 6944 14148 6953
rect 14556 6944 14608 6996
rect 14832 6944 14884 6996
rect 7288 6876 7340 6928
rect 7840 6876 7892 6928
rect 8484 6876 8536 6928
rect 7472 6808 7524 6860
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 8484 6783 8536 6792
rect 8484 6749 8493 6783
rect 8493 6749 8527 6783
rect 8527 6749 8536 6783
rect 8484 6740 8536 6749
rect 9036 6851 9088 6860
rect 9036 6817 9045 6851
rect 9045 6817 9079 6851
rect 9079 6817 9088 6851
rect 9036 6808 9088 6817
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 8668 6672 8720 6724
rect 8024 6604 8076 6656
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 9588 6672 9640 6724
rect 10140 6740 10192 6792
rect 11612 6808 11664 6860
rect 12348 6876 12400 6928
rect 12164 6808 12216 6860
rect 9864 6715 9916 6724
rect 9864 6681 9873 6715
rect 9873 6681 9907 6715
rect 9907 6681 9916 6715
rect 9864 6672 9916 6681
rect 12072 6715 12124 6724
rect 12072 6681 12081 6715
rect 12081 6681 12115 6715
rect 12115 6681 12124 6715
rect 12072 6672 12124 6681
rect 12348 6783 12400 6792
rect 12348 6749 12357 6783
rect 12357 6749 12391 6783
rect 12391 6749 12400 6783
rect 12348 6740 12400 6749
rect 13360 6808 13412 6860
rect 12808 6672 12860 6724
rect 17316 6740 17368 6792
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 11152 6604 11204 6656
rect 11612 6647 11664 6656
rect 11612 6613 11639 6647
rect 11639 6613 11664 6647
rect 11612 6604 11664 6613
rect 11980 6604 12032 6656
rect 12348 6604 12400 6656
rect 4519 6502 4571 6554
rect 4583 6502 4635 6554
rect 4647 6502 4699 6554
rect 4711 6502 4763 6554
rect 4775 6502 4827 6554
rect 8498 6502 8550 6554
rect 8562 6502 8614 6554
rect 8626 6502 8678 6554
rect 8690 6502 8742 6554
rect 8754 6502 8806 6554
rect 12477 6502 12529 6554
rect 12541 6502 12593 6554
rect 12605 6502 12657 6554
rect 12669 6502 12721 6554
rect 12733 6502 12785 6554
rect 16456 6502 16508 6554
rect 16520 6502 16572 6554
rect 16584 6502 16636 6554
rect 16648 6502 16700 6554
rect 16712 6502 16764 6554
rect 8852 6400 8904 6452
rect 10232 6400 10284 6452
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8484 6264 8536 6316
rect 9864 6264 9916 6316
rect 14648 6400 14700 6452
rect 8208 6128 8260 6180
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 11520 6307 11572 6316
rect 11520 6273 11529 6307
rect 11529 6273 11563 6307
rect 11563 6273 11572 6307
rect 11520 6264 11572 6273
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 11428 6196 11480 6248
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 11152 6060 11204 6112
rect 3859 5958 3911 6010
rect 3923 5958 3975 6010
rect 3987 5958 4039 6010
rect 4051 5958 4103 6010
rect 4115 5958 4167 6010
rect 7838 5958 7890 6010
rect 7902 5958 7954 6010
rect 7966 5958 8018 6010
rect 8030 5958 8082 6010
rect 8094 5958 8146 6010
rect 11817 5958 11869 6010
rect 11881 5958 11933 6010
rect 11945 5958 11997 6010
rect 12009 5958 12061 6010
rect 12073 5958 12125 6010
rect 15796 5958 15848 6010
rect 15860 5958 15912 6010
rect 15924 5958 15976 6010
rect 15988 5958 16040 6010
rect 16052 5958 16104 6010
rect 11520 5899 11572 5908
rect 11520 5865 11529 5899
rect 11529 5865 11563 5899
rect 11563 5865 11572 5899
rect 11520 5856 11572 5865
rect 11428 5831 11480 5840
rect 11428 5797 11437 5831
rect 11437 5797 11471 5831
rect 11471 5797 11480 5831
rect 11428 5788 11480 5797
rect 11152 5652 11204 5704
rect 10968 5584 11020 5636
rect 11244 5584 11296 5636
rect 12256 5584 12308 5636
rect 4519 5414 4571 5466
rect 4583 5414 4635 5466
rect 4647 5414 4699 5466
rect 4711 5414 4763 5466
rect 4775 5414 4827 5466
rect 8498 5414 8550 5466
rect 8562 5414 8614 5466
rect 8626 5414 8678 5466
rect 8690 5414 8742 5466
rect 8754 5414 8806 5466
rect 12477 5414 12529 5466
rect 12541 5414 12593 5466
rect 12605 5414 12657 5466
rect 12669 5414 12721 5466
rect 12733 5414 12785 5466
rect 16456 5414 16508 5466
rect 16520 5414 16572 5466
rect 16584 5414 16636 5466
rect 16648 5414 16700 5466
rect 16712 5414 16764 5466
rect 3859 4870 3911 4922
rect 3923 4870 3975 4922
rect 3987 4870 4039 4922
rect 4051 4870 4103 4922
rect 4115 4870 4167 4922
rect 7838 4870 7890 4922
rect 7902 4870 7954 4922
rect 7966 4870 8018 4922
rect 8030 4870 8082 4922
rect 8094 4870 8146 4922
rect 11817 4870 11869 4922
rect 11881 4870 11933 4922
rect 11945 4870 11997 4922
rect 12009 4870 12061 4922
rect 12073 4870 12125 4922
rect 15796 4870 15848 4922
rect 15860 4870 15912 4922
rect 15924 4870 15976 4922
rect 15988 4870 16040 4922
rect 16052 4870 16104 4922
rect 4519 4326 4571 4378
rect 4583 4326 4635 4378
rect 4647 4326 4699 4378
rect 4711 4326 4763 4378
rect 4775 4326 4827 4378
rect 8498 4326 8550 4378
rect 8562 4326 8614 4378
rect 8626 4326 8678 4378
rect 8690 4326 8742 4378
rect 8754 4326 8806 4378
rect 12477 4326 12529 4378
rect 12541 4326 12593 4378
rect 12605 4326 12657 4378
rect 12669 4326 12721 4378
rect 12733 4326 12785 4378
rect 16456 4326 16508 4378
rect 16520 4326 16572 4378
rect 16584 4326 16636 4378
rect 16648 4326 16700 4378
rect 16712 4326 16764 4378
rect 3859 3782 3911 3834
rect 3923 3782 3975 3834
rect 3987 3782 4039 3834
rect 4051 3782 4103 3834
rect 4115 3782 4167 3834
rect 7838 3782 7890 3834
rect 7902 3782 7954 3834
rect 7966 3782 8018 3834
rect 8030 3782 8082 3834
rect 8094 3782 8146 3834
rect 11817 3782 11869 3834
rect 11881 3782 11933 3834
rect 11945 3782 11997 3834
rect 12009 3782 12061 3834
rect 12073 3782 12125 3834
rect 15796 3782 15848 3834
rect 15860 3782 15912 3834
rect 15924 3782 15976 3834
rect 15988 3782 16040 3834
rect 16052 3782 16104 3834
rect 4519 3238 4571 3290
rect 4583 3238 4635 3290
rect 4647 3238 4699 3290
rect 4711 3238 4763 3290
rect 4775 3238 4827 3290
rect 8498 3238 8550 3290
rect 8562 3238 8614 3290
rect 8626 3238 8678 3290
rect 8690 3238 8742 3290
rect 8754 3238 8806 3290
rect 12477 3238 12529 3290
rect 12541 3238 12593 3290
rect 12605 3238 12657 3290
rect 12669 3238 12721 3290
rect 12733 3238 12785 3290
rect 16456 3238 16508 3290
rect 16520 3238 16572 3290
rect 16584 3238 16636 3290
rect 16648 3238 16700 3290
rect 16712 3238 16764 3290
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 10324 2796 10376 2848
rect 3859 2694 3911 2746
rect 3923 2694 3975 2746
rect 3987 2694 4039 2746
rect 4051 2694 4103 2746
rect 4115 2694 4167 2746
rect 7838 2694 7890 2746
rect 7902 2694 7954 2746
rect 7966 2694 8018 2746
rect 8030 2694 8082 2746
rect 8094 2694 8146 2746
rect 11817 2694 11869 2746
rect 11881 2694 11933 2746
rect 11945 2694 11997 2746
rect 12009 2694 12061 2746
rect 12073 2694 12125 2746
rect 15796 2694 15848 2746
rect 15860 2694 15912 2746
rect 15924 2694 15976 2746
rect 15988 2694 16040 2746
rect 16052 2694 16104 2746
rect 9128 2592 9180 2644
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 7748 2524 7800 2576
rect 12164 2524 12216 2576
rect 9036 2456 9088 2508
rect 10140 2499 10192 2508
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 12808 2456 12860 2508
rect 7748 2388 7800 2440
rect 8392 2388 8444 2440
rect 9496 2388 9548 2440
rect 10968 2388 11020 2440
rect 12256 2388 12308 2440
rect 11612 2320 11664 2372
rect 9680 2252 9732 2304
rect 4519 2150 4571 2202
rect 4583 2150 4635 2202
rect 4647 2150 4699 2202
rect 4711 2150 4763 2202
rect 4775 2150 4827 2202
rect 8498 2150 8550 2202
rect 8562 2150 8614 2202
rect 8626 2150 8678 2202
rect 8690 2150 8742 2202
rect 8754 2150 8806 2202
rect 12477 2150 12529 2202
rect 12541 2150 12593 2202
rect 12605 2150 12657 2202
rect 12669 2150 12721 2202
rect 12733 2150 12785 2202
rect 16456 2150 16508 2202
rect 16520 2150 16572 2202
rect 16584 2150 16636 2202
rect 16648 2150 16700 2202
rect 16712 2150 16764 2202
<< metal2 >>
rect 9034 19200 9090 20000
rect 9678 19200 9734 20000
rect 10322 19200 10378 20000
rect 10966 19200 11022 20000
rect 11610 19200 11666 20000
rect 12254 19200 12310 20000
rect 3859 17980 4167 17989
rect 3859 17978 3865 17980
rect 3921 17978 3945 17980
rect 4001 17978 4025 17980
rect 4081 17978 4105 17980
rect 4161 17978 4167 17980
rect 3921 17926 3923 17978
rect 4103 17926 4105 17978
rect 3859 17924 3865 17926
rect 3921 17924 3945 17926
rect 4001 17924 4025 17926
rect 4081 17924 4105 17926
rect 4161 17924 4167 17926
rect 3859 17915 4167 17924
rect 7838 17980 8146 17989
rect 7838 17978 7844 17980
rect 7900 17978 7924 17980
rect 7980 17978 8004 17980
rect 8060 17978 8084 17980
rect 8140 17978 8146 17980
rect 7900 17926 7902 17978
rect 8082 17926 8084 17978
rect 7838 17924 7844 17926
rect 7900 17924 7924 17926
rect 7980 17924 8004 17926
rect 8060 17924 8084 17926
rect 8140 17924 8146 17926
rect 7838 17915 8146 17924
rect 9048 17678 9076 19200
rect 9692 17678 9720 19200
rect 10336 17882 10364 19200
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 4519 17436 4827 17445
rect 4519 17434 4525 17436
rect 4581 17434 4605 17436
rect 4661 17434 4685 17436
rect 4741 17434 4765 17436
rect 4821 17434 4827 17436
rect 4581 17382 4583 17434
rect 4763 17382 4765 17434
rect 4519 17380 4525 17382
rect 4581 17380 4605 17382
rect 4661 17380 4685 17382
rect 4741 17380 4765 17382
rect 4821 17380 4827 17382
rect 4519 17371 4827 17380
rect 8498 17436 8806 17445
rect 8498 17434 8504 17436
rect 8560 17434 8584 17436
rect 8640 17434 8664 17436
rect 8720 17434 8744 17436
rect 8800 17434 8806 17436
rect 8560 17382 8562 17434
rect 8742 17382 8744 17434
rect 8498 17380 8504 17382
rect 8560 17380 8584 17382
rect 8640 17380 8664 17382
rect 8720 17380 8744 17382
rect 8800 17380 8806 17382
rect 8498 17371 8806 17380
rect 3859 16892 4167 16901
rect 3859 16890 3865 16892
rect 3921 16890 3945 16892
rect 4001 16890 4025 16892
rect 4081 16890 4105 16892
rect 4161 16890 4167 16892
rect 3921 16838 3923 16890
rect 4103 16838 4105 16890
rect 3859 16836 3865 16838
rect 3921 16836 3945 16838
rect 4001 16836 4025 16838
rect 4081 16836 4105 16838
rect 4161 16836 4167 16838
rect 3859 16827 4167 16836
rect 7838 16892 8146 16901
rect 7838 16890 7844 16892
rect 7900 16890 7924 16892
rect 7980 16890 8004 16892
rect 8060 16890 8084 16892
rect 8140 16890 8146 16892
rect 7900 16838 7902 16890
rect 8082 16838 8084 16890
rect 7838 16836 7844 16838
rect 7900 16836 7924 16838
rect 7980 16836 8004 16838
rect 8060 16836 8084 16838
rect 8140 16836 8146 16838
rect 7838 16827 8146 16836
rect 4519 16348 4827 16357
rect 4519 16346 4525 16348
rect 4581 16346 4605 16348
rect 4661 16346 4685 16348
rect 4741 16346 4765 16348
rect 4821 16346 4827 16348
rect 4581 16294 4583 16346
rect 4763 16294 4765 16346
rect 4519 16292 4525 16294
rect 4581 16292 4605 16294
rect 4661 16292 4685 16294
rect 4741 16292 4765 16294
rect 4821 16292 4827 16294
rect 4519 16283 4827 16292
rect 8498 16348 8806 16357
rect 8498 16346 8504 16348
rect 8560 16346 8584 16348
rect 8640 16346 8664 16348
rect 8720 16346 8744 16348
rect 8800 16346 8806 16348
rect 8560 16294 8562 16346
rect 8742 16294 8744 16346
rect 8498 16292 8504 16294
rect 8560 16292 8584 16294
rect 8640 16292 8664 16294
rect 8720 16292 8744 16294
rect 8800 16292 8806 16294
rect 8498 16283 8806 16292
rect 3859 15804 4167 15813
rect 3859 15802 3865 15804
rect 3921 15802 3945 15804
rect 4001 15802 4025 15804
rect 4081 15802 4105 15804
rect 4161 15802 4167 15804
rect 3921 15750 3923 15802
rect 4103 15750 4105 15802
rect 3859 15748 3865 15750
rect 3921 15748 3945 15750
rect 4001 15748 4025 15750
rect 4081 15748 4105 15750
rect 4161 15748 4167 15750
rect 3859 15739 4167 15748
rect 7838 15804 8146 15813
rect 7838 15802 7844 15804
rect 7900 15802 7924 15804
rect 7980 15802 8004 15804
rect 8060 15802 8084 15804
rect 8140 15802 8146 15804
rect 7900 15750 7902 15802
rect 8082 15750 8084 15802
rect 7838 15748 7844 15750
rect 7900 15748 7924 15750
rect 7980 15748 8004 15750
rect 8060 15748 8084 15750
rect 8140 15748 8146 15750
rect 7838 15739 8146 15748
rect 4519 15260 4827 15269
rect 4519 15258 4525 15260
rect 4581 15258 4605 15260
rect 4661 15258 4685 15260
rect 4741 15258 4765 15260
rect 4821 15258 4827 15260
rect 4581 15206 4583 15258
rect 4763 15206 4765 15258
rect 4519 15204 4525 15206
rect 4581 15204 4605 15206
rect 4661 15204 4685 15206
rect 4741 15204 4765 15206
rect 4821 15204 4827 15206
rect 4519 15195 4827 15204
rect 8498 15260 8806 15269
rect 8498 15258 8504 15260
rect 8560 15258 8584 15260
rect 8640 15258 8664 15260
rect 8720 15258 8744 15260
rect 8800 15258 8806 15260
rect 8560 15206 8562 15258
rect 8742 15206 8744 15258
rect 8498 15204 8504 15206
rect 8560 15204 8584 15206
rect 8640 15204 8664 15206
rect 8720 15204 8744 15206
rect 8800 15204 8806 15206
rect 8498 15195 8806 15204
rect 3859 14716 4167 14725
rect 3859 14714 3865 14716
rect 3921 14714 3945 14716
rect 4001 14714 4025 14716
rect 4081 14714 4105 14716
rect 4161 14714 4167 14716
rect 3921 14662 3923 14714
rect 4103 14662 4105 14714
rect 3859 14660 3865 14662
rect 3921 14660 3945 14662
rect 4001 14660 4025 14662
rect 4081 14660 4105 14662
rect 4161 14660 4167 14662
rect 3859 14651 4167 14660
rect 7838 14716 8146 14725
rect 7838 14714 7844 14716
rect 7900 14714 7924 14716
rect 7980 14714 8004 14716
rect 8060 14714 8084 14716
rect 8140 14714 8146 14716
rect 7900 14662 7902 14714
rect 8082 14662 8084 14714
rect 7838 14660 7844 14662
rect 7900 14660 7924 14662
rect 7980 14660 8004 14662
rect 8060 14660 8084 14662
rect 8140 14660 8146 14662
rect 7838 14651 8146 14660
rect 4519 14172 4827 14181
rect 4519 14170 4525 14172
rect 4581 14170 4605 14172
rect 4661 14170 4685 14172
rect 4741 14170 4765 14172
rect 4821 14170 4827 14172
rect 4581 14118 4583 14170
rect 4763 14118 4765 14170
rect 4519 14116 4525 14118
rect 4581 14116 4605 14118
rect 4661 14116 4685 14118
rect 4741 14116 4765 14118
rect 4821 14116 4827 14118
rect 4519 14107 4827 14116
rect 8498 14172 8806 14181
rect 8498 14170 8504 14172
rect 8560 14170 8584 14172
rect 8640 14170 8664 14172
rect 8720 14170 8744 14172
rect 8800 14170 8806 14172
rect 8560 14118 8562 14170
rect 8742 14118 8744 14170
rect 8498 14116 8504 14118
rect 8560 14116 8584 14118
rect 8640 14116 8664 14118
rect 8720 14116 8744 14118
rect 8800 14116 8806 14118
rect 8498 14107 8806 14116
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 3859 13628 4167 13637
rect 3859 13626 3865 13628
rect 3921 13626 3945 13628
rect 4001 13626 4025 13628
rect 4081 13626 4105 13628
rect 4161 13626 4167 13628
rect 3921 13574 3923 13626
rect 4103 13574 4105 13626
rect 3859 13572 3865 13574
rect 3921 13572 3945 13574
rect 4001 13572 4025 13574
rect 4081 13572 4105 13574
rect 4161 13572 4167 13574
rect 3859 13563 4167 13572
rect 7838 13628 8146 13637
rect 7838 13626 7844 13628
rect 7900 13626 7924 13628
rect 7980 13626 8004 13628
rect 8060 13626 8084 13628
rect 8140 13626 8146 13628
rect 7900 13574 7902 13626
rect 8082 13574 8084 13626
rect 7838 13572 7844 13574
rect 7900 13572 7924 13574
rect 7980 13572 8004 13574
rect 8060 13572 8084 13574
rect 8140 13572 8146 13574
rect 7838 13563 8146 13572
rect 8588 13530 8616 13874
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 4519 13084 4827 13093
rect 4519 13082 4525 13084
rect 4581 13082 4605 13084
rect 4661 13082 4685 13084
rect 4741 13082 4765 13084
rect 4821 13082 4827 13084
rect 4581 13030 4583 13082
rect 4763 13030 4765 13082
rect 4519 13028 4525 13030
rect 4581 13028 4605 13030
rect 4661 13028 4685 13030
rect 4741 13028 4765 13030
rect 4821 13028 4827 13030
rect 4519 13019 4827 13028
rect 6748 12850 6776 13126
rect 8498 13084 8806 13093
rect 8498 13082 8504 13084
rect 8560 13082 8584 13084
rect 8640 13082 8664 13084
rect 8720 13082 8744 13084
rect 8800 13082 8806 13084
rect 8560 13030 8562 13082
rect 8742 13030 8744 13082
rect 8498 13028 8504 13030
rect 8560 13028 8584 13030
rect 8640 13028 8664 13030
rect 8720 13028 8744 13030
rect 8800 13028 8806 13030
rect 8498 13019 8806 13028
rect 8956 12986 8984 13262
rect 9048 12986 9076 13330
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 12345 2452 12582
rect 3859 12540 4167 12549
rect 3859 12538 3865 12540
rect 3921 12538 3945 12540
rect 4001 12538 4025 12540
rect 4081 12538 4105 12540
rect 4161 12538 4167 12540
rect 3921 12486 3923 12538
rect 4103 12486 4105 12538
rect 3859 12484 3865 12486
rect 3921 12484 3945 12486
rect 4001 12484 4025 12486
rect 4081 12484 4105 12486
rect 4161 12484 4167 12486
rect 3859 12475 4167 12484
rect 6932 12442 6960 12718
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7116 12442 7144 12650
rect 7392 12442 7420 12854
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 7838 12540 8146 12549
rect 7838 12538 7844 12540
rect 7900 12538 7924 12540
rect 7980 12538 8004 12540
rect 8060 12538 8084 12540
rect 8140 12538 8146 12540
rect 7900 12486 7902 12538
rect 8082 12486 8084 12538
rect 7838 12484 7844 12486
rect 7900 12484 7924 12486
rect 7980 12484 8004 12486
rect 8060 12484 8084 12486
rect 8140 12484 8146 12486
rect 7838 12475 8146 12484
rect 8588 12442 8616 12786
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 2410 12336 2466 12345
rect 2410 12271 2466 12280
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 4519 11996 4827 12005
rect 4519 11994 4525 11996
rect 4581 11994 4605 11996
rect 4661 11994 4685 11996
rect 4741 11994 4765 11996
rect 4821 11994 4827 11996
rect 4581 11942 4583 11994
rect 4763 11942 4765 11994
rect 4519 11940 4525 11942
rect 4581 11940 4605 11942
rect 4661 11940 4685 11942
rect 4741 11940 4765 11942
rect 4821 11940 4827 11942
rect 4519 11931 4827 11940
rect 1214 11656 1270 11665
rect 1214 11591 1216 11600
rect 1268 11591 1270 11600
rect 1216 11562 1268 11568
rect 3859 11452 4167 11461
rect 3859 11450 3865 11452
rect 3921 11450 3945 11452
rect 4001 11450 4025 11452
rect 4081 11450 4105 11452
rect 4161 11450 4167 11452
rect 3921 11398 3923 11450
rect 4103 11398 4105 11450
rect 3859 11396 3865 11398
rect 3921 11396 3945 11398
rect 4001 11396 4025 11398
rect 4081 11396 4105 11398
rect 4161 11396 4167 11398
rect 3859 11387 4167 11396
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2332 10985 2360 11086
rect 2318 10976 2374 10985
rect 2318 10911 2374 10920
rect 4519 10908 4827 10917
rect 4519 10906 4525 10908
rect 4581 10906 4605 10908
rect 4661 10906 4685 10908
rect 4741 10906 4765 10908
rect 4821 10906 4827 10908
rect 4581 10854 4583 10906
rect 4763 10854 4765 10906
rect 4519 10852 4525 10854
rect 4581 10852 4605 10854
rect 4661 10852 4685 10854
rect 4741 10852 4765 10854
rect 4821 10852 4827 10854
rect 4519 10843 4827 10852
rect 5920 10606 5948 11222
rect 6380 11082 6408 12174
rect 7668 11354 7696 12242
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 12102 8248 12174
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 7838 11452 8146 11461
rect 7838 11450 7844 11452
rect 7900 11450 7924 11452
rect 7980 11450 8004 11452
rect 8060 11450 8084 11452
rect 8140 11450 8146 11452
rect 7900 11398 7902 11450
rect 8082 11398 8084 11450
rect 7838 11396 7844 11398
rect 7900 11396 7924 11398
rect 7980 11396 8004 11398
rect 8060 11396 8084 11398
rect 8140 11396 8146 11398
rect 7838 11387 8146 11396
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 8220 11218 8248 12038
rect 8498 11996 8806 12005
rect 8498 11994 8504 11996
rect 8560 11994 8584 11996
rect 8640 11994 8664 11996
rect 8720 11994 8744 11996
rect 8800 11994 8806 11996
rect 8560 11942 8562 11994
rect 8742 11942 8744 11994
rect 8498 11940 8504 11942
rect 8560 11940 8584 11942
rect 8640 11940 8664 11942
rect 8720 11940 8744 11942
rect 8800 11940 8806 11942
rect 8498 11931 8806 11940
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8680 11354 8708 11698
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6380 10810 6408 11018
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6656 10674 6684 10950
rect 7024 10810 7052 11086
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 1124 10600 1176 10606
rect 1124 10542 1176 10548
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 1136 10305 1164 10542
rect 3859 10364 4167 10373
rect 3859 10362 3865 10364
rect 3921 10362 3945 10364
rect 4001 10362 4025 10364
rect 4081 10362 4105 10364
rect 4161 10362 4167 10364
rect 3921 10310 3923 10362
rect 4103 10310 4105 10362
rect 3859 10308 3865 10310
rect 3921 10308 3945 10310
rect 4001 10308 4025 10310
rect 4081 10308 4105 10310
rect 4161 10308 4167 10310
rect 1122 10296 1178 10305
rect 3859 10299 4167 10308
rect 5920 10266 5948 10542
rect 1122 10231 1178 10240
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 6472 10062 6500 10610
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 4519 9820 4827 9829
rect 4519 9818 4525 9820
rect 4581 9818 4605 9820
rect 4661 9818 4685 9820
rect 4741 9818 4765 9820
rect 4821 9818 4827 9820
rect 4581 9766 4583 9818
rect 4763 9766 4765 9818
rect 4519 9764 4525 9766
rect 4581 9764 4605 9766
rect 4661 9764 4685 9766
rect 4741 9764 4765 9766
rect 4821 9764 4827 9766
rect 4519 9755 4827 9764
rect 7116 9382 7144 11154
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 7208 10266 7236 11086
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 3859 9276 4167 9285
rect 3859 9274 3865 9276
rect 3921 9274 3945 9276
rect 4001 9274 4025 9276
rect 4081 9274 4105 9276
rect 4161 9274 4167 9276
rect 3921 9222 3923 9274
rect 4103 9222 4105 9274
rect 3859 9220 3865 9222
rect 3921 9220 3945 9222
rect 4001 9220 4025 9222
rect 4081 9220 4105 9222
rect 4161 9220 4167 9222
rect 3859 9211 4167 9220
rect 7116 9110 7144 9318
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 1214 8936 1270 8945
rect 1214 8871 1216 8880
rect 1268 8871 1270 8880
rect 6828 8900 6880 8906
rect 1216 8842 1268 8848
rect 6828 8842 6880 8848
rect 4519 8732 4827 8741
rect 4519 8730 4525 8732
rect 4581 8730 4605 8732
rect 4661 8730 4685 8732
rect 4741 8730 4765 8732
rect 4821 8730 4827 8732
rect 4581 8678 4583 8730
rect 4763 8678 4765 8730
rect 4519 8676 4525 8678
rect 4581 8676 4605 8678
rect 4661 8676 4685 8678
rect 4741 8676 4765 8678
rect 4821 8676 4827 8678
rect 4519 8667 4827 8676
rect 6840 8498 6868 8842
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 3859 8188 4167 8197
rect 3859 8186 3865 8188
rect 3921 8186 3945 8188
rect 4001 8186 4025 8188
rect 4081 8186 4105 8188
rect 4161 8186 4167 8188
rect 3921 8134 3923 8186
rect 4103 8134 4105 8186
rect 3859 8132 3865 8134
rect 3921 8132 3945 8134
rect 4001 8132 4025 8134
rect 4081 8132 4105 8134
rect 4161 8132 4167 8134
rect 3859 8123 4167 8132
rect 4519 7644 4827 7653
rect 4519 7642 4525 7644
rect 4581 7642 4605 7644
rect 4661 7642 4685 7644
rect 4741 7642 4765 7644
rect 4821 7642 4827 7644
rect 4581 7590 4583 7642
rect 4763 7590 4765 7642
rect 4519 7588 4525 7590
rect 4581 7588 4605 7590
rect 4661 7588 4685 7590
rect 4741 7588 4765 7590
rect 4821 7588 4827 7590
rect 4519 7579 4827 7588
rect 7300 7410 7328 8570
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 3859 7100 4167 7109
rect 3859 7098 3865 7100
rect 3921 7098 3945 7100
rect 4001 7098 4025 7100
rect 4081 7098 4105 7100
rect 4161 7098 4167 7100
rect 3921 7046 3923 7098
rect 4103 7046 4105 7098
rect 3859 7044 3865 7046
rect 3921 7044 3945 7046
rect 4001 7044 4025 7046
rect 4081 7044 4105 7046
rect 4161 7044 4167 7046
rect 3859 7035 4167 7044
rect 7300 6934 7328 7346
rect 7392 7002 7420 11086
rect 8498 10908 8806 10917
rect 8498 10906 8504 10908
rect 8560 10906 8584 10908
rect 8640 10906 8664 10908
rect 8720 10906 8744 10908
rect 8800 10906 8806 10908
rect 8560 10854 8562 10906
rect 8742 10854 8744 10906
rect 8498 10852 8504 10854
rect 8560 10852 8584 10854
rect 8640 10852 8664 10854
rect 8720 10852 8744 10854
rect 8800 10852 8806 10854
rect 8498 10843 8806 10852
rect 7472 10668 7524 10674
rect 7748 10668 7800 10674
rect 7524 10628 7696 10656
rect 7472 10610 7524 10616
rect 7668 10470 7696 10628
rect 8484 10668 8536 10674
rect 7748 10610 7800 10616
rect 8404 10628 8484 10656
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9110 7604 9862
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7472 8832 7524 8838
rect 7524 8780 7604 8786
rect 7472 8774 7604 8780
rect 7484 8758 7604 8774
rect 7576 8566 7604 8758
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 7206 7512 8230
rect 7576 7478 7604 8502
rect 7668 8294 7696 10406
rect 7760 9926 7788 10610
rect 7838 10364 8146 10373
rect 7838 10362 7844 10364
rect 7900 10362 7924 10364
rect 7980 10362 8004 10364
rect 8060 10362 8084 10364
rect 8140 10362 8146 10364
rect 7900 10310 7902 10362
rect 8082 10310 8084 10362
rect 7838 10308 7844 10310
rect 7900 10308 7924 10310
rect 7980 10308 8004 10310
rect 8060 10308 8084 10310
rect 8140 10308 8146 10310
rect 7838 10299 8146 10308
rect 8404 10130 8432 10628
rect 8484 10610 8536 10616
rect 8576 10668 8628 10674
rect 8864 10656 8892 11086
rect 8576 10610 8628 10616
rect 8772 10628 8892 10656
rect 8588 10554 8616 10610
rect 8496 10526 8616 10554
rect 8496 10470 8524 10526
rect 8772 10470 8800 10628
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8496 10198 8524 10406
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 8404 9674 8432 10066
rect 8588 10062 8616 10406
rect 8864 10062 8892 10406
rect 8956 10266 8984 11086
rect 9048 10742 9076 12106
rect 9140 11354 9168 13738
rect 9416 12306 9444 17546
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9508 13870 9536 14010
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9508 13326 9536 13806
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13394 9904 13670
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 10060 12850 10088 17478
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10152 13326 10180 13874
rect 10612 13870 10640 17750
rect 10980 17678 11008 19200
rect 11624 17678 11652 19200
rect 11817 17980 12125 17989
rect 11817 17978 11823 17980
rect 11879 17978 11903 17980
rect 11959 17978 11983 17980
rect 12039 17978 12063 17980
rect 12119 17978 12125 17980
rect 11879 17926 11881 17978
rect 12061 17926 12063 17978
rect 11817 17924 11823 17926
rect 11879 17924 11903 17926
rect 11959 17924 11983 17926
rect 12039 17924 12063 17926
rect 12119 17924 12125 17926
rect 11817 17915 12125 17924
rect 12268 17882 12296 19200
rect 15796 17980 16104 17989
rect 15796 17978 15802 17980
rect 15858 17978 15882 17980
rect 15938 17978 15962 17980
rect 16018 17978 16042 17980
rect 16098 17978 16104 17980
rect 15858 17926 15860 17978
rect 16040 17926 16042 17978
rect 15796 17924 15802 17926
rect 15858 17924 15882 17926
rect 15938 17924 15962 17926
rect 16018 17924 16042 17926
rect 16098 17924 16104 17926
rect 15796 17915 16104 17924
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10612 13326 10640 13806
rect 11072 13734 11100 14350
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13462 11100 13670
rect 11164 13530 11192 13806
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11256 13326 11284 14010
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9232 11830 9260 12174
rect 9324 11898 9352 12174
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8864 9926 8892 9998
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8498 9820 8806 9829
rect 8498 9818 8504 9820
rect 8560 9818 8584 9820
rect 8640 9818 8664 9820
rect 8720 9818 8744 9820
rect 8800 9818 8806 9820
rect 8560 9766 8562 9818
rect 8742 9766 8744 9818
rect 8498 9764 8504 9766
rect 8560 9764 8584 9766
rect 8640 9764 8664 9766
rect 8720 9764 8744 9766
rect 8800 9764 8806 9766
rect 8498 9755 8806 9764
rect 8312 9646 8432 9674
rect 7838 9276 8146 9285
rect 7838 9274 7844 9276
rect 7900 9274 7924 9276
rect 7980 9274 8004 9276
rect 8060 9274 8084 9276
rect 8140 9274 8146 9276
rect 7900 9222 7902 9274
rect 8082 9222 8084 9274
rect 7838 9220 7844 9222
rect 7900 9220 7924 9222
rect 7980 9220 8004 9222
rect 8060 9220 8084 9222
rect 8140 9220 8146 9222
rect 7838 9211 8146 9220
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8036 8634 8064 8910
rect 8220 8838 8248 9114
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8220 8378 8248 8774
rect 7944 8362 8248 8378
rect 8312 8362 8340 9646
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8680 9042 8708 9522
rect 8956 9178 8984 9522
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 9178 9076 9454
rect 9232 9450 9260 11766
rect 9968 11762 9996 12242
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9784 10674 9812 11018
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9876 10674 9904 10950
rect 10060 10810 10088 12786
rect 10152 12442 10180 13262
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10612 11762 10640 13262
rect 11348 12238 11376 17478
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10336 11014 10364 11698
rect 10704 11694 10732 12174
rect 11440 11898 11468 17546
rect 12477 17436 12785 17445
rect 12477 17434 12483 17436
rect 12539 17434 12563 17436
rect 12619 17434 12643 17436
rect 12699 17434 12723 17436
rect 12779 17434 12785 17436
rect 12539 17382 12541 17434
rect 12721 17382 12723 17434
rect 12477 17380 12483 17382
rect 12539 17380 12563 17382
rect 12619 17380 12643 17382
rect 12699 17380 12723 17382
rect 12779 17380 12785 17382
rect 12477 17371 12785 17380
rect 11817 16892 12125 16901
rect 11817 16890 11823 16892
rect 11879 16890 11903 16892
rect 11959 16890 11983 16892
rect 12039 16890 12063 16892
rect 12119 16890 12125 16892
rect 11879 16838 11881 16890
rect 12061 16838 12063 16890
rect 11817 16836 11823 16838
rect 11879 16836 11903 16838
rect 11959 16836 11983 16838
rect 12039 16836 12063 16838
rect 12119 16836 12125 16838
rect 11817 16827 12125 16836
rect 12477 16348 12785 16357
rect 12477 16346 12483 16348
rect 12539 16346 12563 16348
rect 12619 16346 12643 16348
rect 12699 16346 12723 16348
rect 12779 16346 12785 16348
rect 12539 16294 12541 16346
rect 12721 16294 12723 16346
rect 12477 16292 12483 16294
rect 12539 16292 12563 16294
rect 12619 16292 12643 16294
rect 12699 16292 12723 16294
rect 12779 16292 12785 16294
rect 12477 16283 12785 16292
rect 11817 15804 12125 15813
rect 11817 15802 11823 15804
rect 11879 15802 11903 15804
rect 11959 15802 11983 15804
rect 12039 15802 12063 15804
rect 12119 15802 12125 15804
rect 11879 15750 11881 15802
rect 12061 15750 12063 15802
rect 11817 15748 11823 15750
rect 11879 15748 11903 15750
rect 11959 15748 11983 15750
rect 12039 15748 12063 15750
rect 12119 15748 12125 15750
rect 11817 15739 12125 15748
rect 12477 15260 12785 15269
rect 12477 15258 12483 15260
rect 12539 15258 12563 15260
rect 12619 15258 12643 15260
rect 12699 15258 12723 15260
rect 12779 15258 12785 15260
rect 12539 15206 12541 15258
rect 12721 15206 12723 15258
rect 12477 15204 12483 15206
rect 12539 15204 12563 15206
rect 12619 15204 12643 15206
rect 12699 15204 12723 15206
rect 12779 15204 12785 15206
rect 12477 15195 12785 15204
rect 11817 14716 12125 14725
rect 11817 14714 11823 14716
rect 11879 14714 11903 14716
rect 11959 14714 11983 14716
rect 12039 14714 12063 14716
rect 12119 14714 12125 14716
rect 11879 14662 11881 14714
rect 12061 14662 12063 14714
rect 11817 14660 11823 14662
rect 11879 14660 11903 14662
rect 11959 14660 11983 14662
rect 12039 14660 12063 14662
rect 12119 14660 12125 14662
rect 11817 14651 12125 14660
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11532 14074 11560 14418
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11150 10732 11630
rect 10888 11354 10916 11698
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11072 11218 11100 11766
rect 11624 11762 11652 14214
rect 12477 14172 12785 14181
rect 12477 14170 12483 14172
rect 12539 14170 12563 14172
rect 12619 14170 12643 14172
rect 12699 14170 12723 14172
rect 12779 14170 12785 14172
rect 12539 14118 12541 14170
rect 12721 14118 12723 14170
rect 12477 14116 12483 14118
rect 12539 14116 12563 14118
rect 12619 14116 12643 14118
rect 12699 14116 12723 14118
rect 12779 14116 12785 14118
rect 12477 14107 12785 14116
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11716 13394 11744 13806
rect 11817 13628 12125 13637
rect 11817 13626 11823 13628
rect 11879 13626 11903 13628
rect 11959 13626 11983 13628
rect 12039 13626 12063 13628
rect 12119 13626 12125 13628
rect 11879 13574 11881 13626
rect 12061 13574 12063 13626
rect 11817 13572 11823 13574
rect 11879 13572 11903 13574
rect 11959 13572 11983 13574
rect 12039 13572 12063 13574
rect 12119 13572 12125 13574
rect 11817 13563 12125 13572
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11817 12540 12125 12549
rect 11817 12538 11823 12540
rect 11879 12538 11903 12540
rect 11959 12538 11983 12540
rect 12039 12538 12063 12540
rect 12119 12538 12125 12540
rect 11879 12486 11881 12538
rect 12061 12486 12063 12538
rect 11817 12484 11823 12486
rect 11879 12484 11903 12486
rect 11959 12484 11983 12486
rect 12039 12484 12063 12486
rect 12119 12484 12125 12486
rect 11817 12475 12125 12484
rect 12176 12442 12204 13806
rect 12477 13084 12785 13093
rect 12477 13082 12483 13084
rect 12539 13082 12563 13084
rect 12619 13082 12643 13084
rect 12699 13082 12723 13084
rect 12779 13082 12785 13084
rect 12539 13030 12541 13082
rect 12721 13030 12723 13082
rect 12477 13028 12483 13030
rect 12539 13028 12563 13030
rect 12619 13028 12643 13030
rect 12699 13028 12723 13030
rect 12779 13028 12785 13030
rect 12477 13019 12785 13028
rect 12820 12442 12848 17614
rect 16456 17436 16764 17445
rect 16456 17434 16462 17436
rect 16518 17434 16542 17436
rect 16598 17434 16622 17436
rect 16678 17434 16702 17436
rect 16758 17434 16764 17436
rect 16518 17382 16520 17434
rect 16700 17382 16702 17434
rect 16456 17380 16462 17382
rect 16518 17380 16542 17382
rect 16598 17380 16622 17382
rect 16678 17380 16702 17382
rect 16758 17380 16764 17382
rect 16456 17371 16764 17380
rect 15796 16892 16104 16901
rect 15796 16890 15802 16892
rect 15858 16890 15882 16892
rect 15938 16890 15962 16892
rect 16018 16890 16042 16892
rect 16098 16890 16104 16892
rect 15858 16838 15860 16890
rect 16040 16838 16042 16890
rect 15796 16836 15802 16838
rect 15858 16836 15882 16838
rect 15938 16836 15962 16838
rect 16018 16836 16042 16838
rect 16098 16836 16104 16838
rect 15796 16827 16104 16836
rect 16456 16348 16764 16357
rect 16456 16346 16462 16348
rect 16518 16346 16542 16348
rect 16598 16346 16622 16348
rect 16678 16346 16702 16348
rect 16758 16346 16764 16348
rect 16518 16294 16520 16346
rect 16700 16294 16702 16346
rect 16456 16292 16462 16294
rect 16518 16292 16542 16294
rect 16598 16292 16622 16294
rect 16678 16292 16702 16294
rect 16758 16292 16764 16294
rect 16456 16283 16764 16292
rect 15796 15804 16104 15813
rect 15796 15802 15802 15804
rect 15858 15802 15882 15804
rect 15938 15802 15962 15804
rect 16018 15802 16042 15804
rect 16098 15802 16104 15804
rect 15858 15750 15860 15802
rect 16040 15750 16042 15802
rect 15796 15748 15802 15750
rect 15858 15748 15882 15750
rect 15938 15748 15962 15750
rect 16018 15748 16042 15750
rect 16098 15748 16104 15750
rect 15796 15739 16104 15748
rect 16456 15260 16764 15269
rect 16456 15258 16462 15260
rect 16518 15258 16542 15260
rect 16598 15258 16622 15260
rect 16678 15258 16702 15260
rect 16758 15258 16764 15260
rect 16518 15206 16520 15258
rect 16700 15206 16702 15258
rect 16456 15204 16462 15206
rect 16518 15204 16542 15206
rect 16598 15204 16622 15206
rect 16678 15204 16702 15206
rect 16758 15204 16764 15206
rect 16456 15195 16764 15204
rect 15796 14716 16104 14725
rect 15796 14714 15802 14716
rect 15858 14714 15882 14716
rect 15938 14714 15962 14716
rect 16018 14714 16042 14716
rect 16098 14714 16104 14716
rect 15858 14662 15860 14714
rect 16040 14662 16042 14714
rect 15796 14660 15802 14662
rect 15858 14660 15882 14662
rect 15938 14660 15962 14662
rect 16018 14660 16042 14662
rect 16098 14660 16104 14662
rect 15796 14651 16104 14660
rect 16456 14172 16764 14181
rect 16456 14170 16462 14172
rect 16518 14170 16542 14172
rect 16598 14170 16622 14172
rect 16678 14170 16702 14172
rect 16758 14170 16764 14172
rect 16518 14118 16520 14170
rect 16700 14118 16702 14170
rect 16456 14116 16462 14118
rect 16518 14116 16542 14118
rect 16598 14116 16622 14118
rect 16678 14116 16702 14118
rect 16758 14116 16764 14118
rect 16456 14107 16764 14116
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13004 13530 13032 13874
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 12268 11898 12296 12174
rect 12477 11996 12785 12005
rect 12477 11994 12483 11996
rect 12539 11994 12563 11996
rect 12619 11994 12643 11996
rect 12699 11994 12723 11996
rect 12779 11994 12785 11996
rect 12539 11942 12541 11994
rect 12721 11942 12723 11994
rect 12477 11940 12483 11942
rect 12539 11940 12563 11942
rect 12619 11940 12643 11942
rect 12699 11940 12723 11942
rect 12779 11940 12785 11942
rect 12477 11931 12785 11940
rect 13188 11898 13216 12174
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 12820 11762 12848 11834
rect 13280 11830 13308 13262
rect 13372 12986 13400 13262
rect 13648 12986 13676 13262
rect 13740 13190 13768 13738
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10692 11144 10744 11150
rect 10612 11104 10692 11132
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10060 10674 10088 10746
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 9324 9654 9352 10610
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8956 8906 8984 8978
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 9048 8838 9076 9114
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8498 8732 8806 8741
rect 8498 8730 8504 8732
rect 8560 8730 8584 8732
rect 8640 8730 8664 8732
rect 8720 8730 8744 8732
rect 8800 8730 8806 8732
rect 8560 8678 8562 8730
rect 8742 8678 8744 8730
rect 8498 8676 8504 8678
rect 8560 8676 8584 8678
rect 8640 8676 8664 8678
rect 8720 8676 8744 8678
rect 8800 8676 8806 8678
rect 8498 8667 8806 8676
rect 9048 8634 9076 8774
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 7932 8356 8248 8362
rect 7984 8350 8248 8356
rect 7932 8298 7984 8304
rect 8220 8294 8248 8350
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7838 8188 8146 8197
rect 7838 8186 7844 8188
rect 7900 8186 7924 8188
rect 7980 8186 8004 8188
rect 8060 8186 8084 8188
rect 8140 8186 8146 8188
rect 7900 8134 7902 8186
rect 8082 8134 8084 8186
rect 7838 8132 7844 8134
rect 7900 8132 7924 8134
rect 7980 8132 8004 8134
rect 8060 8132 8084 8134
rect 8140 8132 8146 8134
rect 7838 8123 8146 8132
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7760 7546 7788 7754
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7564 7472 7616 7478
rect 7852 7426 7880 7482
rect 7564 7414 7616 7420
rect 7760 7398 7880 7426
rect 8208 7404 8260 7410
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7484 6866 7512 7142
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7668 6798 7696 7142
rect 7760 7002 7788 7398
rect 8208 7346 8260 7352
rect 7838 7100 8146 7109
rect 7838 7098 7844 7100
rect 7900 7098 7924 7100
rect 7980 7098 8004 7100
rect 8060 7098 8084 7100
rect 8140 7098 8146 7100
rect 7900 7046 7902 7098
rect 8082 7046 8084 7098
rect 7838 7044 7844 7046
rect 7900 7044 7924 7046
rect 7980 7044 8004 7046
rect 8060 7044 8084 7046
rect 8140 7044 8146 7046
rect 7838 7035 8146 7044
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7840 6928 7892 6934
rect 7760 6876 7840 6882
rect 7760 6870 7892 6876
rect 7760 6854 7880 6870
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 4519 6556 4827 6565
rect 4519 6554 4525 6556
rect 4581 6554 4605 6556
rect 4661 6554 4685 6556
rect 4741 6554 4765 6556
rect 4821 6554 4827 6556
rect 4581 6502 4583 6554
rect 4763 6502 4765 6554
rect 4519 6500 4525 6502
rect 4581 6500 4605 6502
rect 4661 6500 4685 6502
rect 4741 6500 4765 6502
rect 4821 6500 4827 6502
rect 4519 6491 4827 6500
rect 3859 6012 4167 6021
rect 3859 6010 3865 6012
rect 3921 6010 3945 6012
rect 4001 6010 4025 6012
rect 4081 6010 4105 6012
rect 4161 6010 4167 6012
rect 3921 5958 3923 6010
rect 4103 5958 4105 6010
rect 3859 5956 3865 5958
rect 3921 5956 3945 5958
rect 4001 5956 4025 5958
rect 4081 5956 4105 5958
rect 4161 5956 4167 5958
rect 3859 5947 4167 5956
rect 4519 5468 4827 5477
rect 4519 5466 4525 5468
rect 4581 5466 4605 5468
rect 4661 5466 4685 5468
rect 4741 5466 4765 5468
rect 4821 5466 4827 5468
rect 4581 5414 4583 5466
rect 4763 5414 4765 5466
rect 4519 5412 4525 5414
rect 4581 5412 4605 5414
rect 4661 5412 4685 5414
rect 4741 5412 4765 5414
rect 4821 5412 4827 5414
rect 4519 5403 4827 5412
rect 3859 4924 4167 4933
rect 3859 4922 3865 4924
rect 3921 4922 3945 4924
rect 4001 4922 4025 4924
rect 4081 4922 4105 4924
rect 4161 4922 4167 4924
rect 3921 4870 3923 4922
rect 4103 4870 4105 4922
rect 3859 4868 3865 4870
rect 3921 4868 3945 4870
rect 4001 4868 4025 4870
rect 4081 4868 4105 4870
rect 4161 4868 4167 4870
rect 3859 4859 4167 4868
rect 4519 4380 4827 4389
rect 4519 4378 4525 4380
rect 4581 4378 4605 4380
rect 4661 4378 4685 4380
rect 4741 4378 4765 4380
rect 4821 4378 4827 4380
rect 4581 4326 4583 4378
rect 4763 4326 4765 4378
rect 4519 4324 4525 4326
rect 4581 4324 4605 4326
rect 4661 4324 4685 4326
rect 4741 4324 4765 4326
rect 4821 4324 4827 4326
rect 4519 4315 4827 4324
rect 3859 3836 4167 3845
rect 3859 3834 3865 3836
rect 3921 3834 3945 3836
rect 4001 3834 4025 3836
rect 4081 3834 4105 3836
rect 4161 3834 4167 3836
rect 3921 3782 3923 3834
rect 4103 3782 4105 3834
rect 3859 3780 3865 3782
rect 3921 3780 3945 3782
rect 4001 3780 4025 3782
rect 4081 3780 4105 3782
rect 4161 3780 4167 3782
rect 3859 3771 4167 3780
rect 4519 3292 4827 3301
rect 4519 3290 4525 3292
rect 4581 3290 4605 3292
rect 4661 3290 4685 3292
rect 4741 3290 4765 3292
rect 4821 3290 4827 3292
rect 4581 3238 4583 3290
rect 4763 3238 4765 3290
rect 4519 3236 4525 3238
rect 4581 3236 4605 3238
rect 4661 3236 4685 3238
rect 4741 3236 4765 3238
rect 4821 3236 4827 3238
rect 4519 3227 4827 3236
rect 3859 2748 4167 2757
rect 3859 2746 3865 2748
rect 3921 2746 3945 2748
rect 4001 2746 4025 2748
rect 4081 2746 4105 2748
rect 4161 2746 4167 2748
rect 3921 2694 3923 2746
rect 4103 2694 4105 2746
rect 3859 2692 3865 2694
rect 3921 2692 3945 2694
rect 4001 2692 4025 2694
rect 4081 2692 4105 2694
rect 4161 2692 4167 2694
rect 3859 2683 4167 2692
rect 7760 2582 7788 6854
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6322 8064 6598
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8220 6186 8248 7346
rect 8404 7342 8432 8502
rect 9140 8498 9168 8978
rect 9416 8974 9444 9998
rect 9876 9654 9904 10610
rect 10244 10266 10272 10610
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10336 9994 10364 10950
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10520 10198 10548 10610
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10508 10056 10560 10062
rect 10612 10044 10640 11104
rect 10692 11086 10744 11092
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10810 10824 10950
rect 11256 10810 11284 11698
rect 11817 11452 12125 11461
rect 11817 11450 11823 11452
rect 11879 11450 11903 11452
rect 11959 11450 11983 11452
rect 12039 11450 12063 11452
rect 12119 11450 12125 11452
rect 11879 11398 11881 11450
rect 12061 11398 12063 11450
rect 11817 11396 11823 11398
rect 11879 11396 11903 11398
rect 11959 11396 11983 11398
rect 12039 11396 12063 11398
rect 12119 11396 12125 11398
rect 11817 11387 12125 11396
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11520 10668 11572 10674
rect 11572 10628 11652 10656
rect 11520 10610 11572 10616
rect 11072 10266 11100 10610
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11348 10198 11376 10610
rect 11624 10538 11652 10628
rect 11612 10532 11664 10538
rect 11612 10474 11664 10480
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11624 10130 11652 10474
rect 11817 10364 12125 10373
rect 11817 10362 11823 10364
rect 11879 10362 11903 10364
rect 11959 10362 11983 10364
rect 12039 10362 12063 10364
rect 12119 10362 12125 10364
rect 11879 10310 11881 10362
rect 12061 10310 12063 10362
rect 11817 10308 11823 10310
rect 11879 10308 11903 10310
rect 11959 10308 11983 10310
rect 12039 10308 12063 10310
rect 12119 10308 12125 10310
rect 11817 10299 12125 10308
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 10560 10016 10640 10044
rect 10692 10056 10744 10062
rect 10508 9998 10560 10004
rect 10692 9998 10744 10004
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9324 8498 9352 8842
rect 9416 8566 9444 8910
rect 9600 8634 9628 9590
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 8498 7644 8806 7653
rect 8498 7642 8504 7644
rect 8560 7642 8584 7644
rect 8640 7642 8664 7644
rect 8720 7642 8744 7644
rect 8800 7642 8806 7644
rect 8560 7590 8562 7642
rect 8742 7590 8744 7642
rect 8498 7588 8504 7590
rect 8560 7588 8584 7590
rect 8640 7588 8664 7590
rect 8720 7588 8744 7590
rect 8800 7588 8806 7590
rect 8498 7579 8806 7588
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 6322 8340 7142
rect 8404 6662 8432 7278
rect 8496 6934 8524 7346
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8496 6798 8524 6870
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8680 6730 8708 7210
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6338 8432 6598
rect 8498 6556 8806 6565
rect 8498 6554 8504 6556
rect 8560 6554 8584 6556
rect 8640 6554 8664 6556
rect 8720 6554 8744 6556
rect 8800 6554 8806 6556
rect 8560 6502 8562 6554
rect 8742 6502 8744 6554
rect 8498 6500 8504 6502
rect 8560 6500 8584 6502
rect 8640 6500 8664 6502
rect 8720 6500 8744 6502
rect 8800 6500 8806 6502
rect 8498 6491 8806 6500
rect 8864 6458 8892 6938
rect 8956 6798 8984 7142
rect 9048 6866 9076 8298
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8404 6322 8524 6338
rect 8300 6316 8352 6322
rect 8404 6316 8536 6322
rect 8404 6310 8484 6316
rect 8300 6258 8352 6264
rect 8484 6258 8536 6264
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 7838 6012 8146 6021
rect 7838 6010 7844 6012
rect 7900 6010 7924 6012
rect 7980 6010 8004 6012
rect 8060 6010 8084 6012
rect 8140 6010 8146 6012
rect 7900 5958 7902 6010
rect 8082 5958 8084 6010
rect 7838 5956 7844 5958
rect 7900 5956 7924 5958
rect 7980 5956 8004 5958
rect 8060 5956 8084 5958
rect 8140 5956 8146 5958
rect 7838 5947 8146 5956
rect 8498 5468 8806 5477
rect 8498 5466 8504 5468
rect 8560 5466 8584 5468
rect 8640 5466 8664 5468
rect 8720 5466 8744 5468
rect 8800 5466 8806 5468
rect 8560 5414 8562 5466
rect 8742 5414 8744 5466
rect 8498 5412 8504 5414
rect 8560 5412 8584 5414
rect 8640 5412 8664 5414
rect 8720 5412 8744 5414
rect 8800 5412 8806 5414
rect 8498 5403 8806 5412
rect 7838 4924 8146 4933
rect 7838 4922 7844 4924
rect 7900 4922 7924 4924
rect 7980 4922 8004 4924
rect 8060 4922 8084 4924
rect 8140 4922 8146 4924
rect 7900 4870 7902 4922
rect 8082 4870 8084 4922
rect 7838 4868 7844 4870
rect 7900 4868 7924 4870
rect 7980 4868 8004 4870
rect 8060 4868 8084 4870
rect 8140 4868 8146 4870
rect 7838 4859 8146 4868
rect 8498 4380 8806 4389
rect 8498 4378 8504 4380
rect 8560 4378 8584 4380
rect 8640 4378 8664 4380
rect 8720 4378 8744 4380
rect 8800 4378 8806 4380
rect 8560 4326 8562 4378
rect 8742 4326 8744 4378
rect 8498 4324 8504 4326
rect 8560 4324 8584 4326
rect 8640 4324 8664 4326
rect 8720 4324 8744 4326
rect 8800 4324 8806 4326
rect 8498 4315 8806 4324
rect 7838 3836 8146 3845
rect 7838 3834 7844 3836
rect 7900 3834 7924 3836
rect 7980 3834 8004 3836
rect 8060 3834 8084 3836
rect 8140 3834 8146 3836
rect 7900 3782 7902 3834
rect 8082 3782 8084 3834
rect 7838 3780 7844 3782
rect 7900 3780 7924 3782
rect 7980 3780 8004 3782
rect 8060 3780 8084 3782
rect 8140 3780 8146 3782
rect 7838 3771 8146 3780
rect 8498 3292 8806 3301
rect 8498 3290 8504 3292
rect 8560 3290 8584 3292
rect 8640 3290 8664 3292
rect 8720 3290 8744 3292
rect 8800 3290 8806 3292
rect 8560 3238 8562 3290
rect 8742 3238 8744 3290
rect 8498 3236 8504 3238
rect 8560 3236 8584 3238
rect 8640 3236 8664 3238
rect 8720 3236 8744 3238
rect 8800 3236 8806 3238
rect 8498 3227 8806 3236
rect 7838 2748 8146 2757
rect 7838 2746 7844 2748
rect 7900 2746 7924 2748
rect 7980 2746 8004 2748
rect 8060 2746 8084 2748
rect 8140 2746 8146 2748
rect 7900 2694 7902 2746
rect 8082 2694 8084 2746
rect 7838 2692 7844 2694
rect 7900 2692 7924 2694
rect 7980 2692 8004 2694
rect 8060 2692 8084 2694
rect 8140 2692 8146 2694
rect 7838 2683 8146 2692
rect 9140 2650 9168 8434
rect 9324 7410 9352 8434
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9692 7478 9720 8026
rect 10152 7954 10180 9318
rect 10244 8498 10272 9590
rect 10520 9586 10548 9862
rect 10704 9722 10732 9998
rect 10796 9926 10824 10066
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10796 9602 10824 9862
rect 10980 9654 11008 9998
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10704 9574 10824 9602
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10336 8956 10364 9046
rect 10508 8968 10560 8974
rect 10336 8928 10508 8956
rect 10508 8910 10560 8916
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8566 10640 8774
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10244 8090 10272 8434
rect 10704 8430 10732 9574
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 8838 10824 9318
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10980 8514 11008 9590
rect 11716 8906 11744 9998
rect 11992 9722 12020 10066
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 11817 9276 12125 9285
rect 11817 9274 11823 9276
rect 11879 9274 11903 9276
rect 11959 9274 11983 9276
rect 12039 9274 12063 9276
rect 12119 9274 12125 9276
rect 11879 9222 11881 9274
rect 12061 9222 12063 9274
rect 11817 9220 11823 9222
rect 11879 9220 11903 9222
rect 11959 9220 11983 9222
rect 12039 9220 12063 9222
rect 12119 9220 12125 9222
rect 11817 9211 12125 9220
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11060 8560 11112 8566
rect 10980 8508 11060 8514
rect 10980 8502 11112 8508
rect 10784 8492 10836 8498
rect 10980 8486 11100 8502
rect 11716 8498 11744 8842
rect 11704 8492 11756 8498
rect 10784 8434 10836 8440
rect 11704 8434 11756 8440
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10612 7954 10640 8366
rect 10140 7948 10192 7954
rect 10140 7890 10192 7896
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10692 7880 10744 7886
rect 10796 7834 10824 8434
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11072 7886 11100 8230
rect 11164 8022 11192 8298
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11256 8090 11284 8230
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11348 7936 11376 8230
rect 11256 7908 11376 7936
rect 10744 7828 10824 7834
rect 10692 7822 10824 7828
rect 11060 7880 11112 7886
rect 11256 7868 11284 7908
rect 11112 7840 11284 7868
rect 11060 7822 11112 7828
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9600 6730 9628 7346
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 4519 2204 4827 2213
rect 4519 2202 4525 2204
rect 4581 2202 4605 2204
rect 4661 2202 4685 2204
rect 4741 2202 4765 2204
rect 4821 2202 4827 2204
rect 4581 2150 4583 2202
rect 4763 2150 4765 2202
rect 4519 2148 4525 2150
rect 4581 2148 4605 2150
rect 4661 2148 4685 2150
rect 4741 2148 4765 2150
rect 4821 2148 4827 2150
rect 4519 2139 4827 2148
rect 7760 800 7788 2382
rect 8404 800 8432 2382
rect 8498 2204 8806 2213
rect 8498 2202 8504 2204
rect 8560 2202 8584 2204
rect 8640 2202 8664 2204
rect 8720 2202 8744 2204
rect 8800 2202 8806 2204
rect 8560 2150 8562 2202
rect 8742 2150 8744 2202
rect 8498 2148 8504 2150
rect 8560 2148 8584 2150
rect 8640 2148 8664 2150
rect 8720 2148 8744 2150
rect 8800 2148 8806 2150
rect 8498 2139 8806 2148
rect 9048 800 9076 2450
rect 9508 2446 9536 6598
rect 9876 6322 9904 6666
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 10152 2514 10180 6734
rect 10244 6458 10272 7822
rect 10704 7806 10824 7822
rect 10692 7744 10744 7750
rect 10796 7732 10824 7806
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 10968 7744 11020 7750
rect 10796 7704 10968 7732
rect 10692 7686 10744 7692
rect 10968 7686 11020 7692
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10704 3058 10732 7686
rect 10980 6322 11008 7686
rect 11348 7546 11376 7754
rect 11532 7750 11560 8298
rect 11716 7750 11744 8434
rect 12176 8378 12204 11154
rect 12452 11098 12480 11698
rect 12360 11070 12480 11098
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12268 9042 12296 9998
rect 12360 9926 12388 11070
rect 12820 11014 12848 11698
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11150 12940 11630
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12477 10908 12785 10917
rect 12477 10906 12483 10908
rect 12539 10906 12563 10908
rect 12619 10906 12643 10908
rect 12699 10906 12723 10908
rect 12779 10906 12785 10908
rect 12539 10854 12541 10906
rect 12721 10854 12723 10906
rect 12477 10852 12483 10854
rect 12539 10852 12563 10854
rect 12619 10852 12643 10854
rect 12699 10852 12723 10854
rect 12779 10852 12785 10854
rect 12477 10843 12785 10852
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10266 12480 10406
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12544 10062 12572 10134
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12636 9994 12664 10610
rect 12820 10470 12848 10950
rect 13004 10554 13032 11698
rect 13096 10810 13124 11698
rect 13188 11626 13216 11698
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12912 10526 13032 10554
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 10062 12848 10406
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12360 9602 12388 9862
rect 12477 9820 12785 9829
rect 12477 9818 12483 9820
rect 12539 9818 12563 9820
rect 12619 9818 12643 9820
rect 12699 9818 12723 9820
rect 12779 9818 12785 9820
rect 12539 9766 12541 9818
rect 12721 9766 12723 9818
rect 12477 9764 12483 9766
rect 12539 9764 12563 9766
rect 12619 9764 12643 9766
rect 12699 9764 12723 9766
rect 12779 9764 12785 9766
rect 12477 9755 12785 9764
rect 12360 9574 12572 9602
rect 12820 9586 12848 9862
rect 12912 9586 12940 10526
rect 13084 10056 13136 10062
rect 13188 10044 13216 11562
rect 13464 11354 13492 11698
rect 13556 11354 13584 12786
rect 13740 11626 13768 12786
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11898 13860 12242
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13556 10062 13584 11018
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13728 10736 13780 10742
rect 13728 10678 13780 10684
rect 13740 10198 13768 10678
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13740 10062 13768 10134
rect 13832 10062 13860 10950
rect 13136 10016 13216 10044
rect 13084 9998 13136 10004
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12544 9466 12572 9574
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12268 8566 12296 8978
rect 12452 8922 12480 9454
rect 12544 9438 13032 9466
rect 12360 8894 12480 8922
rect 12360 8634 12388 8894
rect 12477 8732 12785 8741
rect 12477 8730 12483 8732
rect 12539 8730 12563 8732
rect 12619 8730 12643 8732
rect 12699 8730 12723 8732
rect 12779 8730 12785 8732
rect 12539 8678 12541 8730
rect 12721 8678 12723 8730
rect 12477 8676 12483 8678
rect 12539 8676 12563 8678
rect 12619 8676 12643 8678
rect 12699 8676 12723 8678
rect 12779 8676 12785 8678
rect 12477 8667 12785 8676
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12176 8350 12388 8378
rect 11817 8188 12125 8197
rect 11817 8186 11823 8188
rect 11879 8186 11903 8188
rect 11959 8186 11983 8188
rect 12039 8186 12063 8188
rect 12119 8186 12125 8188
rect 11879 8134 11881 8186
rect 12061 8134 12063 8186
rect 11817 8132 11823 8134
rect 11879 8132 11903 8134
rect 11959 8132 11983 8134
rect 12039 8132 12063 8134
rect 12119 8132 12125 8134
rect 11817 8123 12125 8132
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 12176 7206 12204 7822
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 11817 7100 12125 7109
rect 11817 7098 11823 7100
rect 11879 7098 11903 7100
rect 11959 7098 11983 7100
rect 12039 7098 12063 7100
rect 12119 7098 12125 7100
rect 11879 7046 11881 7098
rect 12061 7046 12063 7098
rect 11817 7044 11823 7046
rect 11879 7044 11903 7046
rect 11959 7044 11983 7046
rect 12039 7044 12063 7046
rect 12119 7044 12125 7046
rect 11817 7035 12125 7044
rect 12176 7002 12204 7142
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 6866 12204 6938
rect 12360 6934 12388 8350
rect 12636 7954 12664 8570
rect 13004 7954 13032 9438
rect 13096 8974 13124 9862
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13096 8498 13124 8910
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13188 8294 13216 10016
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13280 8566 13308 9930
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13372 8430 13400 8774
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13556 8090 13584 8298
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13648 8022 13676 8230
rect 13832 8090 13860 8434
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 12624 7948 12676 7954
rect 12808 7948 12860 7954
rect 12624 7890 12676 7896
rect 12728 7908 12808 7936
rect 12728 7750 12756 7908
rect 12808 7890 12860 7896
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12477 7644 12785 7653
rect 12477 7642 12483 7644
rect 12539 7642 12563 7644
rect 12619 7642 12643 7644
rect 12699 7642 12723 7644
rect 12779 7642 12785 7644
rect 12539 7590 12541 7642
rect 12721 7590 12723 7642
rect 12477 7588 12483 7590
rect 12539 7588 12563 7590
rect 12619 7588 12643 7590
rect 12699 7588 12723 7590
rect 12779 7588 12785 7590
rect 12477 7579 12785 7588
rect 13372 7410 13400 7890
rect 13924 7546 13952 11086
rect 14016 9518 14044 13874
rect 15796 13628 16104 13637
rect 15796 13626 15802 13628
rect 15858 13626 15882 13628
rect 15938 13626 15962 13628
rect 16018 13626 16042 13628
rect 16098 13626 16104 13628
rect 15858 13574 15860 13626
rect 16040 13574 16042 13626
rect 15796 13572 15802 13574
rect 15858 13572 15882 13574
rect 15938 13572 15962 13574
rect 16018 13572 16042 13574
rect 16098 13572 16104 13574
rect 15796 13563 16104 13572
rect 16456 13084 16764 13093
rect 16456 13082 16462 13084
rect 16518 13082 16542 13084
rect 16598 13082 16622 13084
rect 16678 13082 16702 13084
rect 16758 13082 16764 13084
rect 16518 13030 16520 13082
rect 16700 13030 16702 13082
rect 16456 13028 16462 13030
rect 16518 13028 16542 13030
rect 16598 13028 16622 13030
rect 16678 13028 16702 13030
rect 16758 13028 16764 13030
rect 16456 13019 16764 13028
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 15796 12540 16104 12549
rect 15796 12538 15802 12540
rect 15858 12538 15882 12540
rect 15938 12538 15962 12540
rect 16018 12538 16042 12540
rect 16098 12538 16104 12540
rect 15858 12486 15860 12538
rect 16040 12486 16042 12538
rect 15796 12484 15802 12486
rect 15858 12484 15882 12486
rect 15938 12484 15962 12486
rect 16018 12484 16042 12486
rect 16098 12484 16104 12486
rect 15796 12475 16104 12484
rect 16500 12345 16528 12718
rect 16486 12336 16542 12345
rect 16486 12271 16542 12280
rect 16456 11996 16764 12005
rect 16456 11994 16462 11996
rect 16518 11994 16542 11996
rect 16598 11994 16622 11996
rect 16678 11994 16702 11996
rect 16758 11994 16764 11996
rect 16518 11942 16520 11994
rect 16700 11942 16702 11994
rect 16456 11940 16462 11942
rect 16518 11940 16542 11942
rect 16598 11940 16622 11942
rect 16678 11940 16702 11942
rect 16758 11940 16764 11942
rect 16456 11931 16764 11940
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14200 11218 14228 11562
rect 14292 11354 14320 11698
rect 17328 11665 17356 11698
rect 17314 11656 17370 11665
rect 14832 11620 14884 11626
rect 17314 11591 17370 11600
rect 14832 11562 14884 11568
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14844 11150 14872 11562
rect 15796 11452 16104 11461
rect 15796 11450 15802 11452
rect 15858 11450 15882 11452
rect 15938 11450 15962 11452
rect 16018 11450 16042 11452
rect 16098 11450 16104 11452
rect 15858 11398 15860 11450
rect 16040 11398 16042 11450
rect 15796 11396 15802 11398
rect 15858 11396 15882 11398
rect 15938 11396 15962 11398
rect 16018 11396 16042 11398
rect 16098 11396 16104 11398
rect 15796 11387 16104 11396
rect 17420 11354 17448 11766
rect 17408 11348 17460 11354
rect 17408 11290 17460 11296
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14476 10674 14504 10950
rect 14936 10674 14964 11222
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17512 10985 17540 11018
rect 17498 10976 17554 10985
rect 16456 10908 16764 10917
rect 17498 10911 17554 10920
rect 16456 10906 16462 10908
rect 16518 10906 16542 10908
rect 16598 10906 16622 10908
rect 16678 10906 16702 10908
rect 16758 10906 16764 10908
rect 16518 10854 16520 10906
rect 16700 10854 16702 10906
rect 16456 10852 16462 10854
rect 16518 10852 16542 10854
rect 16598 10852 16622 10854
rect 16678 10852 16702 10854
rect 16758 10852 16764 10854
rect 16456 10843 16764 10852
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 14844 10266 14872 10474
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14936 10198 14964 10610
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 15028 10062 15056 10406
rect 15120 10130 15148 10406
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15488 10062 15516 10474
rect 15796 10364 16104 10373
rect 15796 10362 15802 10364
rect 15858 10362 15882 10364
rect 15938 10362 15962 10364
rect 16018 10362 16042 10364
rect 16098 10362 16104 10364
rect 15858 10310 15860 10362
rect 16040 10310 16042 10362
rect 15796 10308 15802 10310
rect 15858 10308 15882 10310
rect 15938 10308 15962 10310
rect 16018 10308 16042 10310
rect 16098 10308 16104 10310
rect 15796 10299 16104 10308
rect 17420 10305 17448 10610
rect 17406 10296 17462 10305
rect 17406 10231 17462 10240
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 9586 14780 9862
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14476 8974 14504 9454
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14568 8922 14596 9454
rect 15212 8974 15240 9998
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15672 9654 15700 9862
rect 16456 9820 16764 9829
rect 16456 9818 16462 9820
rect 16518 9818 16542 9820
rect 16598 9818 16622 9820
rect 16678 9818 16702 9820
rect 16758 9818 16764 9820
rect 16518 9766 16520 9818
rect 16700 9766 16702 9818
rect 16456 9764 16462 9766
rect 16518 9764 16542 9766
rect 16598 9764 16622 9766
rect 16678 9764 16702 9766
rect 16758 9764 16764 9766
rect 16456 9755 16764 9764
rect 17328 9654 17356 9998
rect 17500 9920 17552 9926
rect 17500 9862 17552 9868
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 17316 9648 17368 9654
rect 17512 9625 17540 9862
rect 17316 9590 17368 9596
rect 17498 9616 17554 9625
rect 17498 9551 17554 9560
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15488 9178 15516 9454
rect 15796 9276 16104 9285
rect 15796 9274 15802 9276
rect 15858 9274 15882 9276
rect 15938 9274 15962 9276
rect 16018 9274 16042 9276
rect 16098 9274 16104 9276
rect 15858 9222 15860 9274
rect 16040 9222 16042 9274
rect 15796 9220 15802 9222
rect 15858 9220 15882 9222
rect 15938 9220 15962 9222
rect 16018 9220 16042 9222
rect 16098 9220 16104 9222
rect 15796 9211 16104 9220
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 14740 8968 14792 8974
rect 14004 8900 14056 8906
rect 14568 8894 14688 8922
rect 14740 8910 14792 8916
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 17498 8936 17554 8945
rect 14004 8842 14056 8848
rect 14016 7886 14044 8842
rect 14660 8838 14688 8894
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14660 8498 14688 8774
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14384 7478 14412 7686
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 11624 6662 11652 6802
rect 12072 6724 12124 6730
rect 12176 6712 12204 6802
rect 12360 6798 12388 6870
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12124 6684 12204 6712
rect 12072 6666 12124 6672
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11164 6322 11192 6598
rect 11992 6322 12020 6598
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 10980 5642 11008 6258
rect 11164 6118 11192 6258
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5710 11192 6054
rect 11440 5846 11468 6190
rect 11532 5914 11560 6258
rect 11817 6012 12125 6021
rect 11817 6010 11823 6012
rect 11879 6010 11903 6012
rect 11959 6010 11983 6012
rect 12039 6010 12063 6012
rect 12119 6010 12125 6012
rect 11879 5958 11881 6010
rect 12061 5958 12063 6010
rect 11817 5956 11823 5958
rect 11879 5956 11903 5958
rect 11959 5956 11983 5958
rect 12039 5956 12063 5958
rect 12119 5956 12125 5958
rect 11817 5947 12125 5956
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 800 9720 2246
rect 10336 800 10364 2790
rect 11256 2650 11284 5578
rect 11817 4924 12125 4933
rect 11817 4922 11823 4924
rect 11879 4922 11903 4924
rect 11959 4922 11983 4924
rect 12039 4922 12063 4924
rect 12119 4922 12125 4924
rect 11879 4870 11881 4922
rect 12061 4870 12063 4922
rect 11817 4868 11823 4870
rect 11879 4868 11903 4870
rect 11959 4868 11983 4870
rect 12039 4868 12063 4870
rect 12119 4868 12125 4870
rect 11817 4859 12125 4868
rect 11817 3836 12125 3845
rect 11817 3834 11823 3836
rect 11879 3834 11903 3836
rect 11959 3834 11983 3836
rect 12039 3834 12063 3836
rect 12119 3834 12125 3836
rect 11879 3782 11881 3834
rect 12061 3782 12063 3834
rect 11817 3780 11823 3782
rect 11879 3780 11903 3782
rect 11959 3780 11983 3782
rect 12039 3780 12063 3782
rect 12119 3780 12125 3782
rect 11817 3771 12125 3780
rect 11817 2748 12125 2757
rect 11817 2746 11823 2748
rect 11879 2746 11903 2748
rect 11959 2746 11983 2748
rect 12039 2746 12063 2748
rect 12119 2746 12125 2748
rect 11879 2694 11881 2746
rect 12061 2694 12063 2746
rect 11817 2692 11823 2694
rect 11879 2692 11903 2694
rect 11959 2692 11983 2694
rect 12039 2692 12063 2694
rect 12119 2692 12125 2694
rect 11817 2683 12125 2692
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 12176 2582 12204 6684
rect 12360 6662 12388 6734
rect 12820 6730 12848 7278
rect 13372 6866 13400 7346
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 7002 14136 7142
rect 14568 7002 14596 7414
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12477 6556 12785 6565
rect 12477 6554 12483 6556
rect 12539 6554 12563 6556
rect 12619 6554 12643 6556
rect 12699 6554 12723 6556
rect 12779 6554 12785 6556
rect 12539 6502 12541 6554
rect 12721 6502 12723 6554
rect 12477 6500 12483 6502
rect 12539 6500 12563 6502
rect 12619 6500 12643 6502
rect 12699 6500 12723 6502
rect 12779 6500 12785 6502
rect 12477 6491 12785 6500
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12268 5642 12296 6190
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 12477 5468 12785 5477
rect 12477 5466 12483 5468
rect 12539 5466 12563 5468
rect 12619 5466 12643 5468
rect 12699 5466 12723 5468
rect 12779 5466 12785 5468
rect 12539 5414 12541 5466
rect 12721 5414 12723 5466
rect 12477 5412 12483 5414
rect 12539 5412 12563 5414
rect 12619 5412 12643 5414
rect 12699 5412 12723 5414
rect 12779 5412 12785 5414
rect 12477 5403 12785 5412
rect 12477 4380 12785 4389
rect 12477 4378 12483 4380
rect 12539 4378 12563 4380
rect 12619 4378 12643 4380
rect 12699 4378 12723 4380
rect 12779 4378 12785 4380
rect 12539 4326 12541 4378
rect 12721 4326 12723 4378
rect 12477 4324 12483 4326
rect 12539 4324 12563 4326
rect 12619 4324 12643 4326
rect 12699 4324 12723 4326
rect 12779 4324 12785 4326
rect 12477 4315 12785 4324
rect 12477 3292 12785 3301
rect 12477 3290 12483 3292
rect 12539 3290 12563 3292
rect 12619 3290 12643 3292
rect 12699 3290 12723 3292
rect 12779 3290 12785 3292
rect 12539 3238 12541 3290
rect 12721 3238 12723 3290
rect 12477 3236 12483 3238
rect 12539 3236 12563 3238
rect 12619 3236 12643 3238
rect 12699 3236 12723 3238
rect 12779 3236 12785 3238
rect 12477 3227 12785 3236
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 12820 2514 12848 6666
rect 14660 6458 14688 8434
rect 14752 8430 14780 8910
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14752 8090 14780 8366
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 15212 7886 15240 8910
rect 17498 8871 17500 8880
rect 17552 8871 17554 8880
rect 17500 8842 17552 8848
rect 16456 8732 16764 8741
rect 16456 8730 16462 8732
rect 16518 8730 16542 8732
rect 16598 8730 16622 8732
rect 16678 8730 16702 8732
rect 16758 8730 16764 8732
rect 16518 8678 16520 8730
rect 16700 8678 16702 8730
rect 16456 8676 16462 8678
rect 16518 8676 16542 8678
rect 16598 8676 16622 8678
rect 16678 8676 16702 8678
rect 16758 8676 16764 8678
rect 16456 8667 16764 8676
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17328 8265 17356 8298
rect 17314 8256 17370 8265
rect 15796 8188 16104 8197
rect 17314 8191 17370 8200
rect 15796 8186 15802 8188
rect 15858 8186 15882 8188
rect 15938 8186 15962 8188
rect 16018 8186 16042 8188
rect 16098 8186 16104 8188
rect 15858 8134 15860 8186
rect 16040 8134 16042 8186
rect 15796 8132 15802 8134
rect 15858 8132 15882 8134
rect 15938 8132 15962 8134
rect 16018 8132 16042 8134
rect 16098 8132 16104 8134
rect 15796 8123 16104 8132
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 14752 7546 14780 7822
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14844 7002 14872 7346
rect 15212 7274 15240 7822
rect 16456 7644 16764 7653
rect 16456 7642 16462 7644
rect 16518 7642 16542 7644
rect 16598 7642 16622 7644
rect 16678 7642 16702 7644
rect 16758 7642 16764 7644
rect 16518 7590 16520 7642
rect 16700 7590 16702 7642
rect 16456 7588 16462 7590
rect 16518 7588 16542 7590
rect 16598 7588 16622 7590
rect 16678 7588 16702 7590
rect 16758 7588 16764 7590
rect 16456 7579 16764 7588
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15796 7100 16104 7109
rect 15796 7098 15802 7100
rect 15858 7098 15882 7100
rect 15938 7098 15962 7100
rect 16018 7098 16042 7100
rect 16098 7098 16104 7100
rect 15858 7046 15860 7098
rect 16040 7046 16042 7098
rect 15796 7044 15802 7046
rect 15858 7044 15882 7046
rect 15938 7044 15962 7046
rect 16018 7044 16042 7046
rect 16098 7044 16104 7046
rect 15796 7035 16104 7044
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 17328 6798 17356 7822
rect 17604 7585 17632 7822
rect 17590 7576 17646 7585
rect 17590 7511 17646 7520
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 16456 6556 16764 6565
rect 16456 6554 16462 6556
rect 16518 6554 16542 6556
rect 16598 6554 16622 6556
rect 16678 6554 16702 6556
rect 16758 6554 16764 6556
rect 16518 6502 16520 6554
rect 16700 6502 16702 6554
rect 16456 6500 16462 6502
rect 16518 6500 16542 6502
rect 16598 6500 16622 6502
rect 16678 6500 16702 6502
rect 16758 6500 16764 6502
rect 16456 6491 16764 6500
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 15796 6012 16104 6021
rect 15796 6010 15802 6012
rect 15858 6010 15882 6012
rect 15938 6010 15962 6012
rect 16018 6010 16042 6012
rect 16098 6010 16104 6012
rect 15858 5958 15860 6010
rect 16040 5958 16042 6010
rect 15796 5956 15802 5958
rect 15858 5956 15882 5958
rect 15938 5956 15962 5958
rect 16018 5956 16042 5958
rect 16098 5956 16104 5958
rect 15796 5947 16104 5956
rect 16456 5468 16764 5477
rect 16456 5466 16462 5468
rect 16518 5466 16542 5468
rect 16598 5466 16622 5468
rect 16678 5466 16702 5468
rect 16758 5466 16764 5468
rect 16518 5414 16520 5466
rect 16700 5414 16702 5466
rect 16456 5412 16462 5414
rect 16518 5412 16542 5414
rect 16598 5412 16622 5414
rect 16678 5412 16702 5414
rect 16758 5412 16764 5414
rect 16456 5403 16764 5412
rect 15796 4924 16104 4933
rect 15796 4922 15802 4924
rect 15858 4922 15882 4924
rect 15938 4922 15962 4924
rect 16018 4922 16042 4924
rect 16098 4922 16104 4924
rect 15858 4870 15860 4922
rect 16040 4870 16042 4922
rect 15796 4868 15802 4870
rect 15858 4868 15882 4870
rect 15938 4868 15962 4870
rect 16018 4868 16042 4870
rect 16098 4868 16104 4870
rect 15796 4859 16104 4868
rect 16456 4380 16764 4389
rect 16456 4378 16462 4380
rect 16518 4378 16542 4380
rect 16598 4378 16622 4380
rect 16678 4378 16702 4380
rect 16758 4378 16764 4380
rect 16518 4326 16520 4378
rect 16700 4326 16702 4378
rect 16456 4324 16462 4326
rect 16518 4324 16542 4326
rect 16598 4324 16622 4326
rect 16678 4324 16702 4326
rect 16758 4324 16764 4326
rect 16456 4315 16764 4324
rect 15796 3836 16104 3845
rect 15796 3834 15802 3836
rect 15858 3834 15882 3836
rect 15938 3834 15962 3836
rect 16018 3834 16042 3836
rect 16098 3834 16104 3836
rect 15858 3782 15860 3834
rect 16040 3782 16042 3834
rect 15796 3780 15802 3782
rect 15858 3780 15882 3782
rect 15938 3780 15962 3782
rect 16018 3780 16042 3782
rect 16098 3780 16104 3782
rect 15796 3771 16104 3780
rect 16456 3292 16764 3301
rect 16456 3290 16462 3292
rect 16518 3290 16542 3292
rect 16598 3290 16622 3292
rect 16678 3290 16702 3292
rect 16758 3290 16764 3292
rect 16518 3238 16520 3290
rect 16700 3238 16702 3290
rect 16456 3236 16462 3238
rect 16518 3236 16542 3238
rect 16598 3236 16622 3238
rect 16678 3236 16702 3238
rect 16758 3236 16764 3238
rect 16456 3227 16764 3236
rect 15796 2748 16104 2757
rect 15796 2746 15802 2748
rect 15858 2746 15882 2748
rect 15938 2746 15962 2748
rect 16018 2746 16042 2748
rect 16098 2746 16104 2748
rect 15858 2694 15860 2746
rect 16040 2694 16042 2746
rect 15796 2692 15802 2694
rect 15858 2692 15882 2694
rect 15938 2692 15962 2694
rect 16018 2692 16042 2694
rect 16098 2692 16104 2694
rect 15796 2683 16104 2692
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 10980 800 11008 2382
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11624 800 11652 2314
rect 12268 800 12296 2382
rect 12477 2204 12785 2213
rect 12477 2202 12483 2204
rect 12539 2202 12563 2204
rect 12619 2202 12643 2204
rect 12699 2202 12723 2204
rect 12779 2202 12785 2204
rect 12539 2150 12541 2202
rect 12721 2150 12723 2202
rect 12477 2148 12483 2150
rect 12539 2148 12563 2150
rect 12619 2148 12643 2150
rect 12699 2148 12723 2150
rect 12779 2148 12785 2150
rect 12477 2139 12785 2148
rect 16456 2204 16764 2213
rect 16456 2202 16462 2204
rect 16518 2202 16542 2204
rect 16598 2202 16622 2204
rect 16678 2202 16702 2204
rect 16758 2202 16764 2204
rect 16518 2150 16520 2202
rect 16700 2150 16702 2202
rect 16456 2148 16462 2150
rect 16518 2148 16542 2150
rect 16598 2148 16622 2150
rect 16678 2148 16702 2150
rect 16758 2148 16764 2150
rect 16456 2139 16764 2148
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
<< via2 >>
rect 3865 17978 3921 17980
rect 3945 17978 4001 17980
rect 4025 17978 4081 17980
rect 4105 17978 4161 17980
rect 3865 17926 3911 17978
rect 3911 17926 3921 17978
rect 3945 17926 3975 17978
rect 3975 17926 3987 17978
rect 3987 17926 4001 17978
rect 4025 17926 4039 17978
rect 4039 17926 4051 17978
rect 4051 17926 4081 17978
rect 4105 17926 4115 17978
rect 4115 17926 4161 17978
rect 3865 17924 3921 17926
rect 3945 17924 4001 17926
rect 4025 17924 4081 17926
rect 4105 17924 4161 17926
rect 7844 17978 7900 17980
rect 7924 17978 7980 17980
rect 8004 17978 8060 17980
rect 8084 17978 8140 17980
rect 7844 17926 7890 17978
rect 7890 17926 7900 17978
rect 7924 17926 7954 17978
rect 7954 17926 7966 17978
rect 7966 17926 7980 17978
rect 8004 17926 8018 17978
rect 8018 17926 8030 17978
rect 8030 17926 8060 17978
rect 8084 17926 8094 17978
rect 8094 17926 8140 17978
rect 7844 17924 7900 17926
rect 7924 17924 7980 17926
rect 8004 17924 8060 17926
rect 8084 17924 8140 17926
rect 4525 17434 4581 17436
rect 4605 17434 4661 17436
rect 4685 17434 4741 17436
rect 4765 17434 4821 17436
rect 4525 17382 4571 17434
rect 4571 17382 4581 17434
rect 4605 17382 4635 17434
rect 4635 17382 4647 17434
rect 4647 17382 4661 17434
rect 4685 17382 4699 17434
rect 4699 17382 4711 17434
rect 4711 17382 4741 17434
rect 4765 17382 4775 17434
rect 4775 17382 4821 17434
rect 4525 17380 4581 17382
rect 4605 17380 4661 17382
rect 4685 17380 4741 17382
rect 4765 17380 4821 17382
rect 8504 17434 8560 17436
rect 8584 17434 8640 17436
rect 8664 17434 8720 17436
rect 8744 17434 8800 17436
rect 8504 17382 8550 17434
rect 8550 17382 8560 17434
rect 8584 17382 8614 17434
rect 8614 17382 8626 17434
rect 8626 17382 8640 17434
rect 8664 17382 8678 17434
rect 8678 17382 8690 17434
rect 8690 17382 8720 17434
rect 8744 17382 8754 17434
rect 8754 17382 8800 17434
rect 8504 17380 8560 17382
rect 8584 17380 8640 17382
rect 8664 17380 8720 17382
rect 8744 17380 8800 17382
rect 3865 16890 3921 16892
rect 3945 16890 4001 16892
rect 4025 16890 4081 16892
rect 4105 16890 4161 16892
rect 3865 16838 3911 16890
rect 3911 16838 3921 16890
rect 3945 16838 3975 16890
rect 3975 16838 3987 16890
rect 3987 16838 4001 16890
rect 4025 16838 4039 16890
rect 4039 16838 4051 16890
rect 4051 16838 4081 16890
rect 4105 16838 4115 16890
rect 4115 16838 4161 16890
rect 3865 16836 3921 16838
rect 3945 16836 4001 16838
rect 4025 16836 4081 16838
rect 4105 16836 4161 16838
rect 7844 16890 7900 16892
rect 7924 16890 7980 16892
rect 8004 16890 8060 16892
rect 8084 16890 8140 16892
rect 7844 16838 7890 16890
rect 7890 16838 7900 16890
rect 7924 16838 7954 16890
rect 7954 16838 7966 16890
rect 7966 16838 7980 16890
rect 8004 16838 8018 16890
rect 8018 16838 8030 16890
rect 8030 16838 8060 16890
rect 8084 16838 8094 16890
rect 8094 16838 8140 16890
rect 7844 16836 7900 16838
rect 7924 16836 7980 16838
rect 8004 16836 8060 16838
rect 8084 16836 8140 16838
rect 4525 16346 4581 16348
rect 4605 16346 4661 16348
rect 4685 16346 4741 16348
rect 4765 16346 4821 16348
rect 4525 16294 4571 16346
rect 4571 16294 4581 16346
rect 4605 16294 4635 16346
rect 4635 16294 4647 16346
rect 4647 16294 4661 16346
rect 4685 16294 4699 16346
rect 4699 16294 4711 16346
rect 4711 16294 4741 16346
rect 4765 16294 4775 16346
rect 4775 16294 4821 16346
rect 4525 16292 4581 16294
rect 4605 16292 4661 16294
rect 4685 16292 4741 16294
rect 4765 16292 4821 16294
rect 8504 16346 8560 16348
rect 8584 16346 8640 16348
rect 8664 16346 8720 16348
rect 8744 16346 8800 16348
rect 8504 16294 8550 16346
rect 8550 16294 8560 16346
rect 8584 16294 8614 16346
rect 8614 16294 8626 16346
rect 8626 16294 8640 16346
rect 8664 16294 8678 16346
rect 8678 16294 8690 16346
rect 8690 16294 8720 16346
rect 8744 16294 8754 16346
rect 8754 16294 8800 16346
rect 8504 16292 8560 16294
rect 8584 16292 8640 16294
rect 8664 16292 8720 16294
rect 8744 16292 8800 16294
rect 3865 15802 3921 15804
rect 3945 15802 4001 15804
rect 4025 15802 4081 15804
rect 4105 15802 4161 15804
rect 3865 15750 3911 15802
rect 3911 15750 3921 15802
rect 3945 15750 3975 15802
rect 3975 15750 3987 15802
rect 3987 15750 4001 15802
rect 4025 15750 4039 15802
rect 4039 15750 4051 15802
rect 4051 15750 4081 15802
rect 4105 15750 4115 15802
rect 4115 15750 4161 15802
rect 3865 15748 3921 15750
rect 3945 15748 4001 15750
rect 4025 15748 4081 15750
rect 4105 15748 4161 15750
rect 7844 15802 7900 15804
rect 7924 15802 7980 15804
rect 8004 15802 8060 15804
rect 8084 15802 8140 15804
rect 7844 15750 7890 15802
rect 7890 15750 7900 15802
rect 7924 15750 7954 15802
rect 7954 15750 7966 15802
rect 7966 15750 7980 15802
rect 8004 15750 8018 15802
rect 8018 15750 8030 15802
rect 8030 15750 8060 15802
rect 8084 15750 8094 15802
rect 8094 15750 8140 15802
rect 7844 15748 7900 15750
rect 7924 15748 7980 15750
rect 8004 15748 8060 15750
rect 8084 15748 8140 15750
rect 4525 15258 4581 15260
rect 4605 15258 4661 15260
rect 4685 15258 4741 15260
rect 4765 15258 4821 15260
rect 4525 15206 4571 15258
rect 4571 15206 4581 15258
rect 4605 15206 4635 15258
rect 4635 15206 4647 15258
rect 4647 15206 4661 15258
rect 4685 15206 4699 15258
rect 4699 15206 4711 15258
rect 4711 15206 4741 15258
rect 4765 15206 4775 15258
rect 4775 15206 4821 15258
rect 4525 15204 4581 15206
rect 4605 15204 4661 15206
rect 4685 15204 4741 15206
rect 4765 15204 4821 15206
rect 8504 15258 8560 15260
rect 8584 15258 8640 15260
rect 8664 15258 8720 15260
rect 8744 15258 8800 15260
rect 8504 15206 8550 15258
rect 8550 15206 8560 15258
rect 8584 15206 8614 15258
rect 8614 15206 8626 15258
rect 8626 15206 8640 15258
rect 8664 15206 8678 15258
rect 8678 15206 8690 15258
rect 8690 15206 8720 15258
rect 8744 15206 8754 15258
rect 8754 15206 8800 15258
rect 8504 15204 8560 15206
rect 8584 15204 8640 15206
rect 8664 15204 8720 15206
rect 8744 15204 8800 15206
rect 3865 14714 3921 14716
rect 3945 14714 4001 14716
rect 4025 14714 4081 14716
rect 4105 14714 4161 14716
rect 3865 14662 3911 14714
rect 3911 14662 3921 14714
rect 3945 14662 3975 14714
rect 3975 14662 3987 14714
rect 3987 14662 4001 14714
rect 4025 14662 4039 14714
rect 4039 14662 4051 14714
rect 4051 14662 4081 14714
rect 4105 14662 4115 14714
rect 4115 14662 4161 14714
rect 3865 14660 3921 14662
rect 3945 14660 4001 14662
rect 4025 14660 4081 14662
rect 4105 14660 4161 14662
rect 7844 14714 7900 14716
rect 7924 14714 7980 14716
rect 8004 14714 8060 14716
rect 8084 14714 8140 14716
rect 7844 14662 7890 14714
rect 7890 14662 7900 14714
rect 7924 14662 7954 14714
rect 7954 14662 7966 14714
rect 7966 14662 7980 14714
rect 8004 14662 8018 14714
rect 8018 14662 8030 14714
rect 8030 14662 8060 14714
rect 8084 14662 8094 14714
rect 8094 14662 8140 14714
rect 7844 14660 7900 14662
rect 7924 14660 7980 14662
rect 8004 14660 8060 14662
rect 8084 14660 8140 14662
rect 4525 14170 4581 14172
rect 4605 14170 4661 14172
rect 4685 14170 4741 14172
rect 4765 14170 4821 14172
rect 4525 14118 4571 14170
rect 4571 14118 4581 14170
rect 4605 14118 4635 14170
rect 4635 14118 4647 14170
rect 4647 14118 4661 14170
rect 4685 14118 4699 14170
rect 4699 14118 4711 14170
rect 4711 14118 4741 14170
rect 4765 14118 4775 14170
rect 4775 14118 4821 14170
rect 4525 14116 4581 14118
rect 4605 14116 4661 14118
rect 4685 14116 4741 14118
rect 4765 14116 4821 14118
rect 8504 14170 8560 14172
rect 8584 14170 8640 14172
rect 8664 14170 8720 14172
rect 8744 14170 8800 14172
rect 8504 14118 8550 14170
rect 8550 14118 8560 14170
rect 8584 14118 8614 14170
rect 8614 14118 8626 14170
rect 8626 14118 8640 14170
rect 8664 14118 8678 14170
rect 8678 14118 8690 14170
rect 8690 14118 8720 14170
rect 8744 14118 8754 14170
rect 8754 14118 8800 14170
rect 8504 14116 8560 14118
rect 8584 14116 8640 14118
rect 8664 14116 8720 14118
rect 8744 14116 8800 14118
rect 3865 13626 3921 13628
rect 3945 13626 4001 13628
rect 4025 13626 4081 13628
rect 4105 13626 4161 13628
rect 3865 13574 3911 13626
rect 3911 13574 3921 13626
rect 3945 13574 3975 13626
rect 3975 13574 3987 13626
rect 3987 13574 4001 13626
rect 4025 13574 4039 13626
rect 4039 13574 4051 13626
rect 4051 13574 4081 13626
rect 4105 13574 4115 13626
rect 4115 13574 4161 13626
rect 3865 13572 3921 13574
rect 3945 13572 4001 13574
rect 4025 13572 4081 13574
rect 4105 13572 4161 13574
rect 7844 13626 7900 13628
rect 7924 13626 7980 13628
rect 8004 13626 8060 13628
rect 8084 13626 8140 13628
rect 7844 13574 7890 13626
rect 7890 13574 7900 13626
rect 7924 13574 7954 13626
rect 7954 13574 7966 13626
rect 7966 13574 7980 13626
rect 8004 13574 8018 13626
rect 8018 13574 8030 13626
rect 8030 13574 8060 13626
rect 8084 13574 8094 13626
rect 8094 13574 8140 13626
rect 7844 13572 7900 13574
rect 7924 13572 7980 13574
rect 8004 13572 8060 13574
rect 8084 13572 8140 13574
rect 4525 13082 4581 13084
rect 4605 13082 4661 13084
rect 4685 13082 4741 13084
rect 4765 13082 4821 13084
rect 4525 13030 4571 13082
rect 4571 13030 4581 13082
rect 4605 13030 4635 13082
rect 4635 13030 4647 13082
rect 4647 13030 4661 13082
rect 4685 13030 4699 13082
rect 4699 13030 4711 13082
rect 4711 13030 4741 13082
rect 4765 13030 4775 13082
rect 4775 13030 4821 13082
rect 4525 13028 4581 13030
rect 4605 13028 4661 13030
rect 4685 13028 4741 13030
rect 4765 13028 4821 13030
rect 8504 13082 8560 13084
rect 8584 13082 8640 13084
rect 8664 13082 8720 13084
rect 8744 13082 8800 13084
rect 8504 13030 8550 13082
rect 8550 13030 8560 13082
rect 8584 13030 8614 13082
rect 8614 13030 8626 13082
rect 8626 13030 8640 13082
rect 8664 13030 8678 13082
rect 8678 13030 8690 13082
rect 8690 13030 8720 13082
rect 8744 13030 8754 13082
rect 8754 13030 8800 13082
rect 8504 13028 8560 13030
rect 8584 13028 8640 13030
rect 8664 13028 8720 13030
rect 8744 13028 8800 13030
rect 3865 12538 3921 12540
rect 3945 12538 4001 12540
rect 4025 12538 4081 12540
rect 4105 12538 4161 12540
rect 3865 12486 3911 12538
rect 3911 12486 3921 12538
rect 3945 12486 3975 12538
rect 3975 12486 3987 12538
rect 3987 12486 4001 12538
rect 4025 12486 4039 12538
rect 4039 12486 4051 12538
rect 4051 12486 4081 12538
rect 4105 12486 4115 12538
rect 4115 12486 4161 12538
rect 3865 12484 3921 12486
rect 3945 12484 4001 12486
rect 4025 12484 4081 12486
rect 4105 12484 4161 12486
rect 7844 12538 7900 12540
rect 7924 12538 7980 12540
rect 8004 12538 8060 12540
rect 8084 12538 8140 12540
rect 7844 12486 7890 12538
rect 7890 12486 7900 12538
rect 7924 12486 7954 12538
rect 7954 12486 7966 12538
rect 7966 12486 7980 12538
rect 8004 12486 8018 12538
rect 8018 12486 8030 12538
rect 8030 12486 8060 12538
rect 8084 12486 8094 12538
rect 8094 12486 8140 12538
rect 7844 12484 7900 12486
rect 7924 12484 7980 12486
rect 8004 12484 8060 12486
rect 8084 12484 8140 12486
rect 2410 12280 2466 12336
rect 4525 11994 4581 11996
rect 4605 11994 4661 11996
rect 4685 11994 4741 11996
rect 4765 11994 4821 11996
rect 4525 11942 4571 11994
rect 4571 11942 4581 11994
rect 4605 11942 4635 11994
rect 4635 11942 4647 11994
rect 4647 11942 4661 11994
rect 4685 11942 4699 11994
rect 4699 11942 4711 11994
rect 4711 11942 4741 11994
rect 4765 11942 4775 11994
rect 4775 11942 4821 11994
rect 4525 11940 4581 11942
rect 4605 11940 4661 11942
rect 4685 11940 4741 11942
rect 4765 11940 4821 11942
rect 1214 11620 1270 11656
rect 1214 11600 1216 11620
rect 1216 11600 1268 11620
rect 1268 11600 1270 11620
rect 3865 11450 3921 11452
rect 3945 11450 4001 11452
rect 4025 11450 4081 11452
rect 4105 11450 4161 11452
rect 3865 11398 3911 11450
rect 3911 11398 3921 11450
rect 3945 11398 3975 11450
rect 3975 11398 3987 11450
rect 3987 11398 4001 11450
rect 4025 11398 4039 11450
rect 4039 11398 4051 11450
rect 4051 11398 4081 11450
rect 4105 11398 4115 11450
rect 4115 11398 4161 11450
rect 3865 11396 3921 11398
rect 3945 11396 4001 11398
rect 4025 11396 4081 11398
rect 4105 11396 4161 11398
rect 2318 10920 2374 10976
rect 4525 10906 4581 10908
rect 4605 10906 4661 10908
rect 4685 10906 4741 10908
rect 4765 10906 4821 10908
rect 4525 10854 4571 10906
rect 4571 10854 4581 10906
rect 4605 10854 4635 10906
rect 4635 10854 4647 10906
rect 4647 10854 4661 10906
rect 4685 10854 4699 10906
rect 4699 10854 4711 10906
rect 4711 10854 4741 10906
rect 4765 10854 4775 10906
rect 4775 10854 4821 10906
rect 4525 10852 4581 10854
rect 4605 10852 4661 10854
rect 4685 10852 4741 10854
rect 4765 10852 4821 10854
rect 7844 11450 7900 11452
rect 7924 11450 7980 11452
rect 8004 11450 8060 11452
rect 8084 11450 8140 11452
rect 7844 11398 7890 11450
rect 7890 11398 7900 11450
rect 7924 11398 7954 11450
rect 7954 11398 7966 11450
rect 7966 11398 7980 11450
rect 8004 11398 8018 11450
rect 8018 11398 8030 11450
rect 8030 11398 8060 11450
rect 8084 11398 8094 11450
rect 8094 11398 8140 11450
rect 7844 11396 7900 11398
rect 7924 11396 7980 11398
rect 8004 11396 8060 11398
rect 8084 11396 8140 11398
rect 8504 11994 8560 11996
rect 8584 11994 8640 11996
rect 8664 11994 8720 11996
rect 8744 11994 8800 11996
rect 8504 11942 8550 11994
rect 8550 11942 8560 11994
rect 8584 11942 8614 11994
rect 8614 11942 8626 11994
rect 8626 11942 8640 11994
rect 8664 11942 8678 11994
rect 8678 11942 8690 11994
rect 8690 11942 8720 11994
rect 8744 11942 8754 11994
rect 8754 11942 8800 11994
rect 8504 11940 8560 11942
rect 8584 11940 8640 11942
rect 8664 11940 8720 11942
rect 8744 11940 8800 11942
rect 3865 10362 3921 10364
rect 3945 10362 4001 10364
rect 4025 10362 4081 10364
rect 4105 10362 4161 10364
rect 3865 10310 3911 10362
rect 3911 10310 3921 10362
rect 3945 10310 3975 10362
rect 3975 10310 3987 10362
rect 3987 10310 4001 10362
rect 4025 10310 4039 10362
rect 4039 10310 4051 10362
rect 4051 10310 4081 10362
rect 4105 10310 4115 10362
rect 4115 10310 4161 10362
rect 3865 10308 3921 10310
rect 3945 10308 4001 10310
rect 4025 10308 4081 10310
rect 4105 10308 4161 10310
rect 1122 10240 1178 10296
rect 4525 9818 4581 9820
rect 4605 9818 4661 9820
rect 4685 9818 4741 9820
rect 4765 9818 4821 9820
rect 4525 9766 4571 9818
rect 4571 9766 4581 9818
rect 4605 9766 4635 9818
rect 4635 9766 4647 9818
rect 4647 9766 4661 9818
rect 4685 9766 4699 9818
rect 4699 9766 4711 9818
rect 4711 9766 4741 9818
rect 4765 9766 4775 9818
rect 4775 9766 4821 9818
rect 4525 9764 4581 9766
rect 4605 9764 4661 9766
rect 4685 9764 4741 9766
rect 4765 9764 4821 9766
rect 3865 9274 3921 9276
rect 3945 9274 4001 9276
rect 4025 9274 4081 9276
rect 4105 9274 4161 9276
rect 3865 9222 3911 9274
rect 3911 9222 3921 9274
rect 3945 9222 3975 9274
rect 3975 9222 3987 9274
rect 3987 9222 4001 9274
rect 4025 9222 4039 9274
rect 4039 9222 4051 9274
rect 4051 9222 4081 9274
rect 4105 9222 4115 9274
rect 4115 9222 4161 9274
rect 3865 9220 3921 9222
rect 3945 9220 4001 9222
rect 4025 9220 4081 9222
rect 4105 9220 4161 9222
rect 1214 8900 1270 8936
rect 1214 8880 1216 8900
rect 1216 8880 1268 8900
rect 1268 8880 1270 8900
rect 4525 8730 4581 8732
rect 4605 8730 4661 8732
rect 4685 8730 4741 8732
rect 4765 8730 4821 8732
rect 4525 8678 4571 8730
rect 4571 8678 4581 8730
rect 4605 8678 4635 8730
rect 4635 8678 4647 8730
rect 4647 8678 4661 8730
rect 4685 8678 4699 8730
rect 4699 8678 4711 8730
rect 4711 8678 4741 8730
rect 4765 8678 4775 8730
rect 4775 8678 4821 8730
rect 4525 8676 4581 8678
rect 4605 8676 4661 8678
rect 4685 8676 4741 8678
rect 4765 8676 4821 8678
rect 3865 8186 3921 8188
rect 3945 8186 4001 8188
rect 4025 8186 4081 8188
rect 4105 8186 4161 8188
rect 3865 8134 3911 8186
rect 3911 8134 3921 8186
rect 3945 8134 3975 8186
rect 3975 8134 3987 8186
rect 3987 8134 4001 8186
rect 4025 8134 4039 8186
rect 4039 8134 4051 8186
rect 4051 8134 4081 8186
rect 4105 8134 4115 8186
rect 4115 8134 4161 8186
rect 3865 8132 3921 8134
rect 3945 8132 4001 8134
rect 4025 8132 4081 8134
rect 4105 8132 4161 8134
rect 4525 7642 4581 7644
rect 4605 7642 4661 7644
rect 4685 7642 4741 7644
rect 4765 7642 4821 7644
rect 4525 7590 4571 7642
rect 4571 7590 4581 7642
rect 4605 7590 4635 7642
rect 4635 7590 4647 7642
rect 4647 7590 4661 7642
rect 4685 7590 4699 7642
rect 4699 7590 4711 7642
rect 4711 7590 4741 7642
rect 4765 7590 4775 7642
rect 4775 7590 4821 7642
rect 4525 7588 4581 7590
rect 4605 7588 4661 7590
rect 4685 7588 4741 7590
rect 4765 7588 4821 7590
rect 3865 7098 3921 7100
rect 3945 7098 4001 7100
rect 4025 7098 4081 7100
rect 4105 7098 4161 7100
rect 3865 7046 3911 7098
rect 3911 7046 3921 7098
rect 3945 7046 3975 7098
rect 3975 7046 3987 7098
rect 3987 7046 4001 7098
rect 4025 7046 4039 7098
rect 4039 7046 4051 7098
rect 4051 7046 4081 7098
rect 4105 7046 4115 7098
rect 4115 7046 4161 7098
rect 3865 7044 3921 7046
rect 3945 7044 4001 7046
rect 4025 7044 4081 7046
rect 4105 7044 4161 7046
rect 8504 10906 8560 10908
rect 8584 10906 8640 10908
rect 8664 10906 8720 10908
rect 8744 10906 8800 10908
rect 8504 10854 8550 10906
rect 8550 10854 8560 10906
rect 8584 10854 8614 10906
rect 8614 10854 8626 10906
rect 8626 10854 8640 10906
rect 8664 10854 8678 10906
rect 8678 10854 8690 10906
rect 8690 10854 8720 10906
rect 8744 10854 8754 10906
rect 8754 10854 8800 10906
rect 8504 10852 8560 10854
rect 8584 10852 8640 10854
rect 8664 10852 8720 10854
rect 8744 10852 8800 10854
rect 7844 10362 7900 10364
rect 7924 10362 7980 10364
rect 8004 10362 8060 10364
rect 8084 10362 8140 10364
rect 7844 10310 7890 10362
rect 7890 10310 7900 10362
rect 7924 10310 7954 10362
rect 7954 10310 7966 10362
rect 7966 10310 7980 10362
rect 8004 10310 8018 10362
rect 8018 10310 8030 10362
rect 8030 10310 8060 10362
rect 8084 10310 8094 10362
rect 8094 10310 8140 10362
rect 7844 10308 7900 10310
rect 7924 10308 7980 10310
rect 8004 10308 8060 10310
rect 8084 10308 8140 10310
rect 11823 17978 11879 17980
rect 11903 17978 11959 17980
rect 11983 17978 12039 17980
rect 12063 17978 12119 17980
rect 11823 17926 11869 17978
rect 11869 17926 11879 17978
rect 11903 17926 11933 17978
rect 11933 17926 11945 17978
rect 11945 17926 11959 17978
rect 11983 17926 11997 17978
rect 11997 17926 12009 17978
rect 12009 17926 12039 17978
rect 12063 17926 12073 17978
rect 12073 17926 12119 17978
rect 11823 17924 11879 17926
rect 11903 17924 11959 17926
rect 11983 17924 12039 17926
rect 12063 17924 12119 17926
rect 15802 17978 15858 17980
rect 15882 17978 15938 17980
rect 15962 17978 16018 17980
rect 16042 17978 16098 17980
rect 15802 17926 15848 17978
rect 15848 17926 15858 17978
rect 15882 17926 15912 17978
rect 15912 17926 15924 17978
rect 15924 17926 15938 17978
rect 15962 17926 15976 17978
rect 15976 17926 15988 17978
rect 15988 17926 16018 17978
rect 16042 17926 16052 17978
rect 16052 17926 16098 17978
rect 15802 17924 15858 17926
rect 15882 17924 15938 17926
rect 15962 17924 16018 17926
rect 16042 17924 16098 17926
rect 8504 9818 8560 9820
rect 8584 9818 8640 9820
rect 8664 9818 8720 9820
rect 8744 9818 8800 9820
rect 8504 9766 8550 9818
rect 8550 9766 8560 9818
rect 8584 9766 8614 9818
rect 8614 9766 8626 9818
rect 8626 9766 8640 9818
rect 8664 9766 8678 9818
rect 8678 9766 8690 9818
rect 8690 9766 8720 9818
rect 8744 9766 8754 9818
rect 8754 9766 8800 9818
rect 8504 9764 8560 9766
rect 8584 9764 8640 9766
rect 8664 9764 8720 9766
rect 8744 9764 8800 9766
rect 7844 9274 7900 9276
rect 7924 9274 7980 9276
rect 8004 9274 8060 9276
rect 8084 9274 8140 9276
rect 7844 9222 7890 9274
rect 7890 9222 7900 9274
rect 7924 9222 7954 9274
rect 7954 9222 7966 9274
rect 7966 9222 7980 9274
rect 8004 9222 8018 9274
rect 8018 9222 8030 9274
rect 8030 9222 8060 9274
rect 8084 9222 8094 9274
rect 8094 9222 8140 9274
rect 7844 9220 7900 9222
rect 7924 9220 7980 9222
rect 8004 9220 8060 9222
rect 8084 9220 8140 9222
rect 12483 17434 12539 17436
rect 12563 17434 12619 17436
rect 12643 17434 12699 17436
rect 12723 17434 12779 17436
rect 12483 17382 12529 17434
rect 12529 17382 12539 17434
rect 12563 17382 12593 17434
rect 12593 17382 12605 17434
rect 12605 17382 12619 17434
rect 12643 17382 12657 17434
rect 12657 17382 12669 17434
rect 12669 17382 12699 17434
rect 12723 17382 12733 17434
rect 12733 17382 12779 17434
rect 12483 17380 12539 17382
rect 12563 17380 12619 17382
rect 12643 17380 12699 17382
rect 12723 17380 12779 17382
rect 11823 16890 11879 16892
rect 11903 16890 11959 16892
rect 11983 16890 12039 16892
rect 12063 16890 12119 16892
rect 11823 16838 11869 16890
rect 11869 16838 11879 16890
rect 11903 16838 11933 16890
rect 11933 16838 11945 16890
rect 11945 16838 11959 16890
rect 11983 16838 11997 16890
rect 11997 16838 12009 16890
rect 12009 16838 12039 16890
rect 12063 16838 12073 16890
rect 12073 16838 12119 16890
rect 11823 16836 11879 16838
rect 11903 16836 11959 16838
rect 11983 16836 12039 16838
rect 12063 16836 12119 16838
rect 12483 16346 12539 16348
rect 12563 16346 12619 16348
rect 12643 16346 12699 16348
rect 12723 16346 12779 16348
rect 12483 16294 12529 16346
rect 12529 16294 12539 16346
rect 12563 16294 12593 16346
rect 12593 16294 12605 16346
rect 12605 16294 12619 16346
rect 12643 16294 12657 16346
rect 12657 16294 12669 16346
rect 12669 16294 12699 16346
rect 12723 16294 12733 16346
rect 12733 16294 12779 16346
rect 12483 16292 12539 16294
rect 12563 16292 12619 16294
rect 12643 16292 12699 16294
rect 12723 16292 12779 16294
rect 11823 15802 11879 15804
rect 11903 15802 11959 15804
rect 11983 15802 12039 15804
rect 12063 15802 12119 15804
rect 11823 15750 11869 15802
rect 11869 15750 11879 15802
rect 11903 15750 11933 15802
rect 11933 15750 11945 15802
rect 11945 15750 11959 15802
rect 11983 15750 11997 15802
rect 11997 15750 12009 15802
rect 12009 15750 12039 15802
rect 12063 15750 12073 15802
rect 12073 15750 12119 15802
rect 11823 15748 11879 15750
rect 11903 15748 11959 15750
rect 11983 15748 12039 15750
rect 12063 15748 12119 15750
rect 12483 15258 12539 15260
rect 12563 15258 12619 15260
rect 12643 15258 12699 15260
rect 12723 15258 12779 15260
rect 12483 15206 12529 15258
rect 12529 15206 12539 15258
rect 12563 15206 12593 15258
rect 12593 15206 12605 15258
rect 12605 15206 12619 15258
rect 12643 15206 12657 15258
rect 12657 15206 12669 15258
rect 12669 15206 12699 15258
rect 12723 15206 12733 15258
rect 12733 15206 12779 15258
rect 12483 15204 12539 15206
rect 12563 15204 12619 15206
rect 12643 15204 12699 15206
rect 12723 15204 12779 15206
rect 11823 14714 11879 14716
rect 11903 14714 11959 14716
rect 11983 14714 12039 14716
rect 12063 14714 12119 14716
rect 11823 14662 11869 14714
rect 11869 14662 11879 14714
rect 11903 14662 11933 14714
rect 11933 14662 11945 14714
rect 11945 14662 11959 14714
rect 11983 14662 11997 14714
rect 11997 14662 12009 14714
rect 12009 14662 12039 14714
rect 12063 14662 12073 14714
rect 12073 14662 12119 14714
rect 11823 14660 11879 14662
rect 11903 14660 11959 14662
rect 11983 14660 12039 14662
rect 12063 14660 12119 14662
rect 12483 14170 12539 14172
rect 12563 14170 12619 14172
rect 12643 14170 12699 14172
rect 12723 14170 12779 14172
rect 12483 14118 12529 14170
rect 12529 14118 12539 14170
rect 12563 14118 12593 14170
rect 12593 14118 12605 14170
rect 12605 14118 12619 14170
rect 12643 14118 12657 14170
rect 12657 14118 12669 14170
rect 12669 14118 12699 14170
rect 12723 14118 12733 14170
rect 12733 14118 12779 14170
rect 12483 14116 12539 14118
rect 12563 14116 12619 14118
rect 12643 14116 12699 14118
rect 12723 14116 12779 14118
rect 11823 13626 11879 13628
rect 11903 13626 11959 13628
rect 11983 13626 12039 13628
rect 12063 13626 12119 13628
rect 11823 13574 11869 13626
rect 11869 13574 11879 13626
rect 11903 13574 11933 13626
rect 11933 13574 11945 13626
rect 11945 13574 11959 13626
rect 11983 13574 11997 13626
rect 11997 13574 12009 13626
rect 12009 13574 12039 13626
rect 12063 13574 12073 13626
rect 12073 13574 12119 13626
rect 11823 13572 11879 13574
rect 11903 13572 11959 13574
rect 11983 13572 12039 13574
rect 12063 13572 12119 13574
rect 11823 12538 11879 12540
rect 11903 12538 11959 12540
rect 11983 12538 12039 12540
rect 12063 12538 12119 12540
rect 11823 12486 11869 12538
rect 11869 12486 11879 12538
rect 11903 12486 11933 12538
rect 11933 12486 11945 12538
rect 11945 12486 11959 12538
rect 11983 12486 11997 12538
rect 11997 12486 12009 12538
rect 12009 12486 12039 12538
rect 12063 12486 12073 12538
rect 12073 12486 12119 12538
rect 11823 12484 11879 12486
rect 11903 12484 11959 12486
rect 11983 12484 12039 12486
rect 12063 12484 12119 12486
rect 12483 13082 12539 13084
rect 12563 13082 12619 13084
rect 12643 13082 12699 13084
rect 12723 13082 12779 13084
rect 12483 13030 12529 13082
rect 12529 13030 12539 13082
rect 12563 13030 12593 13082
rect 12593 13030 12605 13082
rect 12605 13030 12619 13082
rect 12643 13030 12657 13082
rect 12657 13030 12669 13082
rect 12669 13030 12699 13082
rect 12723 13030 12733 13082
rect 12733 13030 12779 13082
rect 12483 13028 12539 13030
rect 12563 13028 12619 13030
rect 12643 13028 12699 13030
rect 12723 13028 12779 13030
rect 16462 17434 16518 17436
rect 16542 17434 16598 17436
rect 16622 17434 16678 17436
rect 16702 17434 16758 17436
rect 16462 17382 16508 17434
rect 16508 17382 16518 17434
rect 16542 17382 16572 17434
rect 16572 17382 16584 17434
rect 16584 17382 16598 17434
rect 16622 17382 16636 17434
rect 16636 17382 16648 17434
rect 16648 17382 16678 17434
rect 16702 17382 16712 17434
rect 16712 17382 16758 17434
rect 16462 17380 16518 17382
rect 16542 17380 16598 17382
rect 16622 17380 16678 17382
rect 16702 17380 16758 17382
rect 15802 16890 15858 16892
rect 15882 16890 15938 16892
rect 15962 16890 16018 16892
rect 16042 16890 16098 16892
rect 15802 16838 15848 16890
rect 15848 16838 15858 16890
rect 15882 16838 15912 16890
rect 15912 16838 15924 16890
rect 15924 16838 15938 16890
rect 15962 16838 15976 16890
rect 15976 16838 15988 16890
rect 15988 16838 16018 16890
rect 16042 16838 16052 16890
rect 16052 16838 16098 16890
rect 15802 16836 15858 16838
rect 15882 16836 15938 16838
rect 15962 16836 16018 16838
rect 16042 16836 16098 16838
rect 16462 16346 16518 16348
rect 16542 16346 16598 16348
rect 16622 16346 16678 16348
rect 16702 16346 16758 16348
rect 16462 16294 16508 16346
rect 16508 16294 16518 16346
rect 16542 16294 16572 16346
rect 16572 16294 16584 16346
rect 16584 16294 16598 16346
rect 16622 16294 16636 16346
rect 16636 16294 16648 16346
rect 16648 16294 16678 16346
rect 16702 16294 16712 16346
rect 16712 16294 16758 16346
rect 16462 16292 16518 16294
rect 16542 16292 16598 16294
rect 16622 16292 16678 16294
rect 16702 16292 16758 16294
rect 15802 15802 15858 15804
rect 15882 15802 15938 15804
rect 15962 15802 16018 15804
rect 16042 15802 16098 15804
rect 15802 15750 15848 15802
rect 15848 15750 15858 15802
rect 15882 15750 15912 15802
rect 15912 15750 15924 15802
rect 15924 15750 15938 15802
rect 15962 15750 15976 15802
rect 15976 15750 15988 15802
rect 15988 15750 16018 15802
rect 16042 15750 16052 15802
rect 16052 15750 16098 15802
rect 15802 15748 15858 15750
rect 15882 15748 15938 15750
rect 15962 15748 16018 15750
rect 16042 15748 16098 15750
rect 16462 15258 16518 15260
rect 16542 15258 16598 15260
rect 16622 15258 16678 15260
rect 16702 15258 16758 15260
rect 16462 15206 16508 15258
rect 16508 15206 16518 15258
rect 16542 15206 16572 15258
rect 16572 15206 16584 15258
rect 16584 15206 16598 15258
rect 16622 15206 16636 15258
rect 16636 15206 16648 15258
rect 16648 15206 16678 15258
rect 16702 15206 16712 15258
rect 16712 15206 16758 15258
rect 16462 15204 16518 15206
rect 16542 15204 16598 15206
rect 16622 15204 16678 15206
rect 16702 15204 16758 15206
rect 15802 14714 15858 14716
rect 15882 14714 15938 14716
rect 15962 14714 16018 14716
rect 16042 14714 16098 14716
rect 15802 14662 15848 14714
rect 15848 14662 15858 14714
rect 15882 14662 15912 14714
rect 15912 14662 15924 14714
rect 15924 14662 15938 14714
rect 15962 14662 15976 14714
rect 15976 14662 15988 14714
rect 15988 14662 16018 14714
rect 16042 14662 16052 14714
rect 16052 14662 16098 14714
rect 15802 14660 15858 14662
rect 15882 14660 15938 14662
rect 15962 14660 16018 14662
rect 16042 14660 16098 14662
rect 16462 14170 16518 14172
rect 16542 14170 16598 14172
rect 16622 14170 16678 14172
rect 16702 14170 16758 14172
rect 16462 14118 16508 14170
rect 16508 14118 16518 14170
rect 16542 14118 16572 14170
rect 16572 14118 16584 14170
rect 16584 14118 16598 14170
rect 16622 14118 16636 14170
rect 16636 14118 16648 14170
rect 16648 14118 16678 14170
rect 16702 14118 16712 14170
rect 16712 14118 16758 14170
rect 16462 14116 16518 14118
rect 16542 14116 16598 14118
rect 16622 14116 16678 14118
rect 16702 14116 16758 14118
rect 12483 11994 12539 11996
rect 12563 11994 12619 11996
rect 12643 11994 12699 11996
rect 12723 11994 12779 11996
rect 12483 11942 12529 11994
rect 12529 11942 12539 11994
rect 12563 11942 12593 11994
rect 12593 11942 12605 11994
rect 12605 11942 12619 11994
rect 12643 11942 12657 11994
rect 12657 11942 12669 11994
rect 12669 11942 12699 11994
rect 12723 11942 12733 11994
rect 12733 11942 12779 11994
rect 12483 11940 12539 11942
rect 12563 11940 12619 11942
rect 12643 11940 12699 11942
rect 12723 11940 12779 11942
rect 8504 8730 8560 8732
rect 8584 8730 8640 8732
rect 8664 8730 8720 8732
rect 8744 8730 8800 8732
rect 8504 8678 8550 8730
rect 8550 8678 8560 8730
rect 8584 8678 8614 8730
rect 8614 8678 8626 8730
rect 8626 8678 8640 8730
rect 8664 8678 8678 8730
rect 8678 8678 8690 8730
rect 8690 8678 8720 8730
rect 8744 8678 8754 8730
rect 8754 8678 8800 8730
rect 8504 8676 8560 8678
rect 8584 8676 8640 8678
rect 8664 8676 8720 8678
rect 8744 8676 8800 8678
rect 7844 8186 7900 8188
rect 7924 8186 7980 8188
rect 8004 8186 8060 8188
rect 8084 8186 8140 8188
rect 7844 8134 7890 8186
rect 7890 8134 7900 8186
rect 7924 8134 7954 8186
rect 7954 8134 7966 8186
rect 7966 8134 7980 8186
rect 8004 8134 8018 8186
rect 8018 8134 8030 8186
rect 8030 8134 8060 8186
rect 8084 8134 8094 8186
rect 8094 8134 8140 8186
rect 7844 8132 7900 8134
rect 7924 8132 7980 8134
rect 8004 8132 8060 8134
rect 8084 8132 8140 8134
rect 7844 7098 7900 7100
rect 7924 7098 7980 7100
rect 8004 7098 8060 7100
rect 8084 7098 8140 7100
rect 7844 7046 7890 7098
rect 7890 7046 7900 7098
rect 7924 7046 7954 7098
rect 7954 7046 7966 7098
rect 7966 7046 7980 7098
rect 8004 7046 8018 7098
rect 8018 7046 8030 7098
rect 8030 7046 8060 7098
rect 8084 7046 8094 7098
rect 8094 7046 8140 7098
rect 7844 7044 7900 7046
rect 7924 7044 7980 7046
rect 8004 7044 8060 7046
rect 8084 7044 8140 7046
rect 4525 6554 4581 6556
rect 4605 6554 4661 6556
rect 4685 6554 4741 6556
rect 4765 6554 4821 6556
rect 4525 6502 4571 6554
rect 4571 6502 4581 6554
rect 4605 6502 4635 6554
rect 4635 6502 4647 6554
rect 4647 6502 4661 6554
rect 4685 6502 4699 6554
rect 4699 6502 4711 6554
rect 4711 6502 4741 6554
rect 4765 6502 4775 6554
rect 4775 6502 4821 6554
rect 4525 6500 4581 6502
rect 4605 6500 4661 6502
rect 4685 6500 4741 6502
rect 4765 6500 4821 6502
rect 3865 6010 3921 6012
rect 3945 6010 4001 6012
rect 4025 6010 4081 6012
rect 4105 6010 4161 6012
rect 3865 5958 3911 6010
rect 3911 5958 3921 6010
rect 3945 5958 3975 6010
rect 3975 5958 3987 6010
rect 3987 5958 4001 6010
rect 4025 5958 4039 6010
rect 4039 5958 4051 6010
rect 4051 5958 4081 6010
rect 4105 5958 4115 6010
rect 4115 5958 4161 6010
rect 3865 5956 3921 5958
rect 3945 5956 4001 5958
rect 4025 5956 4081 5958
rect 4105 5956 4161 5958
rect 4525 5466 4581 5468
rect 4605 5466 4661 5468
rect 4685 5466 4741 5468
rect 4765 5466 4821 5468
rect 4525 5414 4571 5466
rect 4571 5414 4581 5466
rect 4605 5414 4635 5466
rect 4635 5414 4647 5466
rect 4647 5414 4661 5466
rect 4685 5414 4699 5466
rect 4699 5414 4711 5466
rect 4711 5414 4741 5466
rect 4765 5414 4775 5466
rect 4775 5414 4821 5466
rect 4525 5412 4581 5414
rect 4605 5412 4661 5414
rect 4685 5412 4741 5414
rect 4765 5412 4821 5414
rect 3865 4922 3921 4924
rect 3945 4922 4001 4924
rect 4025 4922 4081 4924
rect 4105 4922 4161 4924
rect 3865 4870 3911 4922
rect 3911 4870 3921 4922
rect 3945 4870 3975 4922
rect 3975 4870 3987 4922
rect 3987 4870 4001 4922
rect 4025 4870 4039 4922
rect 4039 4870 4051 4922
rect 4051 4870 4081 4922
rect 4105 4870 4115 4922
rect 4115 4870 4161 4922
rect 3865 4868 3921 4870
rect 3945 4868 4001 4870
rect 4025 4868 4081 4870
rect 4105 4868 4161 4870
rect 4525 4378 4581 4380
rect 4605 4378 4661 4380
rect 4685 4378 4741 4380
rect 4765 4378 4821 4380
rect 4525 4326 4571 4378
rect 4571 4326 4581 4378
rect 4605 4326 4635 4378
rect 4635 4326 4647 4378
rect 4647 4326 4661 4378
rect 4685 4326 4699 4378
rect 4699 4326 4711 4378
rect 4711 4326 4741 4378
rect 4765 4326 4775 4378
rect 4775 4326 4821 4378
rect 4525 4324 4581 4326
rect 4605 4324 4661 4326
rect 4685 4324 4741 4326
rect 4765 4324 4821 4326
rect 3865 3834 3921 3836
rect 3945 3834 4001 3836
rect 4025 3834 4081 3836
rect 4105 3834 4161 3836
rect 3865 3782 3911 3834
rect 3911 3782 3921 3834
rect 3945 3782 3975 3834
rect 3975 3782 3987 3834
rect 3987 3782 4001 3834
rect 4025 3782 4039 3834
rect 4039 3782 4051 3834
rect 4051 3782 4081 3834
rect 4105 3782 4115 3834
rect 4115 3782 4161 3834
rect 3865 3780 3921 3782
rect 3945 3780 4001 3782
rect 4025 3780 4081 3782
rect 4105 3780 4161 3782
rect 4525 3290 4581 3292
rect 4605 3290 4661 3292
rect 4685 3290 4741 3292
rect 4765 3290 4821 3292
rect 4525 3238 4571 3290
rect 4571 3238 4581 3290
rect 4605 3238 4635 3290
rect 4635 3238 4647 3290
rect 4647 3238 4661 3290
rect 4685 3238 4699 3290
rect 4699 3238 4711 3290
rect 4711 3238 4741 3290
rect 4765 3238 4775 3290
rect 4775 3238 4821 3290
rect 4525 3236 4581 3238
rect 4605 3236 4661 3238
rect 4685 3236 4741 3238
rect 4765 3236 4821 3238
rect 3865 2746 3921 2748
rect 3945 2746 4001 2748
rect 4025 2746 4081 2748
rect 4105 2746 4161 2748
rect 3865 2694 3911 2746
rect 3911 2694 3921 2746
rect 3945 2694 3975 2746
rect 3975 2694 3987 2746
rect 3987 2694 4001 2746
rect 4025 2694 4039 2746
rect 4039 2694 4051 2746
rect 4051 2694 4081 2746
rect 4105 2694 4115 2746
rect 4115 2694 4161 2746
rect 3865 2692 3921 2694
rect 3945 2692 4001 2694
rect 4025 2692 4081 2694
rect 4105 2692 4161 2694
rect 11823 11450 11879 11452
rect 11903 11450 11959 11452
rect 11983 11450 12039 11452
rect 12063 11450 12119 11452
rect 11823 11398 11869 11450
rect 11869 11398 11879 11450
rect 11903 11398 11933 11450
rect 11933 11398 11945 11450
rect 11945 11398 11959 11450
rect 11983 11398 11997 11450
rect 11997 11398 12009 11450
rect 12009 11398 12039 11450
rect 12063 11398 12073 11450
rect 12073 11398 12119 11450
rect 11823 11396 11879 11398
rect 11903 11396 11959 11398
rect 11983 11396 12039 11398
rect 12063 11396 12119 11398
rect 11823 10362 11879 10364
rect 11903 10362 11959 10364
rect 11983 10362 12039 10364
rect 12063 10362 12119 10364
rect 11823 10310 11869 10362
rect 11869 10310 11879 10362
rect 11903 10310 11933 10362
rect 11933 10310 11945 10362
rect 11945 10310 11959 10362
rect 11983 10310 11997 10362
rect 11997 10310 12009 10362
rect 12009 10310 12039 10362
rect 12063 10310 12073 10362
rect 12073 10310 12119 10362
rect 11823 10308 11879 10310
rect 11903 10308 11959 10310
rect 11983 10308 12039 10310
rect 12063 10308 12119 10310
rect 8504 7642 8560 7644
rect 8584 7642 8640 7644
rect 8664 7642 8720 7644
rect 8744 7642 8800 7644
rect 8504 7590 8550 7642
rect 8550 7590 8560 7642
rect 8584 7590 8614 7642
rect 8614 7590 8626 7642
rect 8626 7590 8640 7642
rect 8664 7590 8678 7642
rect 8678 7590 8690 7642
rect 8690 7590 8720 7642
rect 8744 7590 8754 7642
rect 8754 7590 8800 7642
rect 8504 7588 8560 7590
rect 8584 7588 8640 7590
rect 8664 7588 8720 7590
rect 8744 7588 8800 7590
rect 8504 6554 8560 6556
rect 8584 6554 8640 6556
rect 8664 6554 8720 6556
rect 8744 6554 8800 6556
rect 8504 6502 8550 6554
rect 8550 6502 8560 6554
rect 8584 6502 8614 6554
rect 8614 6502 8626 6554
rect 8626 6502 8640 6554
rect 8664 6502 8678 6554
rect 8678 6502 8690 6554
rect 8690 6502 8720 6554
rect 8744 6502 8754 6554
rect 8754 6502 8800 6554
rect 8504 6500 8560 6502
rect 8584 6500 8640 6502
rect 8664 6500 8720 6502
rect 8744 6500 8800 6502
rect 7844 6010 7900 6012
rect 7924 6010 7980 6012
rect 8004 6010 8060 6012
rect 8084 6010 8140 6012
rect 7844 5958 7890 6010
rect 7890 5958 7900 6010
rect 7924 5958 7954 6010
rect 7954 5958 7966 6010
rect 7966 5958 7980 6010
rect 8004 5958 8018 6010
rect 8018 5958 8030 6010
rect 8030 5958 8060 6010
rect 8084 5958 8094 6010
rect 8094 5958 8140 6010
rect 7844 5956 7900 5958
rect 7924 5956 7980 5958
rect 8004 5956 8060 5958
rect 8084 5956 8140 5958
rect 8504 5466 8560 5468
rect 8584 5466 8640 5468
rect 8664 5466 8720 5468
rect 8744 5466 8800 5468
rect 8504 5414 8550 5466
rect 8550 5414 8560 5466
rect 8584 5414 8614 5466
rect 8614 5414 8626 5466
rect 8626 5414 8640 5466
rect 8664 5414 8678 5466
rect 8678 5414 8690 5466
rect 8690 5414 8720 5466
rect 8744 5414 8754 5466
rect 8754 5414 8800 5466
rect 8504 5412 8560 5414
rect 8584 5412 8640 5414
rect 8664 5412 8720 5414
rect 8744 5412 8800 5414
rect 7844 4922 7900 4924
rect 7924 4922 7980 4924
rect 8004 4922 8060 4924
rect 8084 4922 8140 4924
rect 7844 4870 7890 4922
rect 7890 4870 7900 4922
rect 7924 4870 7954 4922
rect 7954 4870 7966 4922
rect 7966 4870 7980 4922
rect 8004 4870 8018 4922
rect 8018 4870 8030 4922
rect 8030 4870 8060 4922
rect 8084 4870 8094 4922
rect 8094 4870 8140 4922
rect 7844 4868 7900 4870
rect 7924 4868 7980 4870
rect 8004 4868 8060 4870
rect 8084 4868 8140 4870
rect 8504 4378 8560 4380
rect 8584 4378 8640 4380
rect 8664 4378 8720 4380
rect 8744 4378 8800 4380
rect 8504 4326 8550 4378
rect 8550 4326 8560 4378
rect 8584 4326 8614 4378
rect 8614 4326 8626 4378
rect 8626 4326 8640 4378
rect 8664 4326 8678 4378
rect 8678 4326 8690 4378
rect 8690 4326 8720 4378
rect 8744 4326 8754 4378
rect 8754 4326 8800 4378
rect 8504 4324 8560 4326
rect 8584 4324 8640 4326
rect 8664 4324 8720 4326
rect 8744 4324 8800 4326
rect 7844 3834 7900 3836
rect 7924 3834 7980 3836
rect 8004 3834 8060 3836
rect 8084 3834 8140 3836
rect 7844 3782 7890 3834
rect 7890 3782 7900 3834
rect 7924 3782 7954 3834
rect 7954 3782 7966 3834
rect 7966 3782 7980 3834
rect 8004 3782 8018 3834
rect 8018 3782 8030 3834
rect 8030 3782 8060 3834
rect 8084 3782 8094 3834
rect 8094 3782 8140 3834
rect 7844 3780 7900 3782
rect 7924 3780 7980 3782
rect 8004 3780 8060 3782
rect 8084 3780 8140 3782
rect 8504 3290 8560 3292
rect 8584 3290 8640 3292
rect 8664 3290 8720 3292
rect 8744 3290 8800 3292
rect 8504 3238 8550 3290
rect 8550 3238 8560 3290
rect 8584 3238 8614 3290
rect 8614 3238 8626 3290
rect 8626 3238 8640 3290
rect 8664 3238 8678 3290
rect 8678 3238 8690 3290
rect 8690 3238 8720 3290
rect 8744 3238 8754 3290
rect 8754 3238 8800 3290
rect 8504 3236 8560 3238
rect 8584 3236 8640 3238
rect 8664 3236 8720 3238
rect 8744 3236 8800 3238
rect 7844 2746 7900 2748
rect 7924 2746 7980 2748
rect 8004 2746 8060 2748
rect 8084 2746 8140 2748
rect 7844 2694 7890 2746
rect 7890 2694 7900 2746
rect 7924 2694 7954 2746
rect 7954 2694 7966 2746
rect 7966 2694 7980 2746
rect 8004 2694 8018 2746
rect 8018 2694 8030 2746
rect 8030 2694 8060 2746
rect 8084 2694 8094 2746
rect 8094 2694 8140 2746
rect 7844 2692 7900 2694
rect 7924 2692 7980 2694
rect 8004 2692 8060 2694
rect 8084 2692 8140 2694
rect 11823 9274 11879 9276
rect 11903 9274 11959 9276
rect 11983 9274 12039 9276
rect 12063 9274 12119 9276
rect 11823 9222 11869 9274
rect 11869 9222 11879 9274
rect 11903 9222 11933 9274
rect 11933 9222 11945 9274
rect 11945 9222 11959 9274
rect 11983 9222 11997 9274
rect 11997 9222 12009 9274
rect 12009 9222 12039 9274
rect 12063 9222 12073 9274
rect 12073 9222 12119 9274
rect 11823 9220 11879 9222
rect 11903 9220 11959 9222
rect 11983 9220 12039 9222
rect 12063 9220 12119 9222
rect 4525 2202 4581 2204
rect 4605 2202 4661 2204
rect 4685 2202 4741 2204
rect 4765 2202 4821 2204
rect 4525 2150 4571 2202
rect 4571 2150 4581 2202
rect 4605 2150 4635 2202
rect 4635 2150 4647 2202
rect 4647 2150 4661 2202
rect 4685 2150 4699 2202
rect 4699 2150 4711 2202
rect 4711 2150 4741 2202
rect 4765 2150 4775 2202
rect 4775 2150 4821 2202
rect 4525 2148 4581 2150
rect 4605 2148 4661 2150
rect 4685 2148 4741 2150
rect 4765 2148 4821 2150
rect 8504 2202 8560 2204
rect 8584 2202 8640 2204
rect 8664 2202 8720 2204
rect 8744 2202 8800 2204
rect 8504 2150 8550 2202
rect 8550 2150 8560 2202
rect 8584 2150 8614 2202
rect 8614 2150 8626 2202
rect 8626 2150 8640 2202
rect 8664 2150 8678 2202
rect 8678 2150 8690 2202
rect 8690 2150 8720 2202
rect 8744 2150 8754 2202
rect 8754 2150 8800 2202
rect 8504 2148 8560 2150
rect 8584 2148 8640 2150
rect 8664 2148 8720 2150
rect 8744 2148 8800 2150
rect 12483 10906 12539 10908
rect 12563 10906 12619 10908
rect 12643 10906 12699 10908
rect 12723 10906 12779 10908
rect 12483 10854 12529 10906
rect 12529 10854 12539 10906
rect 12563 10854 12593 10906
rect 12593 10854 12605 10906
rect 12605 10854 12619 10906
rect 12643 10854 12657 10906
rect 12657 10854 12669 10906
rect 12669 10854 12699 10906
rect 12723 10854 12733 10906
rect 12733 10854 12779 10906
rect 12483 10852 12539 10854
rect 12563 10852 12619 10854
rect 12643 10852 12699 10854
rect 12723 10852 12779 10854
rect 12483 9818 12539 9820
rect 12563 9818 12619 9820
rect 12643 9818 12699 9820
rect 12723 9818 12779 9820
rect 12483 9766 12529 9818
rect 12529 9766 12539 9818
rect 12563 9766 12593 9818
rect 12593 9766 12605 9818
rect 12605 9766 12619 9818
rect 12643 9766 12657 9818
rect 12657 9766 12669 9818
rect 12669 9766 12699 9818
rect 12723 9766 12733 9818
rect 12733 9766 12779 9818
rect 12483 9764 12539 9766
rect 12563 9764 12619 9766
rect 12643 9764 12699 9766
rect 12723 9764 12779 9766
rect 12483 8730 12539 8732
rect 12563 8730 12619 8732
rect 12643 8730 12699 8732
rect 12723 8730 12779 8732
rect 12483 8678 12529 8730
rect 12529 8678 12539 8730
rect 12563 8678 12593 8730
rect 12593 8678 12605 8730
rect 12605 8678 12619 8730
rect 12643 8678 12657 8730
rect 12657 8678 12669 8730
rect 12669 8678 12699 8730
rect 12723 8678 12733 8730
rect 12733 8678 12779 8730
rect 12483 8676 12539 8678
rect 12563 8676 12619 8678
rect 12643 8676 12699 8678
rect 12723 8676 12779 8678
rect 11823 8186 11879 8188
rect 11903 8186 11959 8188
rect 11983 8186 12039 8188
rect 12063 8186 12119 8188
rect 11823 8134 11869 8186
rect 11869 8134 11879 8186
rect 11903 8134 11933 8186
rect 11933 8134 11945 8186
rect 11945 8134 11959 8186
rect 11983 8134 11997 8186
rect 11997 8134 12009 8186
rect 12009 8134 12039 8186
rect 12063 8134 12073 8186
rect 12073 8134 12119 8186
rect 11823 8132 11879 8134
rect 11903 8132 11959 8134
rect 11983 8132 12039 8134
rect 12063 8132 12119 8134
rect 11823 7098 11879 7100
rect 11903 7098 11959 7100
rect 11983 7098 12039 7100
rect 12063 7098 12119 7100
rect 11823 7046 11869 7098
rect 11869 7046 11879 7098
rect 11903 7046 11933 7098
rect 11933 7046 11945 7098
rect 11945 7046 11959 7098
rect 11983 7046 11997 7098
rect 11997 7046 12009 7098
rect 12009 7046 12039 7098
rect 12063 7046 12073 7098
rect 12073 7046 12119 7098
rect 11823 7044 11879 7046
rect 11903 7044 11959 7046
rect 11983 7044 12039 7046
rect 12063 7044 12119 7046
rect 12483 7642 12539 7644
rect 12563 7642 12619 7644
rect 12643 7642 12699 7644
rect 12723 7642 12779 7644
rect 12483 7590 12529 7642
rect 12529 7590 12539 7642
rect 12563 7590 12593 7642
rect 12593 7590 12605 7642
rect 12605 7590 12619 7642
rect 12643 7590 12657 7642
rect 12657 7590 12669 7642
rect 12669 7590 12699 7642
rect 12723 7590 12733 7642
rect 12733 7590 12779 7642
rect 12483 7588 12539 7590
rect 12563 7588 12619 7590
rect 12643 7588 12699 7590
rect 12723 7588 12779 7590
rect 15802 13626 15858 13628
rect 15882 13626 15938 13628
rect 15962 13626 16018 13628
rect 16042 13626 16098 13628
rect 15802 13574 15848 13626
rect 15848 13574 15858 13626
rect 15882 13574 15912 13626
rect 15912 13574 15924 13626
rect 15924 13574 15938 13626
rect 15962 13574 15976 13626
rect 15976 13574 15988 13626
rect 15988 13574 16018 13626
rect 16042 13574 16052 13626
rect 16052 13574 16098 13626
rect 15802 13572 15858 13574
rect 15882 13572 15938 13574
rect 15962 13572 16018 13574
rect 16042 13572 16098 13574
rect 16462 13082 16518 13084
rect 16542 13082 16598 13084
rect 16622 13082 16678 13084
rect 16702 13082 16758 13084
rect 16462 13030 16508 13082
rect 16508 13030 16518 13082
rect 16542 13030 16572 13082
rect 16572 13030 16584 13082
rect 16584 13030 16598 13082
rect 16622 13030 16636 13082
rect 16636 13030 16648 13082
rect 16648 13030 16678 13082
rect 16702 13030 16712 13082
rect 16712 13030 16758 13082
rect 16462 13028 16518 13030
rect 16542 13028 16598 13030
rect 16622 13028 16678 13030
rect 16702 13028 16758 13030
rect 15802 12538 15858 12540
rect 15882 12538 15938 12540
rect 15962 12538 16018 12540
rect 16042 12538 16098 12540
rect 15802 12486 15848 12538
rect 15848 12486 15858 12538
rect 15882 12486 15912 12538
rect 15912 12486 15924 12538
rect 15924 12486 15938 12538
rect 15962 12486 15976 12538
rect 15976 12486 15988 12538
rect 15988 12486 16018 12538
rect 16042 12486 16052 12538
rect 16052 12486 16098 12538
rect 15802 12484 15858 12486
rect 15882 12484 15938 12486
rect 15962 12484 16018 12486
rect 16042 12484 16098 12486
rect 16486 12280 16542 12336
rect 16462 11994 16518 11996
rect 16542 11994 16598 11996
rect 16622 11994 16678 11996
rect 16702 11994 16758 11996
rect 16462 11942 16508 11994
rect 16508 11942 16518 11994
rect 16542 11942 16572 11994
rect 16572 11942 16584 11994
rect 16584 11942 16598 11994
rect 16622 11942 16636 11994
rect 16636 11942 16648 11994
rect 16648 11942 16678 11994
rect 16702 11942 16712 11994
rect 16712 11942 16758 11994
rect 16462 11940 16518 11942
rect 16542 11940 16598 11942
rect 16622 11940 16678 11942
rect 16702 11940 16758 11942
rect 17314 11600 17370 11656
rect 15802 11450 15858 11452
rect 15882 11450 15938 11452
rect 15962 11450 16018 11452
rect 16042 11450 16098 11452
rect 15802 11398 15848 11450
rect 15848 11398 15858 11450
rect 15882 11398 15912 11450
rect 15912 11398 15924 11450
rect 15924 11398 15938 11450
rect 15962 11398 15976 11450
rect 15976 11398 15988 11450
rect 15988 11398 16018 11450
rect 16042 11398 16052 11450
rect 16052 11398 16098 11450
rect 15802 11396 15858 11398
rect 15882 11396 15938 11398
rect 15962 11396 16018 11398
rect 16042 11396 16098 11398
rect 17498 10920 17554 10976
rect 16462 10906 16518 10908
rect 16542 10906 16598 10908
rect 16622 10906 16678 10908
rect 16702 10906 16758 10908
rect 16462 10854 16508 10906
rect 16508 10854 16518 10906
rect 16542 10854 16572 10906
rect 16572 10854 16584 10906
rect 16584 10854 16598 10906
rect 16622 10854 16636 10906
rect 16636 10854 16648 10906
rect 16648 10854 16678 10906
rect 16702 10854 16712 10906
rect 16712 10854 16758 10906
rect 16462 10852 16518 10854
rect 16542 10852 16598 10854
rect 16622 10852 16678 10854
rect 16702 10852 16758 10854
rect 15802 10362 15858 10364
rect 15882 10362 15938 10364
rect 15962 10362 16018 10364
rect 16042 10362 16098 10364
rect 15802 10310 15848 10362
rect 15848 10310 15858 10362
rect 15882 10310 15912 10362
rect 15912 10310 15924 10362
rect 15924 10310 15938 10362
rect 15962 10310 15976 10362
rect 15976 10310 15988 10362
rect 15988 10310 16018 10362
rect 16042 10310 16052 10362
rect 16052 10310 16098 10362
rect 15802 10308 15858 10310
rect 15882 10308 15938 10310
rect 15962 10308 16018 10310
rect 16042 10308 16098 10310
rect 17406 10240 17462 10296
rect 16462 9818 16518 9820
rect 16542 9818 16598 9820
rect 16622 9818 16678 9820
rect 16702 9818 16758 9820
rect 16462 9766 16508 9818
rect 16508 9766 16518 9818
rect 16542 9766 16572 9818
rect 16572 9766 16584 9818
rect 16584 9766 16598 9818
rect 16622 9766 16636 9818
rect 16636 9766 16648 9818
rect 16648 9766 16678 9818
rect 16702 9766 16712 9818
rect 16712 9766 16758 9818
rect 16462 9764 16518 9766
rect 16542 9764 16598 9766
rect 16622 9764 16678 9766
rect 16702 9764 16758 9766
rect 17498 9560 17554 9616
rect 15802 9274 15858 9276
rect 15882 9274 15938 9276
rect 15962 9274 16018 9276
rect 16042 9274 16098 9276
rect 15802 9222 15848 9274
rect 15848 9222 15858 9274
rect 15882 9222 15912 9274
rect 15912 9222 15924 9274
rect 15924 9222 15938 9274
rect 15962 9222 15976 9274
rect 15976 9222 15988 9274
rect 15988 9222 16018 9274
rect 16042 9222 16052 9274
rect 16052 9222 16098 9274
rect 15802 9220 15858 9222
rect 15882 9220 15938 9222
rect 15962 9220 16018 9222
rect 16042 9220 16098 9222
rect 11823 6010 11879 6012
rect 11903 6010 11959 6012
rect 11983 6010 12039 6012
rect 12063 6010 12119 6012
rect 11823 5958 11869 6010
rect 11869 5958 11879 6010
rect 11903 5958 11933 6010
rect 11933 5958 11945 6010
rect 11945 5958 11959 6010
rect 11983 5958 11997 6010
rect 11997 5958 12009 6010
rect 12009 5958 12039 6010
rect 12063 5958 12073 6010
rect 12073 5958 12119 6010
rect 11823 5956 11879 5958
rect 11903 5956 11959 5958
rect 11983 5956 12039 5958
rect 12063 5956 12119 5958
rect 11823 4922 11879 4924
rect 11903 4922 11959 4924
rect 11983 4922 12039 4924
rect 12063 4922 12119 4924
rect 11823 4870 11869 4922
rect 11869 4870 11879 4922
rect 11903 4870 11933 4922
rect 11933 4870 11945 4922
rect 11945 4870 11959 4922
rect 11983 4870 11997 4922
rect 11997 4870 12009 4922
rect 12009 4870 12039 4922
rect 12063 4870 12073 4922
rect 12073 4870 12119 4922
rect 11823 4868 11879 4870
rect 11903 4868 11959 4870
rect 11983 4868 12039 4870
rect 12063 4868 12119 4870
rect 11823 3834 11879 3836
rect 11903 3834 11959 3836
rect 11983 3834 12039 3836
rect 12063 3834 12119 3836
rect 11823 3782 11869 3834
rect 11869 3782 11879 3834
rect 11903 3782 11933 3834
rect 11933 3782 11945 3834
rect 11945 3782 11959 3834
rect 11983 3782 11997 3834
rect 11997 3782 12009 3834
rect 12009 3782 12039 3834
rect 12063 3782 12073 3834
rect 12073 3782 12119 3834
rect 11823 3780 11879 3782
rect 11903 3780 11959 3782
rect 11983 3780 12039 3782
rect 12063 3780 12119 3782
rect 11823 2746 11879 2748
rect 11903 2746 11959 2748
rect 11983 2746 12039 2748
rect 12063 2746 12119 2748
rect 11823 2694 11869 2746
rect 11869 2694 11879 2746
rect 11903 2694 11933 2746
rect 11933 2694 11945 2746
rect 11945 2694 11959 2746
rect 11983 2694 11997 2746
rect 11997 2694 12009 2746
rect 12009 2694 12039 2746
rect 12063 2694 12073 2746
rect 12073 2694 12119 2746
rect 11823 2692 11879 2694
rect 11903 2692 11959 2694
rect 11983 2692 12039 2694
rect 12063 2692 12119 2694
rect 12483 6554 12539 6556
rect 12563 6554 12619 6556
rect 12643 6554 12699 6556
rect 12723 6554 12779 6556
rect 12483 6502 12529 6554
rect 12529 6502 12539 6554
rect 12563 6502 12593 6554
rect 12593 6502 12605 6554
rect 12605 6502 12619 6554
rect 12643 6502 12657 6554
rect 12657 6502 12669 6554
rect 12669 6502 12699 6554
rect 12723 6502 12733 6554
rect 12733 6502 12779 6554
rect 12483 6500 12539 6502
rect 12563 6500 12619 6502
rect 12643 6500 12699 6502
rect 12723 6500 12779 6502
rect 12483 5466 12539 5468
rect 12563 5466 12619 5468
rect 12643 5466 12699 5468
rect 12723 5466 12779 5468
rect 12483 5414 12529 5466
rect 12529 5414 12539 5466
rect 12563 5414 12593 5466
rect 12593 5414 12605 5466
rect 12605 5414 12619 5466
rect 12643 5414 12657 5466
rect 12657 5414 12669 5466
rect 12669 5414 12699 5466
rect 12723 5414 12733 5466
rect 12733 5414 12779 5466
rect 12483 5412 12539 5414
rect 12563 5412 12619 5414
rect 12643 5412 12699 5414
rect 12723 5412 12779 5414
rect 12483 4378 12539 4380
rect 12563 4378 12619 4380
rect 12643 4378 12699 4380
rect 12723 4378 12779 4380
rect 12483 4326 12529 4378
rect 12529 4326 12539 4378
rect 12563 4326 12593 4378
rect 12593 4326 12605 4378
rect 12605 4326 12619 4378
rect 12643 4326 12657 4378
rect 12657 4326 12669 4378
rect 12669 4326 12699 4378
rect 12723 4326 12733 4378
rect 12733 4326 12779 4378
rect 12483 4324 12539 4326
rect 12563 4324 12619 4326
rect 12643 4324 12699 4326
rect 12723 4324 12779 4326
rect 12483 3290 12539 3292
rect 12563 3290 12619 3292
rect 12643 3290 12699 3292
rect 12723 3290 12779 3292
rect 12483 3238 12529 3290
rect 12529 3238 12539 3290
rect 12563 3238 12593 3290
rect 12593 3238 12605 3290
rect 12605 3238 12619 3290
rect 12643 3238 12657 3290
rect 12657 3238 12669 3290
rect 12669 3238 12699 3290
rect 12723 3238 12733 3290
rect 12733 3238 12779 3290
rect 12483 3236 12539 3238
rect 12563 3236 12619 3238
rect 12643 3236 12699 3238
rect 12723 3236 12779 3238
rect 17498 8900 17554 8936
rect 17498 8880 17500 8900
rect 17500 8880 17552 8900
rect 17552 8880 17554 8900
rect 16462 8730 16518 8732
rect 16542 8730 16598 8732
rect 16622 8730 16678 8732
rect 16702 8730 16758 8732
rect 16462 8678 16508 8730
rect 16508 8678 16518 8730
rect 16542 8678 16572 8730
rect 16572 8678 16584 8730
rect 16584 8678 16598 8730
rect 16622 8678 16636 8730
rect 16636 8678 16648 8730
rect 16648 8678 16678 8730
rect 16702 8678 16712 8730
rect 16712 8678 16758 8730
rect 16462 8676 16518 8678
rect 16542 8676 16598 8678
rect 16622 8676 16678 8678
rect 16702 8676 16758 8678
rect 17314 8200 17370 8256
rect 15802 8186 15858 8188
rect 15882 8186 15938 8188
rect 15962 8186 16018 8188
rect 16042 8186 16098 8188
rect 15802 8134 15848 8186
rect 15848 8134 15858 8186
rect 15882 8134 15912 8186
rect 15912 8134 15924 8186
rect 15924 8134 15938 8186
rect 15962 8134 15976 8186
rect 15976 8134 15988 8186
rect 15988 8134 16018 8186
rect 16042 8134 16052 8186
rect 16052 8134 16098 8186
rect 15802 8132 15858 8134
rect 15882 8132 15938 8134
rect 15962 8132 16018 8134
rect 16042 8132 16098 8134
rect 16462 7642 16518 7644
rect 16542 7642 16598 7644
rect 16622 7642 16678 7644
rect 16702 7642 16758 7644
rect 16462 7590 16508 7642
rect 16508 7590 16518 7642
rect 16542 7590 16572 7642
rect 16572 7590 16584 7642
rect 16584 7590 16598 7642
rect 16622 7590 16636 7642
rect 16636 7590 16648 7642
rect 16648 7590 16678 7642
rect 16702 7590 16712 7642
rect 16712 7590 16758 7642
rect 16462 7588 16518 7590
rect 16542 7588 16598 7590
rect 16622 7588 16678 7590
rect 16702 7588 16758 7590
rect 15802 7098 15858 7100
rect 15882 7098 15938 7100
rect 15962 7098 16018 7100
rect 16042 7098 16098 7100
rect 15802 7046 15848 7098
rect 15848 7046 15858 7098
rect 15882 7046 15912 7098
rect 15912 7046 15924 7098
rect 15924 7046 15938 7098
rect 15962 7046 15976 7098
rect 15976 7046 15988 7098
rect 15988 7046 16018 7098
rect 16042 7046 16052 7098
rect 16052 7046 16098 7098
rect 15802 7044 15858 7046
rect 15882 7044 15938 7046
rect 15962 7044 16018 7046
rect 16042 7044 16098 7046
rect 17590 7520 17646 7576
rect 16462 6554 16518 6556
rect 16542 6554 16598 6556
rect 16622 6554 16678 6556
rect 16702 6554 16758 6556
rect 16462 6502 16508 6554
rect 16508 6502 16518 6554
rect 16542 6502 16572 6554
rect 16572 6502 16584 6554
rect 16584 6502 16598 6554
rect 16622 6502 16636 6554
rect 16636 6502 16648 6554
rect 16648 6502 16678 6554
rect 16702 6502 16712 6554
rect 16712 6502 16758 6554
rect 16462 6500 16518 6502
rect 16542 6500 16598 6502
rect 16622 6500 16678 6502
rect 16702 6500 16758 6502
rect 15802 6010 15858 6012
rect 15882 6010 15938 6012
rect 15962 6010 16018 6012
rect 16042 6010 16098 6012
rect 15802 5958 15848 6010
rect 15848 5958 15858 6010
rect 15882 5958 15912 6010
rect 15912 5958 15924 6010
rect 15924 5958 15938 6010
rect 15962 5958 15976 6010
rect 15976 5958 15988 6010
rect 15988 5958 16018 6010
rect 16042 5958 16052 6010
rect 16052 5958 16098 6010
rect 15802 5956 15858 5958
rect 15882 5956 15938 5958
rect 15962 5956 16018 5958
rect 16042 5956 16098 5958
rect 16462 5466 16518 5468
rect 16542 5466 16598 5468
rect 16622 5466 16678 5468
rect 16702 5466 16758 5468
rect 16462 5414 16508 5466
rect 16508 5414 16518 5466
rect 16542 5414 16572 5466
rect 16572 5414 16584 5466
rect 16584 5414 16598 5466
rect 16622 5414 16636 5466
rect 16636 5414 16648 5466
rect 16648 5414 16678 5466
rect 16702 5414 16712 5466
rect 16712 5414 16758 5466
rect 16462 5412 16518 5414
rect 16542 5412 16598 5414
rect 16622 5412 16678 5414
rect 16702 5412 16758 5414
rect 15802 4922 15858 4924
rect 15882 4922 15938 4924
rect 15962 4922 16018 4924
rect 16042 4922 16098 4924
rect 15802 4870 15848 4922
rect 15848 4870 15858 4922
rect 15882 4870 15912 4922
rect 15912 4870 15924 4922
rect 15924 4870 15938 4922
rect 15962 4870 15976 4922
rect 15976 4870 15988 4922
rect 15988 4870 16018 4922
rect 16042 4870 16052 4922
rect 16052 4870 16098 4922
rect 15802 4868 15858 4870
rect 15882 4868 15938 4870
rect 15962 4868 16018 4870
rect 16042 4868 16098 4870
rect 16462 4378 16518 4380
rect 16542 4378 16598 4380
rect 16622 4378 16678 4380
rect 16702 4378 16758 4380
rect 16462 4326 16508 4378
rect 16508 4326 16518 4378
rect 16542 4326 16572 4378
rect 16572 4326 16584 4378
rect 16584 4326 16598 4378
rect 16622 4326 16636 4378
rect 16636 4326 16648 4378
rect 16648 4326 16678 4378
rect 16702 4326 16712 4378
rect 16712 4326 16758 4378
rect 16462 4324 16518 4326
rect 16542 4324 16598 4326
rect 16622 4324 16678 4326
rect 16702 4324 16758 4326
rect 15802 3834 15858 3836
rect 15882 3834 15938 3836
rect 15962 3834 16018 3836
rect 16042 3834 16098 3836
rect 15802 3782 15848 3834
rect 15848 3782 15858 3834
rect 15882 3782 15912 3834
rect 15912 3782 15924 3834
rect 15924 3782 15938 3834
rect 15962 3782 15976 3834
rect 15976 3782 15988 3834
rect 15988 3782 16018 3834
rect 16042 3782 16052 3834
rect 16052 3782 16098 3834
rect 15802 3780 15858 3782
rect 15882 3780 15938 3782
rect 15962 3780 16018 3782
rect 16042 3780 16098 3782
rect 16462 3290 16518 3292
rect 16542 3290 16598 3292
rect 16622 3290 16678 3292
rect 16702 3290 16758 3292
rect 16462 3238 16508 3290
rect 16508 3238 16518 3290
rect 16542 3238 16572 3290
rect 16572 3238 16584 3290
rect 16584 3238 16598 3290
rect 16622 3238 16636 3290
rect 16636 3238 16648 3290
rect 16648 3238 16678 3290
rect 16702 3238 16712 3290
rect 16712 3238 16758 3290
rect 16462 3236 16518 3238
rect 16542 3236 16598 3238
rect 16622 3236 16678 3238
rect 16702 3236 16758 3238
rect 15802 2746 15858 2748
rect 15882 2746 15938 2748
rect 15962 2746 16018 2748
rect 16042 2746 16098 2748
rect 15802 2694 15848 2746
rect 15848 2694 15858 2746
rect 15882 2694 15912 2746
rect 15912 2694 15924 2746
rect 15924 2694 15938 2746
rect 15962 2694 15976 2746
rect 15976 2694 15988 2746
rect 15988 2694 16018 2746
rect 16042 2694 16052 2746
rect 16052 2694 16098 2746
rect 15802 2692 15858 2694
rect 15882 2692 15938 2694
rect 15962 2692 16018 2694
rect 16042 2692 16098 2694
rect 12483 2202 12539 2204
rect 12563 2202 12619 2204
rect 12643 2202 12699 2204
rect 12723 2202 12779 2204
rect 12483 2150 12529 2202
rect 12529 2150 12539 2202
rect 12563 2150 12593 2202
rect 12593 2150 12605 2202
rect 12605 2150 12619 2202
rect 12643 2150 12657 2202
rect 12657 2150 12669 2202
rect 12669 2150 12699 2202
rect 12723 2150 12733 2202
rect 12733 2150 12779 2202
rect 12483 2148 12539 2150
rect 12563 2148 12619 2150
rect 12643 2148 12699 2150
rect 12723 2148 12779 2150
rect 16462 2202 16518 2204
rect 16542 2202 16598 2204
rect 16622 2202 16678 2204
rect 16702 2202 16758 2204
rect 16462 2150 16508 2202
rect 16508 2150 16518 2202
rect 16542 2150 16572 2202
rect 16572 2150 16584 2202
rect 16584 2150 16598 2202
rect 16622 2150 16636 2202
rect 16636 2150 16648 2202
rect 16648 2150 16678 2202
rect 16702 2150 16712 2202
rect 16712 2150 16758 2202
rect 16462 2148 16518 2150
rect 16542 2148 16598 2150
rect 16622 2148 16678 2150
rect 16702 2148 16758 2150
<< metal3 >>
rect 3855 17984 4171 17985
rect 3855 17920 3861 17984
rect 3925 17920 3941 17984
rect 4005 17920 4021 17984
rect 4085 17920 4101 17984
rect 4165 17920 4171 17984
rect 3855 17919 4171 17920
rect 7834 17984 8150 17985
rect 7834 17920 7840 17984
rect 7904 17920 7920 17984
rect 7984 17920 8000 17984
rect 8064 17920 8080 17984
rect 8144 17920 8150 17984
rect 7834 17919 8150 17920
rect 11813 17984 12129 17985
rect 11813 17920 11819 17984
rect 11883 17920 11899 17984
rect 11963 17920 11979 17984
rect 12043 17920 12059 17984
rect 12123 17920 12129 17984
rect 11813 17919 12129 17920
rect 15792 17984 16108 17985
rect 15792 17920 15798 17984
rect 15862 17920 15878 17984
rect 15942 17920 15958 17984
rect 16022 17920 16038 17984
rect 16102 17920 16108 17984
rect 15792 17919 16108 17920
rect 4515 17440 4831 17441
rect 4515 17376 4521 17440
rect 4585 17376 4601 17440
rect 4665 17376 4681 17440
rect 4745 17376 4761 17440
rect 4825 17376 4831 17440
rect 4515 17375 4831 17376
rect 8494 17440 8810 17441
rect 8494 17376 8500 17440
rect 8564 17376 8580 17440
rect 8644 17376 8660 17440
rect 8724 17376 8740 17440
rect 8804 17376 8810 17440
rect 8494 17375 8810 17376
rect 12473 17440 12789 17441
rect 12473 17376 12479 17440
rect 12543 17376 12559 17440
rect 12623 17376 12639 17440
rect 12703 17376 12719 17440
rect 12783 17376 12789 17440
rect 12473 17375 12789 17376
rect 16452 17440 16768 17441
rect 16452 17376 16458 17440
rect 16522 17376 16538 17440
rect 16602 17376 16618 17440
rect 16682 17376 16698 17440
rect 16762 17376 16768 17440
rect 16452 17375 16768 17376
rect 3855 16896 4171 16897
rect 3855 16832 3861 16896
rect 3925 16832 3941 16896
rect 4005 16832 4021 16896
rect 4085 16832 4101 16896
rect 4165 16832 4171 16896
rect 3855 16831 4171 16832
rect 7834 16896 8150 16897
rect 7834 16832 7840 16896
rect 7904 16832 7920 16896
rect 7984 16832 8000 16896
rect 8064 16832 8080 16896
rect 8144 16832 8150 16896
rect 7834 16831 8150 16832
rect 11813 16896 12129 16897
rect 11813 16832 11819 16896
rect 11883 16832 11899 16896
rect 11963 16832 11979 16896
rect 12043 16832 12059 16896
rect 12123 16832 12129 16896
rect 11813 16831 12129 16832
rect 15792 16896 16108 16897
rect 15792 16832 15798 16896
rect 15862 16832 15878 16896
rect 15942 16832 15958 16896
rect 16022 16832 16038 16896
rect 16102 16832 16108 16896
rect 15792 16831 16108 16832
rect 4515 16352 4831 16353
rect 4515 16288 4521 16352
rect 4585 16288 4601 16352
rect 4665 16288 4681 16352
rect 4745 16288 4761 16352
rect 4825 16288 4831 16352
rect 4515 16287 4831 16288
rect 8494 16352 8810 16353
rect 8494 16288 8500 16352
rect 8564 16288 8580 16352
rect 8644 16288 8660 16352
rect 8724 16288 8740 16352
rect 8804 16288 8810 16352
rect 8494 16287 8810 16288
rect 12473 16352 12789 16353
rect 12473 16288 12479 16352
rect 12543 16288 12559 16352
rect 12623 16288 12639 16352
rect 12703 16288 12719 16352
rect 12783 16288 12789 16352
rect 12473 16287 12789 16288
rect 16452 16352 16768 16353
rect 16452 16288 16458 16352
rect 16522 16288 16538 16352
rect 16602 16288 16618 16352
rect 16682 16288 16698 16352
rect 16762 16288 16768 16352
rect 16452 16287 16768 16288
rect 3855 15808 4171 15809
rect 3855 15744 3861 15808
rect 3925 15744 3941 15808
rect 4005 15744 4021 15808
rect 4085 15744 4101 15808
rect 4165 15744 4171 15808
rect 3855 15743 4171 15744
rect 7834 15808 8150 15809
rect 7834 15744 7840 15808
rect 7904 15744 7920 15808
rect 7984 15744 8000 15808
rect 8064 15744 8080 15808
rect 8144 15744 8150 15808
rect 7834 15743 8150 15744
rect 11813 15808 12129 15809
rect 11813 15744 11819 15808
rect 11883 15744 11899 15808
rect 11963 15744 11979 15808
rect 12043 15744 12059 15808
rect 12123 15744 12129 15808
rect 11813 15743 12129 15744
rect 15792 15808 16108 15809
rect 15792 15744 15798 15808
rect 15862 15744 15878 15808
rect 15942 15744 15958 15808
rect 16022 15744 16038 15808
rect 16102 15744 16108 15808
rect 15792 15743 16108 15744
rect 4515 15264 4831 15265
rect 4515 15200 4521 15264
rect 4585 15200 4601 15264
rect 4665 15200 4681 15264
rect 4745 15200 4761 15264
rect 4825 15200 4831 15264
rect 4515 15199 4831 15200
rect 8494 15264 8810 15265
rect 8494 15200 8500 15264
rect 8564 15200 8580 15264
rect 8644 15200 8660 15264
rect 8724 15200 8740 15264
rect 8804 15200 8810 15264
rect 8494 15199 8810 15200
rect 12473 15264 12789 15265
rect 12473 15200 12479 15264
rect 12543 15200 12559 15264
rect 12623 15200 12639 15264
rect 12703 15200 12719 15264
rect 12783 15200 12789 15264
rect 12473 15199 12789 15200
rect 16452 15264 16768 15265
rect 16452 15200 16458 15264
rect 16522 15200 16538 15264
rect 16602 15200 16618 15264
rect 16682 15200 16698 15264
rect 16762 15200 16768 15264
rect 16452 15199 16768 15200
rect 3855 14720 4171 14721
rect 3855 14656 3861 14720
rect 3925 14656 3941 14720
rect 4005 14656 4021 14720
rect 4085 14656 4101 14720
rect 4165 14656 4171 14720
rect 3855 14655 4171 14656
rect 7834 14720 8150 14721
rect 7834 14656 7840 14720
rect 7904 14656 7920 14720
rect 7984 14656 8000 14720
rect 8064 14656 8080 14720
rect 8144 14656 8150 14720
rect 7834 14655 8150 14656
rect 11813 14720 12129 14721
rect 11813 14656 11819 14720
rect 11883 14656 11899 14720
rect 11963 14656 11979 14720
rect 12043 14656 12059 14720
rect 12123 14656 12129 14720
rect 11813 14655 12129 14656
rect 15792 14720 16108 14721
rect 15792 14656 15798 14720
rect 15862 14656 15878 14720
rect 15942 14656 15958 14720
rect 16022 14656 16038 14720
rect 16102 14656 16108 14720
rect 15792 14655 16108 14656
rect 4515 14176 4831 14177
rect 4515 14112 4521 14176
rect 4585 14112 4601 14176
rect 4665 14112 4681 14176
rect 4745 14112 4761 14176
rect 4825 14112 4831 14176
rect 4515 14111 4831 14112
rect 8494 14176 8810 14177
rect 8494 14112 8500 14176
rect 8564 14112 8580 14176
rect 8644 14112 8660 14176
rect 8724 14112 8740 14176
rect 8804 14112 8810 14176
rect 8494 14111 8810 14112
rect 12473 14176 12789 14177
rect 12473 14112 12479 14176
rect 12543 14112 12559 14176
rect 12623 14112 12639 14176
rect 12703 14112 12719 14176
rect 12783 14112 12789 14176
rect 12473 14111 12789 14112
rect 16452 14176 16768 14177
rect 16452 14112 16458 14176
rect 16522 14112 16538 14176
rect 16602 14112 16618 14176
rect 16682 14112 16698 14176
rect 16762 14112 16768 14176
rect 16452 14111 16768 14112
rect 3855 13632 4171 13633
rect 3855 13568 3861 13632
rect 3925 13568 3941 13632
rect 4005 13568 4021 13632
rect 4085 13568 4101 13632
rect 4165 13568 4171 13632
rect 3855 13567 4171 13568
rect 7834 13632 8150 13633
rect 7834 13568 7840 13632
rect 7904 13568 7920 13632
rect 7984 13568 8000 13632
rect 8064 13568 8080 13632
rect 8144 13568 8150 13632
rect 7834 13567 8150 13568
rect 11813 13632 12129 13633
rect 11813 13568 11819 13632
rect 11883 13568 11899 13632
rect 11963 13568 11979 13632
rect 12043 13568 12059 13632
rect 12123 13568 12129 13632
rect 11813 13567 12129 13568
rect 15792 13632 16108 13633
rect 15792 13568 15798 13632
rect 15862 13568 15878 13632
rect 15942 13568 15958 13632
rect 16022 13568 16038 13632
rect 16102 13568 16108 13632
rect 15792 13567 16108 13568
rect 4515 13088 4831 13089
rect 4515 13024 4521 13088
rect 4585 13024 4601 13088
rect 4665 13024 4681 13088
rect 4745 13024 4761 13088
rect 4825 13024 4831 13088
rect 4515 13023 4831 13024
rect 8494 13088 8810 13089
rect 8494 13024 8500 13088
rect 8564 13024 8580 13088
rect 8644 13024 8660 13088
rect 8724 13024 8740 13088
rect 8804 13024 8810 13088
rect 8494 13023 8810 13024
rect 12473 13088 12789 13089
rect 12473 13024 12479 13088
rect 12543 13024 12559 13088
rect 12623 13024 12639 13088
rect 12703 13024 12719 13088
rect 12783 13024 12789 13088
rect 12473 13023 12789 13024
rect 16452 13088 16768 13089
rect 16452 13024 16458 13088
rect 16522 13024 16538 13088
rect 16602 13024 16618 13088
rect 16682 13024 16698 13088
rect 16762 13024 16768 13088
rect 16452 13023 16768 13024
rect 3855 12544 4171 12545
rect 3855 12480 3861 12544
rect 3925 12480 3941 12544
rect 4005 12480 4021 12544
rect 4085 12480 4101 12544
rect 4165 12480 4171 12544
rect 3855 12479 4171 12480
rect 7834 12544 8150 12545
rect 7834 12480 7840 12544
rect 7904 12480 7920 12544
rect 7984 12480 8000 12544
rect 8064 12480 8080 12544
rect 8144 12480 8150 12544
rect 7834 12479 8150 12480
rect 11813 12544 12129 12545
rect 11813 12480 11819 12544
rect 11883 12480 11899 12544
rect 11963 12480 11979 12544
rect 12043 12480 12059 12544
rect 12123 12480 12129 12544
rect 11813 12479 12129 12480
rect 15792 12544 16108 12545
rect 15792 12480 15798 12544
rect 15862 12480 15878 12544
rect 15942 12480 15958 12544
rect 16022 12480 16038 12544
rect 16102 12480 16108 12544
rect 15792 12479 16108 12480
rect 0 12338 800 12368
rect 2405 12338 2471 12341
rect 0 12336 2471 12338
rect 0 12280 2410 12336
rect 2466 12280 2471 12336
rect 0 12278 2471 12280
rect 0 12248 800 12278
rect 2405 12275 2471 12278
rect 16481 12338 16547 12341
rect 19200 12338 20000 12368
rect 16481 12336 20000 12338
rect 16481 12280 16486 12336
rect 16542 12280 20000 12336
rect 16481 12278 20000 12280
rect 16481 12275 16547 12278
rect 19200 12248 20000 12278
rect 4515 12000 4831 12001
rect 4515 11936 4521 12000
rect 4585 11936 4601 12000
rect 4665 11936 4681 12000
rect 4745 11936 4761 12000
rect 4825 11936 4831 12000
rect 4515 11935 4831 11936
rect 8494 12000 8810 12001
rect 8494 11936 8500 12000
rect 8564 11936 8580 12000
rect 8644 11936 8660 12000
rect 8724 11936 8740 12000
rect 8804 11936 8810 12000
rect 8494 11935 8810 11936
rect 12473 12000 12789 12001
rect 12473 11936 12479 12000
rect 12543 11936 12559 12000
rect 12623 11936 12639 12000
rect 12703 11936 12719 12000
rect 12783 11936 12789 12000
rect 12473 11935 12789 11936
rect 16452 12000 16768 12001
rect 16452 11936 16458 12000
rect 16522 11936 16538 12000
rect 16602 11936 16618 12000
rect 16682 11936 16698 12000
rect 16762 11936 16768 12000
rect 16452 11935 16768 11936
rect 0 11658 800 11688
rect 1209 11658 1275 11661
rect 0 11656 1275 11658
rect 0 11600 1214 11656
rect 1270 11600 1275 11656
rect 0 11598 1275 11600
rect 0 11568 800 11598
rect 1209 11595 1275 11598
rect 17309 11658 17375 11661
rect 19200 11658 20000 11688
rect 17309 11656 20000 11658
rect 17309 11600 17314 11656
rect 17370 11600 20000 11656
rect 17309 11598 20000 11600
rect 17309 11595 17375 11598
rect 19200 11568 20000 11598
rect 3855 11456 4171 11457
rect 3855 11392 3861 11456
rect 3925 11392 3941 11456
rect 4005 11392 4021 11456
rect 4085 11392 4101 11456
rect 4165 11392 4171 11456
rect 3855 11391 4171 11392
rect 7834 11456 8150 11457
rect 7834 11392 7840 11456
rect 7904 11392 7920 11456
rect 7984 11392 8000 11456
rect 8064 11392 8080 11456
rect 8144 11392 8150 11456
rect 7834 11391 8150 11392
rect 11813 11456 12129 11457
rect 11813 11392 11819 11456
rect 11883 11392 11899 11456
rect 11963 11392 11979 11456
rect 12043 11392 12059 11456
rect 12123 11392 12129 11456
rect 11813 11391 12129 11392
rect 15792 11456 16108 11457
rect 15792 11392 15798 11456
rect 15862 11392 15878 11456
rect 15942 11392 15958 11456
rect 16022 11392 16038 11456
rect 16102 11392 16108 11456
rect 15792 11391 16108 11392
rect 0 10978 800 11008
rect 2313 10978 2379 10981
rect 0 10976 2379 10978
rect 0 10920 2318 10976
rect 2374 10920 2379 10976
rect 0 10918 2379 10920
rect 0 10888 800 10918
rect 2313 10915 2379 10918
rect 17493 10978 17559 10981
rect 19200 10978 20000 11008
rect 17493 10976 20000 10978
rect 17493 10920 17498 10976
rect 17554 10920 20000 10976
rect 17493 10918 20000 10920
rect 17493 10915 17559 10918
rect 4515 10912 4831 10913
rect 4515 10848 4521 10912
rect 4585 10848 4601 10912
rect 4665 10848 4681 10912
rect 4745 10848 4761 10912
rect 4825 10848 4831 10912
rect 4515 10847 4831 10848
rect 8494 10912 8810 10913
rect 8494 10848 8500 10912
rect 8564 10848 8580 10912
rect 8644 10848 8660 10912
rect 8724 10848 8740 10912
rect 8804 10848 8810 10912
rect 8494 10847 8810 10848
rect 12473 10912 12789 10913
rect 12473 10848 12479 10912
rect 12543 10848 12559 10912
rect 12623 10848 12639 10912
rect 12703 10848 12719 10912
rect 12783 10848 12789 10912
rect 12473 10847 12789 10848
rect 16452 10912 16768 10913
rect 16452 10848 16458 10912
rect 16522 10848 16538 10912
rect 16602 10848 16618 10912
rect 16682 10848 16698 10912
rect 16762 10848 16768 10912
rect 19200 10888 20000 10918
rect 16452 10847 16768 10848
rect 3855 10368 4171 10369
rect 0 10298 800 10328
rect 3855 10304 3861 10368
rect 3925 10304 3941 10368
rect 4005 10304 4021 10368
rect 4085 10304 4101 10368
rect 4165 10304 4171 10368
rect 3855 10303 4171 10304
rect 7834 10368 8150 10369
rect 7834 10304 7840 10368
rect 7904 10304 7920 10368
rect 7984 10304 8000 10368
rect 8064 10304 8080 10368
rect 8144 10304 8150 10368
rect 7834 10303 8150 10304
rect 11813 10368 12129 10369
rect 11813 10304 11819 10368
rect 11883 10304 11899 10368
rect 11963 10304 11979 10368
rect 12043 10304 12059 10368
rect 12123 10304 12129 10368
rect 11813 10303 12129 10304
rect 15792 10368 16108 10369
rect 15792 10304 15798 10368
rect 15862 10304 15878 10368
rect 15942 10304 15958 10368
rect 16022 10304 16038 10368
rect 16102 10304 16108 10368
rect 15792 10303 16108 10304
rect 1117 10298 1183 10301
rect 0 10296 1183 10298
rect 0 10240 1122 10296
rect 1178 10240 1183 10296
rect 0 10238 1183 10240
rect 0 10208 800 10238
rect 1117 10235 1183 10238
rect 17401 10298 17467 10301
rect 19200 10298 20000 10328
rect 17401 10296 20000 10298
rect 17401 10240 17406 10296
rect 17462 10240 20000 10296
rect 17401 10238 20000 10240
rect 17401 10235 17467 10238
rect 19200 10208 20000 10238
rect 4515 9824 4831 9825
rect 4515 9760 4521 9824
rect 4585 9760 4601 9824
rect 4665 9760 4681 9824
rect 4745 9760 4761 9824
rect 4825 9760 4831 9824
rect 4515 9759 4831 9760
rect 8494 9824 8810 9825
rect 8494 9760 8500 9824
rect 8564 9760 8580 9824
rect 8644 9760 8660 9824
rect 8724 9760 8740 9824
rect 8804 9760 8810 9824
rect 8494 9759 8810 9760
rect 12473 9824 12789 9825
rect 12473 9760 12479 9824
rect 12543 9760 12559 9824
rect 12623 9760 12639 9824
rect 12703 9760 12719 9824
rect 12783 9760 12789 9824
rect 12473 9759 12789 9760
rect 16452 9824 16768 9825
rect 16452 9760 16458 9824
rect 16522 9760 16538 9824
rect 16602 9760 16618 9824
rect 16682 9760 16698 9824
rect 16762 9760 16768 9824
rect 16452 9759 16768 9760
rect 17493 9618 17559 9621
rect 19200 9618 20000 9648
rect 17493 9616 20000 9618
rect 17493 9560 17498 9616
rect 17554 9560 20000 9616
rect 17493 9558 20000 9560
rect 17493 9555 17559 9558
rect 19200 9528 20000 9558
rect 3855 9280 4171 9281
rect 3855 9216 3861 9280
rect 3925 9216 3941 9280
rect 4005 9216 4021 9280
rect 4085 9216 4101 9280
rect 4165 9216 4171 9280
rect 3855 9215 4171 9216
rect 7834 9280 8150 9281
rect 7834 9216 7840 9280
rect 7904 9216 7920 9280
rect 7984 9216 8000 9280
rect 8064 9216 8080 9280
rect 8144 9216 8150 9280
rect 7834 9215 8150 9216
rect 11813 9280 12129 9281
rect 11813 9216 11819 9280
rect 11883 9216 11899 9280
rect 11963 9216 11979 9280
rect 12043 9216 12059 9280
rect 12123 9216 12129 9280
rect 11813 9215 12129 9216
rect 15792 9280 16108 9281
rect 15792 9216 15798 9280
rect 15862 9216 15878 9280
rect 15942 9216 15958 9280
rect 16022 9216 16038 9280
rect 16102 9216 16108 9280
rect 15792 9215 16108 9216
rect 0 8938 800 8968
rect 1209 8938 1275 8941
rect 0 8936 1275 8938
rect 0 8880 1214 8936
rect 1270 8880 1275 8936
rect 0 8878 1275 8880
rect 0 8848 800 8878
rect 1209 8875 1275 8878
rect 17493 8938 17559 8941
rect 19200 8938 20000 8968
rect 17493 8936 20000 8938
rect 17493 8880 17498 8936
rect 17554 8880 20000 8936
rect 17493 8878 20000 8880
rect 17493 8875 17559 8878
rect 19200 8848 20000 8878
rect 4515 8736 4831 8737
rect 4515 8672 4521 8736
rect 4585 8672 4601 8736
rect 4665 8672 4681 8736
rect 4745 8672 4761 8736
rect 4825 8672 4831 8736
rect 4515 8671 4831 8672
rect 8494 8736 8810 8737
rect 8494 8672 8500 8736
rect 8564 8672 8580 8736
rect 8644 8672 8660 8736
rect 8724 8672 8740 8736
rect 8804 8672 8810 8736
rect 8494 8671 8810 8672
rect 12473 8736 12789 8737
rect 12473 8672 12479 8736
rect 12543 8672 12559 8736
rect 12623 8672 12639 8736
rect 12703 8672 12719 8736
rect 12783 8672 12789 8736
rect 12473 8671 12789 8672
rect 16452 8736 16768 8737
rect 16452 8672 16458 8736
rect 16522 8672 16538 8736
rect 16602 8672 16618 8736
rect 16682 8672 16698 8736
rect 16762 8672 16768 8736
rect 16452 8671 16768 8672
rect 17309 8258 17375 8261
rect 19200 8258 20000 8288
rect 17309 8256 20000 8258
rect 17309 8200 17314 8256
rect 17370 8200 20000 8256
rect 17309 8198 20000 8200
rect 17309 8195 17375 8198
rect 3855 8192 4171 8193
rect 3855 8128 3861 8192
rect 3925 8128 3941 8192
rect 4005 8128 4021 8192
rect 4085 8128 4101 8192
rect 4165 8128 4171 8192
rect 3855 8127 4171 8128
rect 7834 8192 8150 8193
rect 7834 8128 7840 8192
rect 7904 8128 7920 8192
rect 7984 8128 8000 8192
rect 8064 8128 8080 8192
rect 8144 8128 8150 8192
rect 7834 8127 8150 8128
rect 11813 8192 12129 8193
rect 11813 8128 11819 8192
rect 11883 8128 11899 8192
rect 11963 8128 11979 8192
rect 12043 8128 12059 8192
rect 12123 8128 12129 8192
rect 11813 8127 12129 8128
rect 15792 8192 16108 8193
rect 15792 8128 15798 8192
rect 15862 8128 15878 8192
rect 15942 8128 15958 8192
rect 16022 8128 16038 8192
rect 16102 8128 16108 8192
rect 19200 8168 20000 8198
rect 15792 8127 16108 8128
rect 4515 7648 4831 7649
rect 4515 7584 4521 7648
rect 4585 7584 4601 7648
rect 4665 7584 4681 7648
rect 4745 7584 4761 7648
rect 4825 7584 4831 7648
rect 4515 7583 4831 7584
rect 8494 7648 8810 7649
rect 8494 7584 8500 7648
rect 8564 7584 8580 7648
rect 8644 7584 8660 7648
rect 8724 7584 8740 7648
rect 8804 7584 8810 7648
rect 8494 7583 8810 7584
rect 12473 7648 12789 7649
rect 12473 7584 12479 7648
rect 12543 7584 12559 7648
rect 12623 7584 12639 7648
rect 12703 7584 12719 7648
rect 12783 7584 12789 7648
rect 12473 7583 12789 7584
rect 16452 7648 16768 7649
rect 16452 7584 16458 7648
rect 16522 7584 16538 7648
rect 16602 7584 16618 7648
rect 16682 7584 16698 7648
rect 16762 7584 16768 7648
rect 16452 7583 16768 7584
rect 17585 7578 17651 7581
rect 19200 7578 20000 7608
rect 17585 7576 20000 7578
rect 17585 7520 17590 7576
rect 17646 7520 20000 7576
rect 17585 7518 20000 7520
rect 17585 7515 17651 7518
rect 19200 7488 20000 7518
rect 3855 7104 4171 7105
rect 3855 7040 3861 7104
rect 3925 7040 3941 7104
rect 4005 7040 4021 7104
rect 4085 7040 4101 7104
rect 4165 7040 4171 7104
rect 3855 7039 4171 7040
rect 7834 7104 8150 7105
rect 7834 7040 7840 7104
rect 7904 7040 7920 7104
rect 7984 7040 8000 7104
rect 8064 7040 8080 7104
rect 8144 7040 8150 7104
rect 7834 7039 8150 7040
rect 11813 7104 12129 7105
rect 11813 7040 11819 7104
rect 11883 7040 11899 7104
rect 11963 7040 11979 7104
rect 12043 7040 12059 7104
rect 12123 7040 12129 7104
rect 11813 7039 12129 7040
rect 15792 7104 16108 7105
rect 15792 7040 15798 7104
rect 15862 7040 15878 7104
rect 15942 7040 15958 7104
rect 16022 7040 16038 7104
rect 16102 7040 16108 7104
rect 15792 7039 16108 7040
rect 4515 6560 4831 6561
rect 4515 6496 4521 6560
rect 4585 6496 4601 6560
rect 4665 6496 4681 6560
rect 4745 6496 4761 6560
rect 4825 6496 4831 6560
rect 4515 6495 4831 6496
rect 8494 6560 8810 6561
rect 8494 6496 8500 6560
rect 8564 6496 8580 6560
rect 8644 6496 8660 6560
rect 8724 6496 8740 6560
rect 8804 6496 8810 6560
rect 8494 6495 8810 6496
rect 12473 6560 12789 6561
rect 12473 6496 12479 6560
rect 12543 6496 12559 6560
rect 12623 6496 12639 6560
rect 12703 6496 12719 6560
rect 12783 6496 12789 6560
rect 12473 6495 12789 6496
rect 16452 6560 16768 6561
rect 16452 6496 16458 6560
rect 16522 6496 16538 6560
rect 16602 6496 16618 6560
rect 16682 6496 16698 6560
rect 16762 6496 16768 6560
rect 16452 6495 16768 6496
rect 3855 6016 4171 6017
rect 3855 5952 3861 6016
rect 3925 5952 3941 6016
rect 4005 5952 4021 6016
rect 4085 5952 4101 6016
rect 4165 5952 4171 6016
rect 3855 5951 4171 5952
rect 7834 6016 8150 6017
rect 7834 5952 7840 6016
rect 7904 5952 7920 6016
rect 7984 5952 8000 6016
rect 8064 5952 8080 6016
rect 8144 5952 8150 6016
rect 7834 5951 8150 5952
rect 11813 6016 12129 6017
rect 11813 5952 11819 6016
rect 11883 5952 11899 6016
rect 11963 5952 11979 6016
rect 12043 5952 12059 6016
rect 12123 5952 12129 6016
rect 11813 5951 12129 5952
rect 15792 6016 16108 6017
rect 15792 5952 15798 6016
rect 15862 5952 15878 6016
rect 15942 5952 15958 6016
rect 16022 5952 16038 6016
rect 16102 5952 16108 6016
rect 15792 5951 16108 5952
rect 4515 5472 4831 5473
rect 4515 5408 4521 5472
rect 4585 5408 4601 5472
rect 4665 5408 4681 5472
rect 4745 5408 4761 5472
rect 4825 5408 4831 5472
rect 4515 5407 4831 5408
rect 8494 5472 8810 5473
rect 8494 5408 8500 5472
rect 8564 5408 8580 5472
rect 8644 5408 8660 5472
rect 8724 5408 8740 5472
rect 8804 5408 8810 5472
rect 8494 5407 8810 5408
rect 12473 5472 12789 5473
rect 12473 5408 12479 5472
rect 12543 5408 12559 5472
rect 12623 5408 12639 5472
rect 12703 5408 12719 5472
rect 12783 5408 12789 5472
rect 12473 5407 12789 5408
rect 16452 5472 16768 5473
rect 16452 5408 16458 5472
rect 16522 5408 16538 5472
rect 16602 5408 16618 5472
rect 16682 5408 16698 5472
rect 16762 5408 16768 5472
rect 16452 5407 16768 5408
rect 3855 4928 4171 4929
rect 3855 4864 3861 4928
rect 3925 4864 3941 4928
rect 4005 4864 4021 4928
rect 4085 4864 4101 4928
rect 4165 4864 4171 4928
rect 3855 4863 4171 4864
rect 7834 4928 8150 4929
rect 7834 4864 7840 4928
rect 7904 4864 7920 4928
rect 7984 4864 8000 4928
rect 8064 4864 8080 4928
rect 8144 4864 8150 4928
rect 7834 4863 8150 4864
rect 11813 4928 12129 4929
rect 11813 4864 11819 4928
rect 11883 4864 11899 4928
rect 11963 4864 11979 4928
rect 12043 4864 12059 4928
rect 12123 4864 12129 4928
rect 11813 4863 12129 4864
rect 15792 4928 16108 4929
rect 15792 4864 15798 4928
rect 15862 4864 15878 4928
rect 15942 4864 15958 4928
rect 16022 4864 16038 4928
rect 16102 4864 16108 4928
rect 15792 4863 16108 4864
rect 4515 4384 4831 4385
rect 4515 4320 4521 4384
rect 4585 4320 4601 4384
rect 4665 4320 4681 4384
rect 4745 4320 4761 4384
rect 4825 4320 4831 4384
rect 4515 4319 4831 4320
rect 8494 4384 8810 4385
rect 8494 4320 8500 4384
rect 8564 4320 8580 4384
rect 8644 4320 8660 4384
rect 8724 4320 8740 4384
rect 8804 4320 8810 4384
rect 8494 4319 8810 4320
rect 12473 4384 12789 4385
rect 12473 4320 12479 4384
rect 12543 4320 12559 4384
rect 12623 4320 12639 4384
rect 12703 4320 12719 4384
rect 12783 4320 12789 4384
rect 12473 4319 12789 4320
rect 16452 4384 16768 4385
rect 16452 4320 16458 4384
rect 16522 4320 16538 4384
rect 16602 4320 16618 4384
rect 16682 4320 16698 4384
rect 16762 4320 16768 4384
rect 16452 4319 16768 4320
rect 3855 3840 4171 3841
rect 3855 3776 3861 3840
rect 3925 3776 3941 3840
rect 4005 3776 4021 3840
rect 4085 3776 4101 3840
rect 4165 3776 4171 3840
rect 3855 3775 4171 3776
rect 7834 3840 8150 3841
rect 7834 3776 7840 3840
rect 7904 3776 7920 3840
rect 7984 3776 8000 3840
rect 8064 3776 8080 3840
rect 8144 3776 8150 3840
rect 7834 3775 8150 3776
rect 11813 3840 12129 3841
rect 11813 3776 11819 3840
rect 11883 3776 11899 3840
rect 11963 3776 11979 3840
rect 12043 3776 12059 3840
rect 12123 3776 12129 3840
rect 11813 3775 12129 3776
rect 15792 3840 16108 3841
rect 15792 3776 15798 3840
rect 15862 3776 15878 3840
rect 15942 3776 15958 3840
rect 16022 3776 16038 3840
rect 16102 3776 16108 3840
rect 15792 3775 16108 3776
rect 4515 3296 4831 3297
rect 4515 3232 4521 3296
rect 4585 3232 4601 3296
rect 4665 3232 4681 3296
rect 4745 3232 4761 3296
rect 4825 3232 4831 3296
rect 4515 3231 4831 3232
rect 8494 3296 8810 3297
rect 8494 3232 8500 3296
rect 8564 3232 8580 3296
rect 8644 3232 8660 3296
rect 8724 3232 8740 3296
rect 8804 3232 8810 3296
rect 8494 3231 8810 3232
rect 12473 3296 12789 3297
rect 12473 3232 12479 3296
rect 12543 3232 12559 3296
rect 12623 3232 12639 3296
rect 12703 3232 12719 3296
rect 12783 3232 12789 3296
rect 12473 3231 12789 3232
rect 16452 3296 16768 3297
rect 16452 3232 16458 3296
rect 16522 3232 16538 3296
rect 16602 3232 16618 3296
rect 16682 3232 16698 3296
rect 16762 3232 16768 3296
rect 16452 3231 16768 3232
rect 3855 2752 4171 2753
rect 3855 2688 3861 2752
rect 3925 2688 3941 2752
rect 4005 2688 4021 2752
rect 4085 2688 4101 2752
rect 4165 2688 4171 2752
rect 3855 2687 4171 2688
rect 7834 2752 8150 2753
rect 7834 2688 7840 2752
rect 7904 2688 7920 2752
rect 7984 2688 8000 2752
rect 8064 2688 8080 2752
rect 8144 2688 8150 2752
rect 7834 2687 8150 2688
rect 11813 2752 12129 2753
rect 11813 2688 11819 2752
rect 11883 2688 11899 2752
rect 11963 2688 11979 2752
rect 12043 2688 12059 2752
rect 12123 2688 12129 2752
rect 11813 2687 12129 2688
rect 15792 2752 16108 2753
rect 15792 2688 15798 2752
rect 15862 2688 15878 2752
rect 15942 2688 15958 2752
rect 16022 2688 16038 2752
rect 16102 2688 16108 2752
rect 15792 2687 16108 2688
rect 4515 2208 4831 2209
rect 4515 2144 4521 2208
rect 4585 2144 4601 2208
rect 4665 2144 4681 2208
rect 4745 2144 4761 2208
rect 4825 2144 4831 2208
rect 4515 2143 4831 2144
rect 8494 2208 8810 2209
rect 8494 2144 8500 2208
rect 8564 2144 8580 2208
rect 8644 2144 8660 2208
rect 8724 2144 8740 2208
rect 8804 2144 8810 2208
rect 8494 2143 8810 2144
rect 12473 2208 12789 2209
rect 12473 2144 12479 2208
rect 12543 2144 12559 2208
rect 12623 2144 12639 2208
rect 12703 2144 12719 2208
rect 12783 2144 12789 2208
rect 12473 2143 12789 2144
rect 16452 2208 16768 2209
rect 16452 2144 16458 2208
rect 16522 2144 16538 2208
rect 16602 2144 16618 2208
rect 16682 2144 16698 2208
rect 16762 2144 16768 2208
rect 16452 2143 16768 2144
<< via3 >>
rect 3861 17980 3925 17984
rect 3861 17924 3865 17980
rect 3865 17924 3921 17980
rect 3921 17924 3925 17980
rect 3861 17920 3925 17924
rect 3941 17980 4005 17984
rect 3941 17924 3945 17980
rect 3945 17924 4001 17980
rect 4001 17924 4005 17980
rect 3941 17920 4005 17924
rect 4021 17980 4085 17984
rect 4021 17924 4025 17980
rect 4025 17924 4081 17980
rect 4081 17924 4085 17980
rect 4021 17920 4085 17924
rect 4101 17980 4165 17984
rect 4101 17924 4105 17980
rect 4105 17924 4161 17980
rect 4161 17924 4165 17980
rect 4101 17920 4165 17924
rect 7840 17980 7904 17984
rect 7840 17924 7844 17980
rect 7844 17924 7900 17980
rect 7900 17924 7904 17980
rect 7840 17920 7904 17924
rect 7920 17980 7984 17984
rect 7920 17924 7924 17980
rect 7924 17924 7980 17980
rect 7980 17924 7984 17980
rect 7920 17920 7984 17924
rect 8000 17980 8064 17984
rect 8000 17924 8004 17980
rect 8004 17924 8060 17980
rect 8060 17924 8064 17980
rect 8000 17920 8064 17924
rect 8080 17980 8144 17984
rect 8080 17924 8084 17980
rect 8084 17924 8140 17980
rect 8140 17924 8144 17980
rect 8080 17920 8144 17924
rect 11819 17980 11883 17984
rect 11819 17924 11823 17980
rect 11823 17924 11879 17980
rect 11879 17924 11883 17980
rect 11819 17920 11883 17924
rect 11899 17980 11963 17984
rect 11899 17924 11903 17980
rect 11903 17924 11959 17980
rect 11959 17924 11963 17980
rect 11899 17920 11963 17924
rect 11979 17980 12043 17984
rect 11979 17924 11983 17980
rect 11983 17924 12039 17980
rect 12039 17924 12043 17980
rect 11979 17920 12043 17924
rect 12059 17980 12123 17984
rect 12059 17924 12063 17980
rect 12063 17924 12119 17980
rect 12119 17924 12123 17980
rect 12059 17920 12123 17924
rect 15798 17980 15862 17984
rect 15798 17924 15802 17980
rect 15802 17924 15858 17980
rect 15858 17924 15862 17980
rect 15798 17920 15862 17924
rect 15878 17980 15942 17984
rect 15878 17924 15882 17980
rect 15882 17924 15938 17980
rect 15938 17924 15942 17980
rect 15878 17920 15942 17924
rect 15958 17980 16022 17984
rect 15958 17924 15962 17980
rect 15962 17924 16018 17980
rect 16018 17924 16022 17980
rect 15958 17920 16022 17924
rect 16038 17980 16102 17984
rect 16038 17924 16042 17980
rect 16042 17924 16098 17980
rect 16098 17924 16102 17980
rect 16038 17920 16102 17924
rect 4521 17436 4585 17440
rect 4521 17380 4525 17436
rect 4525 17380 4581 17436
rect 4581 17380 4585 17436
rect 4521 17376 4585 17380
rect 4601 17436 4665 17440
rect 4601 17380 4605 17436
rect 4605 17380 4661 17436
rect 4661 17380 4665 17436
rect 4601 17376 4665 17380
rect 4681 17436 4745 17440
rect 4681 17380 4685 17436
rect 4685 17380 4741 17436
rect 4741 17380 4745 17436
rect 4681 17376 4745 17380
rect 4761 17436 4825 17440
rect 4761 17380 4765 17436
rect 4765 17380 4821 17436
rect 4821 17380 4825 17436
rect 4761 17376 4825 17380
rect 8500 17436 8564 17440
rect 8500 17380 8504 17436
rect 8504 17380 8560 17436
rect 8560 17380 8564 17436
rect 8500 17376 8564 17380
rect 8580 17436 8644 17440
rect 8580 17380 8584 17436
rect 8584 17380 8640 17436
rect 8640 17380 8644 17436
rect 8580 17376 8644 17380
rect 8660 17436 8724 17440
rect 8660 17380 8664 17436
rect 8664 17380 8720 17436
rect 8720 17380 8724 17436
rect 8660 17376 8724 17380
rect 8740 17436 8804 17440
rect 8740 17380 8744 17436
rect 8744 17380 8800 17436
rect 8800 17380 8804 17436
rect 8740 17376 8804 17380
rect 12479 17436 12543 17440
rect 12479 17380 12483 17436
rect 12483 17380 12539 17436
rect 12539 17380 12543 17436
rect 12479 17376 12543 17380
rect 12559 17436 12623 17440
rect 12559 17380 12563 17436
rect 12563 17380 12619 17436
rect 12619 17380 12623 17436
rect 12559 17376 12623 17380
rect 12639 17436 12703 17440
rect 12639 17380 12643 17436
rect 12643 17380 12699 17436
rect 12699 17380 12703 17436
rect 12639 17376 12703 17380
rect 12719 17436 12783 17440
rect 12719 17380 12723 17436
rect 12723 17380 12779 17436
rect 12779 17380 12783 17436
rect 12719 17376 12783 17380
rect 16458 17436 16522 17440
rect 16458 17380 16462 17436
rect 16462 17380 16518 17436
rect 16518 17380 16522 17436
rect 16458 17376 16522 17380
rect 16538 17436 16602 17440
rect 16538 17380 16542 17436
rect 16542 17380 16598 17436
rect 16598 17380 16602 17436
rect 16538 17376 16602 17380
rect 16618 17436 16682 17440
rect 16618 17380 16622 17436
rect 16622 17380 16678 17436
rect 16678 17380 16682 17436
rect 16618 17376 16682 17380
rect 16698 17436 16762 17440
rect 16698 17380 16702 17436
rect 16702 17380 16758 17436
rect 16758 17380 16762 17436
rect 16698 17376 16762 17380
rect 3861 16892 3925 16896
rect 3861 16836 3865 16892
rect 3865 16836 3921 16892
rect 3921 16836 3925 16892
rect 3861 16832 3925 16836
rect 3941 16892 4005 16896
rect 3941 16836 3945 16892
rect 3945 16836 4001 16892
rect 4001 16836 4005 16892
rect 3941 16832 4005 16836
rect 4021 16892 4085 16896
rect 4021 16836 4025 16892
rect 4025 16836 4081 16892
rect 4081 16836 4085 16892
rect 4021 16832 4085 16836
rect 4101 16892 4165 16896
rect 4101 16836 4105 16892
rect 4105 16836 4161 16892
rect 4161 16836 4165 16892
rect 4101 16832 4165 16836
rect 7840 16892 7904 16896
rect 7840 16836 7844 16892
rect 7844 16836 7900 16892
rect 7900 16836 7904 16892
rect 7840 16832 7904 16836
rect 7920 16892 7984 16896
rect 7920 16836 7924 16892
rect 7924 16836 7980 16892
rect 7980 16836 7984 16892
rect 7920 16832 7984 16836
rect 8000 16892 8064 16896
rect 8000 16836 8004 16892
rect 8004 16836 8060 16892
rect 8060 16836 8064 16892
rect 8000 16832 8064 16836
rect 8080 16892 8144 16896
rect 8080 16836 8084 16892
rect 8084 16836 8140 16892
rect 8140 16836 8144 16892
rect 8080 16832 8144 16836
rect 11819 16892 11883 16896
rect 11819 16836 11823 16892
rect 11823 16836 11879 16892
rect 11879 16836 11883 16892
rect 11819 16832 11883 16836
rect 11899 16892 11963 16896
rect 11899 16836 11903 16892
rect 11903 16836 11959 16892
rect 11959 16836 11963 16892
rect 11899 16832 11963 16836
rect 11979 16892 12043 16896
rect 11979 16836 11983 16892
rect 11983 16836 12039 16892
rect 12039 16836 12043 16892
rect 11979 16832 12043 16836
rect 12059 16892 12123 16896
rect 12059 16836 12063 16892
rect 12063 16836 12119 16892
rect 12119 16836 12123 16892
rect 12059 16832 12123 16836
rect 15798 16892 15862 16896
rect 15798 16836 15802 16892
rect 15802 16836 15858 16892
rect 15858 16836 15862 16892
rect 15798 16832 15862 16836
rect 15878 16892 15942 16896
rect 15878 16836 15882 16892
rect 15882 16836 15938 16892
rect 15938 16836 15942 16892
rect 15878 16832 15942 16836
rect 15958 16892 16022 16896
rect 15958 16836 15962 16892
rect 15962 16836 16018 16892
rect 16018 16836 16022 16892
rect 15958 16832 16022 16836
rect 16038 16892 16102 16896
rect 16038 16836 16042 16892
rect 16042 16836 16098 16892
rect 16098 16836 16102 16892
rect 16038 16832 16102 16836
rect 4521 16348 4585 16352
rect 4521 16292 4525 16348
rect 4525 16292 4581 16348
rect 4581 16292 4585 16348
rect 4521 16288 4585 16292
rect 4601 16348 4665 16352
rect 4601 16292 4605 16348
rect 4605 16292 4661 16348
rect 4661 16292 4665 16348
rect 4601 16288 4665 16292
rect 4681 16348 4745 16352
rect 4681 16292 4685 16348
rect 4685 16292 4741 16348
rect 4741 16292 4745 16348
rect 4681 16288 4745 16292
rect 4761 16348 4825 16352
rect 4761 16292 4765 16348
rect 4765 16292 4821 16348
rect 4821 16292 4825 16348
rect 4761 16288 4825 16292
rect 8500 16348 8564 16352
rect 8500 16292 8504 16348
rect 8504 16292 8560 16348
rect 8560 16292 8564 16348
rect 8500 16288 8564 16292
rect 8580 16348 8644 16352
rect 8580 16292 8584 16348
rect 8584 16292 8640 16348
rect 8640 16292 8644 16348
rect 8580 16288 8644 16292
rect 8660 16348 8724 16352
rect 8660 16292 8664 16348
rect 8664 16292 8720 16348
rect 8720 16292 8724 16348
rect 8660 16288 8724 16292
rect 8740 16348 8804 16352
rect 8740 16292 8744 16348
rect 8744 16292 8800 16348
rect 8800 16292 8804 16348
rect 8740 16288 8804 16292
rect 12479 16348 12543 16352
rect 12479 16292 12483 16348
rect 12483 16292 12539 16348
rect 12539 16292 12543 16348
rect 12479 16288 12543 16292
rect 12559 16348 12623 16352
rect 12559 16292 12563 16348
rect 12563 16292 12619 16348
rect 12619 16292 12623 16348
rect 12559 16288 12623 16292
rect 12639 16348 12703 16352
rect 12639 16292 12643 16348
rect 12643 16292 12699 16348
rect 12699 16292 12703 16348
rect 12639 16288 12703 16292
rect 12719 16348 12783 16352
rect 12719 16292 12723 16348
rect 12723 16292 12779 16348
rect 12779 16292 12783 16348
rect 12719 16288 12783 16292
rect 16458 16348 16522 16352
rect 16458 16292 16462 16348
rect 16462 16292 16518 16348
rect 16518 16292 16522 16348
rect 16458 16288 16522 16292
rect 16538 16348 16602 16352
rect 16538 16292 16542 16348
rect 16542 16292 16598 16348
rect 16598 16292 16602 16348
rect 16538 16288 16602 16292
rect 16618 16348 16682 16352
rect 16618 16292 16622 16348
rect 16622 16292 16678 16348
rect 16678 16292 16682 16348
rect 16618 16288 16682 16292
rect 16698 16348 16762 16352
rect 16698 16292 16702 16348
rect 16702 16292 16758 16348
rect 16758 16292 16762 16348
rect 16698 16288 16762 16292
rect 3861 15804 3925 15808
rect 3861 15748 3865 15804
rect 3865 15748 3921 15804
rect 3921 15748 3925 15804
rect 3861 15744 3925 15748
rect 3941 15804 4005 15808
rect 3941 15748 3945 15804
rect 3945 15748 4001 15804
rect 4001 15748 4005 15804
rect 3941 15744 4005 15748
rect 4021 15804 4085 15808
rect 4021 15748 4025 15804
rect 4025 15748 4081 15804
rect 4081 15748 4085 15804
rect 4021 15744 4085 15748
rect 4101 15804 4165 15808
rect 4101 15748 4105 15804
rect 4105 15748 4161 15804
rect 4161 15748 4165 15804
rect 4101 15744 4165 15748
rect 7840 15804 7904 15808
rect 7840 15748 7844 15804
rect 7844 15748 7900 15804
rect 7900 15748 7904 15804
rect 7840 15744 7904 15748
rect 7920 15804 7984 15808
rect 7920 15748 7924 15804
rect 7924 15748 7980 15804
rect 7980 15748 7984 15804
rect 7920 15744 7984 15748
rect 8000 15804 8064 15808
rect 8000 15748 8004 15804
rect 8004 15748 8060 15804
rect 8060 15748 8064 15804
rect 8000 15744 8064 15748
rect 8080 15804 8144 15808
rect 8080 15748 8084 15804
rect 8084 15748 8140 15804
rect 8140 15748 8144 15804
rect 8080 15744 8144 15748
rect 11819 15804 11883 15808
rect 11819 15748 11823 15804
rect 11823 15748 11879 15804
rect 11879 15748 11883 15804
rect 11819 15744 11883 15748
rect 11899 15804 11963 15808
rect 11899 15748 11903 15804
rect 11903 15748 11959 15804
rect 11959 15748 11963 15804
rect 11899 15744 11963 15748
rect 11979 15804 12043 15808
rect 11979 15748 11983 15804
rect 11983 15748 12039 15804
rect 12039 15748 12043 15804
rect 11979 15744 12043 15748
rect 12059 15804 12123 15808
rect 12059 15748 12063 15804
rect 12063 15748 12119 15804
rect 12119 15748 12123 15804
rect 12059 15744 12123 15748
rect 15798 15804 15862 15808
rect 15798 15748 15802 15804
rect 15802 15748 15858 15804
rect 15858 15748 15862 15804
rect 15798 15744 15862 15748
rect 15878 15804 15942 15808
rect 15878 15748 15882 15804
rect 15882 15748 15938 15804
rect 15938 15748 15942 15804
rect 15878 15744 15942 15748
rect 15958 15804 16022 15808
rect 15958 15748 15962 15804
rect 15962 15748 16018 15804
rect 16018 15748 16022 15804
rect 15958 15744 16022 15748
rect 16038 15804 16102 15808
rect 16038 15748 16042 15804
rect 16042 15748 16098 15804
rect 16098 15748 16102 15804
rect 16038 15744 16102 15748
rect 4521 15260 4585 15264
rect 4521 15204 4525 15260
rect 4525 15204 4581 15260
rect 4581 15204 4585 15260
rect 4521 15200 4585 15204
rect 4601 15260 4665 15264
rect 4601 15204 4605 15260
rect 4605 15204 4661 15260
rect 4661 15204 4665 15260
rect 4601 15200 4665 15204
rect 4681 15260 4745 15264
rect 4681 15204 4685 15260
rect 4685 15204 4741 15260
rect 4741 15204 4745 15260
rect 4681 15200 4745 15204
rect 4761 15260 4825 15264
rect 4761 15204 4765 15260
rect 4765 15204 4821 15260
rect 4821 15204 4825 15260
rect 4761 15200 4825 15204
rect 8500 15260 8564 15264
rect 8500 15204 8504 15260
rect 8504 15204 8560 15260
rect 8560 15204 8564 15260
rect 8500 15200 8564 15204
rect 8580 15260 8644 15264
rect 8580 15204 8584 15260
rect 8584 15204 8640 15260
rect 8640 15204 8644 15260
rect 8580 15200 8644 15204
rect 8660 15260 8724 15264
rect 8660 15204 8664 15260
rect 8664 15204 8720 15260
rect 8720 15204 8724 15260
rect 8660 15200 8724 15204
rect 8740 15260 8804 15264
rect 8740 15204 8744 15260
rect 8744 15204 8800 15260
rect 8800 15204 8804 15260
rect 8740 15200 8804 15204
rect 12479 15260 12543 15264
rect 12479 15204 12483 15260
rect 12483 15204 12539 15260
rect 12539 15204 12543 15260
rect 12479 15200 12543 15204
rect 12559 15260 12623 15264
rect 12559 15204 12563 15260
rect 12563 15204 12619 15260
rect 12619 15204 12623 15260
rect 12559 15200 12623 15204
rect 12639 15260 12703 15264
rect 12639 15204 12643 15260
rect 12643 15204 12699 15260
rect 12699 15204 12703 15260
rect 12639 15200 12703 15204
rect 12719 15260 12783 15264
rect 12719 15204 12723 15260
rect 12723 15204 12779 15260
rect 12779 15204 12783 15260
rect 12719 15200 12783 15204
rect 16458 15260 16522 15264
rect 16458 15204 16462 15260
rect 16462 15204 16518 15260
rect 16518 15204 16522 15260
rect 16458 15200 16522 15204
rect 16538 15260 16602 15264
rect 16538 15204 16542 15260
rect 16542 15204 16598 15260
rect 16598 15204 16602 15260
rect 16538 15200 16602 15204
rect 16618 15260 16682 15264
rect 16618 15204 16622 15260
rect 16622 15204 16678 15260
rect 16678 15204 16682 15260
rect 16618 15200 16682 15204
rect 16698 15260 16762 15264
rect 16698 15204 16702 15260
rect 16702 15204 16758 15260
rect 16758 15204 16762 15260
rect 16698 15200 16762 15204
rect 3861 14716 3925 14720
rect 3861 14660 3865 14716
rect 3865 14660 3921 14716
rect 3921 14660 3925 14716
rect 3861 14656 3925 14660
rect 3941 14716 4005 14720
rect 3941 14660 3945 14716
rect 3945 14660 4001 14716
rect 4001 14660 4005 14716
rect 3941 14656 4005 14660
rect 4021 14716 4085 14720
rect 4021 14660 4025 14716
rect 4025 14660 4081 14716
rect 4081 14660 4085 14716
rect 4021 14656 4085 14660
rect 4101 14716 4165 14720
rect 4101 14660 4105 14716
rect 4105 14660 4161 14716
rect 4161 14660 4165 14716
rect 4101 14656 4165 14660
rect 7840 14716 7904 14720
rect 7840 14660 7844 14716
rect 7844 14660 7900 14716
rect 7900 14660 7904 14716
rect 7840 14656 7904 14660
rect 7920 14716 7984 14720
rect 7920 14660 7924 14716
rect 7924 14660 7980 14716
rect 7980 14660 7984 14716
rect 7920 14656 7984 14660
rect 8000 14716 8064 14720
rect 8000 14660 8004 14716
rect 8004 14660 8060 14716
rect 8060 14660 8064 14716
rect 8000 14656 8064 14660
rect 8080 14716 8144 14720
rect 8080 14660 8084 14716
rect 8084 14660 8140 14716
rect 8140 14660 8144 14716
rect 8080 14656 8144 14660
rect 11819 14716 11883 14720
rect 11819 14660 11823 14716
rect 11823 14660 11879 14716
rect 11879 14660 11883 14716
rect 11819 14656 11883 14660
rect 11899 14716 11963 14720
rect 11899 14660 11903 14716
rect 11903 14660 11959 14716
rect 11959 14660 11963 14716
rect 11899 14656 11963 14660
rect 11979 14716 12043 14720
rect 11979 14660 11983 14716
rect 11983 14660 12039 14716
rect 12039 14660 12043 14716
rect 11979 14656 12043 14660
rect 12059 14716 12123 14720
rect 12059 14660 12063 14716
rect 12063 14660 12119 14716
rect 12119 14660 12123 14716
rect 12059 14656 12123 14660
rect 15798 14716 15862 14720
rect 15798 14660 15802 14716
rect 15802 14660 15858 14716
rect 15858 14660 15862 14716
rect 15798 14656 15862 14660
rect 15878 14716 15942 14720
rect 15878 14660 15882 14716
rect 15882 14660 15938 14716
rect 15938 14660 15942 14716
rect 15878 14656 15942 14660
rect 15958 14716 16022 14720
rect 15958 14660 15962 14716
rect 15962 14660 16018 14716
rect 16018 14660 16022 14716
rect 15958 14656 16022 14660
rect 16038 14716 16102 14720
rect 16038 14660 16042 14716
rect 16042 14660 16098 14716
rect 16098 14660 16102 14716
rect 16038 14656 16102 14660
rect 4521 14172 4585 14176
rect 4521 14116 4525 14172
rect 4525 14116 4581 14172
rect 4581 14116 4585 14172
rect 4521 14112 4585 14116
rect 4601 14172 4665 14176
rect 4601 14116 4605 14172
rect 4605 14116 4661 14172
rect 4661 14116 4665 14172
rect 4601 14112 4665 14116
rect 4681 14172 4745 14176
rect 4681 14116 4685 14172
rect 4685 14116 4741 14172
rect 4741 14116 4745 14172
rect 4681 14112 4745 14116
rect 4761 14172 4825 14176
rect 4761 14116 4765 14172
rect 4765 14116 4821 14172
rect 4821 14116 4825 14172
rect 4761 14112 4825 14116
rect 8500 14172 8564 14176
rect 8500 14116 8504 14172
rect 8504 14116 8560 14172
rect 8560 14116 8564 14172
rect 8500 14112 8564 14116
rect 8580 14172 8644 14176
rect 8580 14116 8584 14172
rect 8584 14116 8640 14172
rect 8640 14116 8644 14172
rect 8580 14112 8644 14116
rect 8660 14172 8724 14176
rect 8660 14116 8664 14172
rect 8664 14116 8720 14172
rect 8720 14116 8724 14172
rect 8660 14112 8724 14116
rect 8740 14172 8804 14176
rect 8740 14116 8744 14172
rect 8744 14116 8800 14172
rect 8800 14116 8804 14172
rect 8740 14112 8804 14116
rect 12479 14172 12543 14176
rect 12479 14116 12483 14172
rect 12483 14116 12539 14172
rect 12539 14116 12543 14172
rect 12479 14112 12543 14116
rect 12559 14172 12623 14176
rect 12559 14116 12563 14172
rect 12563 14116 12619 14172
rect 12619 14116 12623 14172
rect 12559 14112 12623 14116
rect 12639 14172 12703 14176
rect 12639 14116 12643 14172
rect 12643 14116 12699 14172
rect 12699 14116 12703 14172
rect 12639 14112 12703 14116
rect 12719 14172 12783 14176
rect 12719 14116 12723 14172
rect 12723 14116 12779 14172
rect 12779 14116 12783 14172
rect 12719 14112 12783 14116
rect 16458 14172 16522 14176
rect 16458 14116 16462 14172
rect 16462 14116 16518 14172
rect 16518 14116 16522 14172
rect 16458 14112 16522 14116
rect 16538 14172 16602 14176
rect 16538 14116 16542 14172
rect 16542 14116 16598 14172
rect 16598 14116 16602 14172
rect 16538 14112 16602 14116
rect 16618 14172 16682 14176
rect 16618 14116 16622 14172
rect 16622 14116 16678 14172
rect 16678 14116 16682 14172
rect 16618 14112 16682 14116
rect 16698 14172 16762 14176
rect 16698 14116 16702 14172
rect 16702 14116 16758 14172
rect 16758 14116 16762 14172
rect 16698 14112 16762 14116
rect 3861 13628 3925 13632
rect 3861 13572 3865 13628
rect 3865 13572 3921 13628
rect 3921 13572 3925 13628
rect 3861 13568 3925 13572
rect 3941 13628 4005 13632
rect 3941 13572 3945 13628
rect 3945 13572 4001 13628
rect 4001 13572 4005 13628
rect 3941 13568 4005 13572
rect 4021 13628 4085 13632
rect 4021 13572 4025 13628
rect 4025 13572 4081 13628
rect 4081 13572 4085 13628
rect 4021 13568 4085 13572
rect 4101 13628 4165 13632
rect 4101 13572 4105 13628
rect 4105 13572 4161 13628
rect 4161 13572 4165 13628
rect 4101 13568 4165 13572
rect 7840 13628 7904 13632
rect 7840 13572 7844 13628
rect 7844 13572 7900 13628
rect 7900 13572 7904 13628
rect 7840 13568 7904 13572
rect 7920 13628 7984 13632
rect 7920 13572 7924 13628
rect 7924 13572 7980 13628
rect 7980 13572 7984 13628
rect 7920 13568 7984 13572
rect 8000 13628 8064 13632
rect 8000 13572 8004 13628
rect 8004 13572 8060 13628
rect 8060 13572 8064 13628
rect 8000 13568 8064 13572
rect 8080 13628 8144 13632
rect 8080 13572 8084 13628
rect 8084 13572 8140 13628
rect 8140 13572 8144 13628
rect 8080 13568 8144 13572
rect 11819 13628 11883 13632
rect 11819 13572 11823 13628
rect 11823 13572 11879 13628
rect 11879 13572 11883 13628
rect 11819 13568 11883 13572
rect 11899 13628 11963 13632
rect 11899 13572 11903 13628
rect 11903 13572 11959 13628
rect 11959 13572 11963 13628
rect 11899 13568 11963 13572
rect 11979 13628 12043 13632
rect 11979 13572 11983 13628
rect 11983 13572 12039 13628
rect 12039 13572 12043 13628
rect 11979 13568 12043 13572
rect 12059 13628 12123 13632
rect 12059 13572 12063 13628
rect 12063 13572 12119 13628
rect 12119 13572 12123 13628
rect 12059 13568 12123 13572
rect 15798 13628 15862 13632
rect 15798 13572 15802 13628
rect 15802 13572 15858 13628
rect 15858 13572 15862 13628
rect 15798 13568 15862 13572
rect 15878 13628 15942 13632
rect 15878 13572 15882 13628
rect 15882 13572 15938 13628
rect 15938 13572 15942 13628
rect 15878 13568 15942 13572
rect 15958 13628 16022 13632
rect 15958 13572 15962 13628
rect 15962 13572 16018 13628
rect 16018 13572 16022 13628
rect 15958 13568 16022 13572
rect 16038 13628 16102 13632
rect 16038 13572 16042 13628
rect 16042 13572 16098 13628
rect 16098 13572 16102 13628
rect 16038 13568 16102 13572
rect 4521 13084 4585 13088
rect 4521 13028 4525 13084
rect 4525 13028 4581 13084
rect 4581 13028 4585 13084
rect 4521 13024 4585 13028
rect 4601 13084 4665 13088
rect 4601 13028 4605 13084
rect 4605 13028 4661 13084
rect 4661 13028 4665 13084
rect 4601 13024 4665 13028
rect 4681 13084 4745 13088
rect 4681 13028 4685 13084
rect 4685 13028 4741 13084
rect 4741 13028 4745 13084
rect 4681 13024 4745 13028
rect 4761 13084 4825 13088
rect 4761 13028 4765 13084
rect 4765 13028 4821 13084
rect 4821 13028 4825 13084
rect 4761 13024 4825 13028
rect 8500 13084 8564 13088
rect 8500 13028 8504 13084
rect 8504 13028 8560 13084
rect 8560 13028 8564 13084
rect 8500 13024 8564 13028
rect 8580 13084 8644 13088
rect 8580 13028 8584 13084
rect 8584 13028 8640 13084
rect 8640 13028 8644 13084
rect 8580 13024 8644 13028
rect 8660 13084 8724 13088
rect 8660 13028 8664 13084
rect 8664 13028 8720 13084
rect 8720 13028 8724 13084
rect 8660 13024 8724 13028
rect 8740 13084 8804 13088
rect 8740 13028 8744 13084
rect 8744 13028 8800 13084
rect 8800 13028 8804 13084
rect 8740 13024 8804 13028
rect 12479 13084 12543 13088
rect 12479 13028 12483 13084
rect 12483 13028 12539 13084
rect 12539 13028 12543 13084
rect 12479 13024 12543 13028
rect 12559 13084 12623 13088
rect 12559 13028 12563 13084
rect 12563 13028 12619 13084
rect 12619 13028 12623 13084
rect 12559 13024 12623 13028
rect 12639 13084 12703 13088
rect 12639 13028 12643 13084
rect 12643 13028 12699 13084
rect 12699 13028 12703 13084
rect 12639 13024 12703 13028
rect 12719 13084 12783 13088
rect 12719 13028 12723 13084
rect 12723 13028 12779 13084
rect 12779 13028 12783 13084
rect 12719 13024 12783 13028
rect 16458 13084 16522 13088
rect 16458 13028 16462 13084
rect 16462 13028 16518 13084
rect 16518 13028 16522 13084
rect 16458 13024 16522 13028
rect 16538 13084 16602 13088
rect 16538 13028 16542 13084
rect 16542 13028 16598 13084
rect 16598 13028 16602 13084
rect 16538 13024 16602 13028
rect 16618 13084 16682 13088
rect 16618 13028 16622 13084
rect 16622 13028 16678 13084
rect 16678 13028 16682 13084
rect 16618 13024 16682 13028
rect 16698 13084 16762 13088
rect 16698 13028 16702 13084
rect 16702 13028 16758 13084
rect 16758 13028 16762 13084
rect 16698 13024 16762 13028
rect 3861 12540 3925 12544
rect 3861 12484 3865 12540
rect 3865 12484 3921 12540
rect 3921 12484 3925 12540
rect 3861 12480 3925 12484
rect 3941 12540 4005 12544
rect 3941 12484 3945 12540
rect 3945 12484 4001 12540
rect 4001 12484 4005 12540
rect 3941 12480 4005 12484
rect 4021 12540 4085 12544
rect 4021 12484 4025 12540
rect 4025 12484 4081 12540
rect 4081 12484 4085 12540
rect 4021 12480 4085 12484
rect 4101 12540 4165 12544
rect 4101 12484 4105 12540
rect 4105 12484 4161 12540
rect 4161 12484 4165 12540
rect 4101 12480 4165 12484
rect 7840 12540 7904 12544
rect 7840 12484 7844 12540
rect 7844 12484 7900 12540
rect 7900 12484 7904 12540
rect 7840 12480 7904 12484
rect 7920 12540 7984 12544
rect 7920 12484 7924 12540
rect 7924 12484 7980 12540
rect 7980 12484 7984 12540
rect 7920 12480 7984 12484
rect 8000 12540 8064 12544
rect 8000 12484 8004 12540
rect 8004 12484 8060 12540
rect 8060 12484 8064 12540
rect 8000 12480 8064 12484
rect 8080 12540 8144 12544
rect 8080 12484 8084 12540
rect 8084 12484 8140 12540
rect 8140 12484 8144 12540
rect 8080 12480 8144 12484
rect 11819 12540 11883 12544
rect 11819 12484 11823 12540
rect 11823 12484 11879 12540
rect 11879 12484 11883 12540
rect 11819 12480 11883 12484
rect 11899 12540 11963 12544
rect 11899 12484 11903 12540
rect 11903 12484 11959 12540
rect 11959 12484 11963 12540
rect 11899 12480 11963 12484
rect 11979 12540 12043 12544
rect 11979 12484 11983 12540
rect 11983 12484 12039 12540
rect 12039 12484 12043 12540
rect 11979 12480 12043 12484
rect 12059 12540 12123 12544
rect 12059 12484 12063 12540
rect 12063 12484 12119 12540
rect 12119 12484 12123 12540
rect 12059 12480 12123 12484
rect 15798 12540 15862 12544
rect 15798 12484 15802 12540
rect 15802 12484 15858 12540
rect 15858 12484 15862 12540
rect 15798 12480 15862 12484
rect 15878 12540 15942 12544
rect 15878 12484 15882 12540
rect 15882 12484 15938 12540
rect 15938 12484 15942 12540
rect 15878 12480 15942 12484
rect 15958 12540 16022 12544
rect 15958 12484 15962 12540
rect 15962 12484 16018 12540
rect 16018 12484 16022 12540
rect 15958 12480 16022 12484
rect 16038 12540 16102 12544
rect 16038 12484 16042 12540
rect 16042 12484 16098 12540
rect 16098 12484 16102 12540
rect 16038 12480 16102 12484
rect 4521 11996 4585 12000
rect 4521 11940 4525 11996
rect 4525 11940 4581 11996
rect 4581 11940 4585 11996
rect 4521 11936 4585 11940
rect 4601 11996 4665 12000
rect 4601 11940 4605 11996
rect 4605 11940 4661 11996
rect 4661 11940 4665 11996
rect 4601 11936 4665 11940
rect 4681 11996 4745 12000
rect 4681 11940 4685 11996
rect 4685 11940 4741 11996
rect 4741 11940 4745 11996
rect 4681 11936 4745 11940
rect 4761 11996 4825 12000
rect 4761 11940 4765 11996
rect 4765 11940 4821 11996
rect 4821 11940 4825 11996
rect 4761 11936 4825 11940
rect 8500 11996 8564 12000
rect 8500 11940 8504 11996
rect 8504 11940 8560 11996
rect 8560 11940 8564 11996
rect 8500 11936 8564 11940
rect 8580 11996 8644 12000
rect 8580 11940 8584 11996
rect 8584 11940 8640 11996
rect 8640 11940 8644 11996
rect 8580 11936 8644 11940
rect 8660 11996 8724 12000
rect 8660 11940 8664 11996
rect 8664 11940 8720 11996
rect 8720 11940 8724 11996
rect 8660 11936 8724 11940
rect 8740 11996 8804 12000
rect 8740 11940 8744 11996
rect 8744 11940 8800 11996
rect 8800 11940 8804 11996
rect 8740 11936 8804 11940
rect 12479 11996 12543 12000
rect 12479 11940 12483 11996
rect 12483 11940 12539 11996
rect 12539 11940 12543 11996
rect 12479 11936 12543 11940
rect 12559 11996 12623 12000
rect 12559 11940 12563 11996
rect 12563 11940 12619 11996
rect 12619 11940 12623 11996
rect 12559 11936 12623 11940
rect 12639 11996 12703 12000
rect 12639 11940 12643 11996
rect 12643 11940 12699 11996
rect 12699 11940 12703 11996
rect 12639 11936 12703 11940
rect 12719 11996 12783 12000
rect 12719 11940 12723 11996
rect 12723 11940 12779 11996
rect 12779 11940 12783 11996
rect 12719 11936 12783 11940
rect 16458 11996 16522 12000
rect 16458 11940 16462 11996
rect 16462 11940 16518 11996
rect 16518 11940 16522 11996
rect 16458 11936 16522 11940
rect 16538 11996 16602 12000
rect 16538 11940 16542 11996
rect 16542 11940 16598 11996
rect 16598 11940 16602 11996
rect 16538 11936 16602 11940
rect 16618 11996 16682 12000
rect 16618 11940 16622 11996
rect 16622 11940 16678 11996
rect 16678 11940 16682 11996
rect 16618 11936 16682 11940
rect 16698 11996 16762 12000
rect 16698 11940 16702 11996
rect 16702 11940 16758 11996
rect 16758 11940 16762 11996
rect 16698 11936 16762 11940
rect 3861 11452 3925 11456
rect 3861 11396 3865 11452
rect 3865 11396 3921 11452
rect 3921 11396 3925 11452
rect 3861 11392 3925 11396
rect 3941 11452 4005 11456
rect 3941 11396 3945 11452
rect 3945 11396 4001 11452
rect 4001 11396 4005 11452
rect 3941 11392 4005 11396
rect 4021 11452 4085 11456
rect 4021 11396 4025 11452
rect 4025 11396 4081 11452
rect 4081 11396 4085 11452
rect 4021 11392 4085 11396
rect 4101 11452 4165 11456
rect 4101 11396 4105 11452
rect 4105 11396 4161 11452
rect 4161 11396 4165 11452
rect 4101 11392 4165 11396
rect 7840 11452 7904 11456
rect 7840 11396 7844 11452
rect 7844 11396 7900 11452
rect 7900 11396 7904 11452
rect 7840 11392 7904 11396
rect 7920 11452 7984 11456
rect 7920 11396 7924 11452
rect 7924 11396 7980 11452
rect 7980 11396 7984 11452
rect 7920 11392 7984 11396
rect 8000 11452 8064 11456
rect 8000 11396 8004 11452
rect 8004 11396 8060 11452
rect 8060 11396 8064 11452
rect 8000 11392 8064 11396
rect 8080 11452 8144 11456
rect 8080 11396 8084 11452
rect 8084 11396 8140 11452
rect 8140 11396 8144 11452
rect 8080 11392 8144 11396
rect 11819 11452 11883 11456
rect 11819 11396 11823 11452
rect 11823 11396 11879 11452
rect 11879 11396 11883 11452
rect 11819 11392 11883 11396
rect 11899 11452 11963 11456
rect 11899 11396 11903 11452
rect 11903 11396 11959 11452
rect 11959 11396 11963 11452
rect 11899 11392 11963 11396
rect 11979 11452 12043 11456
rect 11979 11396 11983 11452
rect 11983 11396 12039 11452
rect 12039 11396 12043 11452
rect 11979 11392 12043 11396
rect 12059 11452 12123 11456
rect 12059 11396 12063 11452
rect 12063 11396 12119 11452
rect 12119 11396 12123 11452
rect 12059 11392 12123 11396
rect 15798 11452 15862 11456
rect 15798 11396 15802 11452
rect 15802 11396 15858 11452
rect 15858 11396 15862 11452
rect 15798 11392 15862 11396
rect 15878 11452 15942 11456
rect 15878 11396 15882 11452
rect 15882 11396 15938 11452
rect 15938 11396 15942 11452
rect 15878 11392 15942 11396
rect 15958 11452 16022 11456
rect 15958 11396 15962 11452
rect 15962 11396 16018 11452
rect 16018 11396 16022 11452
rect 15958 11392 16022 11396
rect 16038 11452 16102 11456
rect 16038 11396 16042 11452
rect 16042 11396 16098 11452
rect 16098 11396 16102 11452
rect 16038 11392 16102 11396
rect 4521 10908 4585 10912
rect 4521 10852 4525 10908
rect 4525 10852 4581 10908
rect 4581 10852 4585 10908
rect 4521 10848 4585 10852
rect 4601 10908 4665 10912
rect 4601 10852 4605 10908
rect 4605 10852 4661 10908
rect 4661 10852 4665 10908
rect 4601 10848 4665 10852
rect 4681 10908 4745 10912
rect 4681 10852 4685 10908
rect 4685 10852 4741 10908
rect 4741 10852 4745 10908
rect 4681 10848 4745 10852
rect 4761 10908 4825 10912
rect 4761 10852 4765 10908
rect 4765 10852 4821 10908
rect 4821 10852 4825 10908
rect 4761 10848 4825 10852
rect 8500 10908 8564 10912
rect 8500 10852 8504 10908
rect 8504 10852 8560 10908
rect 8560 10852 8564 10908
rect 8500 10848 8564 10852
rect 8580 10908 8644 10912
rect 8580 10852 8584 10908
rect 8584 10852 8640 10908
rect 8640 10852 8644 10908
rect 8580 10848 8644 10852
rect 8660 10908 8724 10912
rect 8660 10852 8664 10908
rect 8664 10852 8720 10908
rect 8720 10852 8724 10908
rect 8660 10848 8724 10852
rect 8740 10908 8804 10912
rect 8740 10852 8744 10908
rect 8744 10852 8800 10908
rect 8800 10852 8804 10908
rect 8740 10848 8804 10852
rect 12479 10908 12543 10912
rect 12479 10852 12483 10908
rect 12483 10852 12539 10908
rect 12539 10852 12543 10908
rect 12479 10848 12543 10852
rect 12559 10908 12623 10912
rect 12559 10852 12563 10908
rect 12563 10852 12619 10908
rect 12619 10852 12623 10908
rect 12559 10848 12623 10852
rect 12639 10908 12703 10912
rect 12639 10852 12643 10908
rect 12643 10852 12699 10908
rect 12699 10852 12703 10908
rect 12639 10848 12703 10852
rect 12719 10908 12783 10912
rect 12719 10852 12723 10908
rect 12723 10852 12779 10908
rect 12779 10852 12783 10908
rect 12719 10848 12783 10852
rect 16458 10908 16522 10912
rect 16458 10852 16462 10908
rect 16462 10852 16518 10908
rect 16518 10852 16522 10908
rect 16458 10848 16522 10852
rect 16538 10908 16602 10912
rect 16538 10852 16542 10908
rect 16542 10852 16598 10908
rect 16598 10852 16602 10908
rect 16538 10848 16602 10852
rect 16618 10908 16682 10912
rect 16618 10852 16622 10908
rect 16622 10852 16678 10908
rect 16678 10852 16682 10908
rect 16618 10848 16682 10852
rect 16698 10908 16762 10912
rect 16698 10852 16702 10908
rect 16702 10852 16758 10908
rect 16758 10852 16762 10908
rect 16698 10848 16762 10852
rect 3861 10364 3925 10368
rect 3861 10308 3865 10364
rect 3865 10308 3921 10364
rect 3921 10308 3925 10364
rect 3861 10304 3925 10308
rect 3941 10364 4005 10368
rect 3941 10308 3945 10364
rect 3945 10308 4001 10364
rect 4001 10308 4005 10364
rect 3941 10304 4005 10308
rect 4021 10364 4085 10368
rect 4021 10308 4025 10364
rect 4025 10308 4081 10364
rect 4081 10308 4085 10364
rect 4021 10304 4085 10308
rect 4101 10364 4165 10368
rect 4101 10308 4105 10364
rect 4105 10308 4161 10364
rect 4161 10308 4165 10364
rect 4101 10304 4165 10308
rect 7840 10364 7904 10368
rect 7840 10308 7844 10364
rect 7844 10308 7900 10364
rect 7900 10308 7904 10364
rect 7840 10304 7904 10308
rect 7920 10364 7984 10368
rect 7920 10308 7924 10364
rect 7924 10308 7980 10364
rect 7980 10308 7984 10364
rect 7920 10304 7984 10308
rect 8000 10364 8064 10368
rect 8000 10308 8004 10364
rect 8004 10308 8060 10364
rect 8060 10308 8064 10364
rect 8000 10304 8064 10308
rect 8080 10364 8144 10368
rect 8080 10308 8084 10364
rect 8084 10308 8140 10364
rect 8140 10308 8144 10364
rect 8080 10304 8144 10308
rect 11819 10364 11883 10368
rect 11819 10308 11823 10364
rect 11823 10308 11879 10364
rect 11879 10308 11883 10364
rect 11819 10304 11883 10308
rect 11899 10364 11963 10368
rect 11899 10308 11903 10364
rect 11903 10308 11959 10364
rect 11959 10308 11963 10364
rect 11899 10304 11963 10308
rect 11979 10364 12043 10368
rect 11979 10308 11983 10364
rect 11983 10308 12039 10364
rect 12039 10308 12043 10364
rect 11979 10304 12043 10308
rect 12059 10364 12123 10368
rect 12059 10308 12063 10364
rect 12063 10308 12119 10364
rect 12119 10308 12123 10364
rect 12059 10304 12123 10308
rect 15798 10364 15862 10368
rect 15798 10308 15802 10364
rect 15802 10308 15858 10364
rect 15858 10308 15862 10364
rect 15798 10304 15862 10308
rect 15878 10364 15942 10368
rect 15878 10308 15882 10364
rect 15882 10308 15938 10364
rect 15938 10308 15942 10364
rect 15878 10304 15942 10308
rect 15958 10364 16022 10368
rect 15958 10308 15962 10364
rect 15962 10308 16018 10364
rect 16018 10308 16022 10364
rect 15958 10304 16022 10308
rect 16038 10364 16102 10368
rect 16038 10308 16042 10364
rect 16042 10308 16098 10364
rect 16098 10308 16102 10364
rect 16038 10304 16102 10308
rect 4521 9820 4585 9824
rect 4521 9764 4525 9820
rect 4525 9764 4581 9820
rect 4581 9764 4585 9820
rect 4521 9760 4585 9764
rect 4601 9820 4665 9824
rect 4601 9764 4605 9820
rect 4605 9764 4661 9820
rect 4661 9764 4665 9820
rect 4601 9760 4665 9764
rect 4681 9820 4745 9824
rect 4681 9764 4685 9820
rect 4685 9764 4741 9820
rect 4741 9764 4745 9820
rect 4681 9760 4745 9764
rect 4761 9820 4825 9824
rect 4761 9764 4765 9820
rect 4765 9764 4821 9820
rect 4821 9764 4825 9820
rect 4761 9760 4825 9764
rect 8500 9820 8564 9824
rect 8500 9764 8504 9820
rect 8504 9764 8560 9820
rect 8560 9764 8564 9820
rect 8500 9760 8564 9764
rect 8580 9820 8644 9824
rect 8580 9764 8584 9820
rect 8584 9764 8640 9820
rect 8640 9764 8644 9820
rect 8580 9760 8644 9764
rect 8660 9820 8724 9824
rect 8660 9764 8664 9820
rect 8664 9764 8720 9820
rect 8720 9764 8724 9820
rect 8660 9760 8724 9764
rect 8740 9820 8804 9824
rect 8740 9764 8744 9820
rect 8744 9764 8800 9820
rect 8800 9764 8804 9820
rect 8740 9760 8804 9764
rect 12479 9820 12543 9824
rect 12479 9764 12483 9820
rect 12483 9764 12539 9820
rect 12539 9764 12543 9820
rect 12479 9760 12543 9764
rect 12559 9820 12623 9824
rect 12559 9764 12563 9820
rect 12563 9764 12619 9820
rect 12619 9764 12623 9820
rect 12559 9760 12623 9764
rect 12639 9820 12703 9824
rect 12639 9764 12643 9820
rect 12643 9764 12699 9820
rect 12699 9764 12703 9820
rect 12639 9760 12703 9764
rect 12719 9820 12783 9824
rect 12719 9764 12723 9820
rect 12723 9764 12779 9820
rect 12779 9764 12783 9820
rect 12719 9760 12783 9764
rect 16458 9820 16522 9824
rect 16458 9764 16462 9820
rect 16462 9764 16518 9820
rect 16518 9764 16522 9820
rect 16458 9760 16522 9764
rect 16538 9820 16602 9824
rect 16538 9764 16542 9820
rect 16542 9764 16598 9820
rect 16598 9764 16602 9820
rect 16538 9760 16602 9764
rect 16618 9820 16682 9824
rect 16618 9764 16622 9820
rect 16622 9764 16678 9820
rect 16678 9764 16682 9820
rect 16618 9760 16682 9764
rect 16698 9820 16762 9824
rect 16698 9764 16702 9820
rect 16702 9764 16758 9820
rect 16758 9764 16762 9820
rect 16698 9760 16762 9764
rect 3861 9276 3925 9280
rect 3861 9220 3865 9276
rect 3865 9220 3921 9276
rect 3921 9220 3925 9276
rect 3861 9216 3925 9220
rect 3941 9276 4005 9280
rect 3941 9220 3945 9276
rect 3945 9220 4001 9276
rect 4001 9220 4005 9276
rect 3941 9216 4005 9220
rect 4021 9276 4085 9280
rect 4021 9220 4025 9276
rect 4025 9220 4081 9276
rect 4081 9220 4085 9276
rect 4021 9216 4085 9220
rect 4101 9276 4165 9280
rect 4101 9220 4105 9276
rect 4105 9220 4161 9276
rect 4161 9220 4165 9276
rect 4101 9216 4165 9220
rect 7840 9276 7904 9280
rect 7840 9220 7844 9276
rect 7844 9220 7900 9276
rect 7900 9220 7904 9276
rect 7840 9216 7904 9220
rect 7920 9276 7984 9280
rect 7920 9220 7924 9276
rect 7924 9220 7980 9276
rect 7980 9220 7984 9276
rect 7920 9216 7984 9220
rect 8000 9276 8064 9280
rect 8000 9220 8004 9276
rect 8004 9220 8060 9276
rect 8060 9220 8064 9276
rect 8000 9216 8064 9220
rect 8080 9276 8144 9280
rect 8080 9220 8084 9276
rect 8084 9220 8140 9276
rect 8140 9220 8144 9276
rect 8080 9216 8144 9220
rect 11819 9276 11883 9280
rect 11819 9220 11823 9276
rect 11823 9220 11879 9276
rect 11879 9220 11883 9276
rect 11819 9216 11883 9220
rect 11899 9276 11963 9280
rect 11899 9220 11903 9276
rect 11903 9220 11959 9276
rect 11959 9220 11963 9276
rect 11899 9216 11963 9220
rect 11979 9276 12043 9280
rect 11979 9220 11983 9276
rect 11983 9220 12039 9276
rect 12039 9220 12043 9276
rect 11979 9216 12043 9220
rect 12059 9276 12123 9280
rect 12059 9220 12063 9276
rect 12063 9220 12119 9276
rect 12119 9220 12123 9276
rect 12059 9216 12123 9220
rect 15798 9276 15862 9280
rect 15798 9220 15802 9276
rect 15802 9220 15858 9276
rect 15858 9220 15862 9276
rect 15798 9216 15862 9220
rect 15878 9276 15942 9280
rect 15878 9220 15882 9276
rect 15882 9220 15938 9276
rect 15938 9220 15942 9276
rect 15878 9216 15942 9220
rect 15958 9276 16022 9280
rect 15958 9220 15962 9276
rect 15962 9220 16018 9276
rect 16018 9220 16022 9276
rect 15958 9216 16022 9220
rect 16038 9276 16102 9280
rect 16038 9220 16042 9276
rect 16042 9220 16098 9276
rect 16098 9220 16102 9276
rect 16038 9216 16102 9220
rect 4521 8732 4585 8736
rect 4521 8676 4525 8732
rect 4525 8676 4581 8732
rect 4581 8676 4585 8732
rect 4521 8672 4585 8676
rect 4601 8732 4665 8736
rect 4601 8676 4605 8732
rect 4605 8676 4661 8732
rect 4661 8676 4665 8732
rect 4601 8672 4665 8676
rect 4681 8732 4745 8736
rect 4681 8676 4685 8732
rect 4685 8676 4741 8732
rect 4741 8676 4745 8732
rect 4681 8672 4745 8676
rect 4761 8732 4825 8736
rect 4761 8676 4765 8732
rect 4765 8676 4821 8732
rect 4821 8676 4825 8732
rect 4761 8672 4825 8676
rect 8500 8732 8564 8736
rect 8500 8676 8504 8732
rect 8504 8676 8560 8732
rect 8560 8676 8564 8732
rect 8500 8672 8564 8676
rect 8580 8732 8644 8736
rect 8580 8676 8584 8732
rect 8584 8676 8640 8732
rect 8640 8676 8644 8732
rect 8580 8672 8644 8676
rect 8660 8732 8724 8736
rect 8660 8676 8664 8732
rect 8664 8676 8720 8732
rect 8720 8676 8724 8732
rect 8660 8672 8724 8676
rect 8740 8732 8804 8736
rect 8740 8676 8744 8732
rect 8744 8676 8800 8732
rect 8800 8676 8804 8732
rect 8740 8672 8804 8676
rect 12479 8732 12543 8736
rect 12479 8676 12483 8732
rect 12483 8676 12539 8732
rect 12539 8676 12543 8732
rect 12479 8672 12543 8676
rect 12559 8732 12623 8736
rect 12559 8676 12563 8732
rect 12563 8676 12619 8732
rect 12619 8676 12623 8732
rect 12559 8672 12623 8676
rect 12639 8732 12703 8736
rect 12639 8676 12643 8732
rect 12643 8676 12699 8732
rect 12699 8676 12703 8732
rect 12639 8672 12703 8676
rect 12719 8732 12783 8736
rect 12719 8676 12723 8732
rect 12723 8676 12779 8732
rect 12779 8676 12783 8732
rect 12719 8672 12783 8676
rect 16458 8732 16522 8736
rect 16458 8676 16462 8732
rect 16462 8676 16518 8732
rect 16518 8676 16522 8732
rect 16458 8672 16522 8676
rect 16538 8732 16602 8736
rect 16538 8676 16542 8732
rect 16542 8676 16598 8732
rect 16598 8676 16602 8732
rect 16538 8672 16602 8676
rect 16618 8732 16682 8736
rect 16618 8676 16622 8732
rect 16622 8676 16678 8732
rect 16678 8676 16682 8732
rect 16618 8672 16682 8676
rect 16698 8732 16762 8736
rect 16698 8676 16702 8732
rect 16702 8676 16758 8732
rect 16758 8676 16762 8732
rect 16698 8672 16762 8676
rect 3861 8188 3925 8192
rect 3861 8132 3865 8188
rect 3865 8132 3921 8188
rect 3921 8132 3925 8188
rect 3861 8128 3925 8132
rect 3941 8188 4005 8192
rect 3941 8132 3945 8188
rect 3945 8132 4001 8188
rect 4001 8132 4005 8188
rect 3941 8128 4005 8132
rect 4021 8188 4085 8192
rect 4021 8132 4025 8188
rect 4025 8132 4081 8188
rect 4081 8132 4085 8188
rect 4021 8128 4085 8132
rect 4101 8188 4165 8192
rect 4101 8132 4105 8188
rect 4105 8132 4161 8188
rect 4161 8132 4165 8188
rect 4101 8128 4165 8132
rect 7840 8188 7904 8192
rect 7840 8132 7844 8188
rect 7844 8132 7900 8188
rect 7900 8132 7904 8188
rect 7840 8128 7904 8132
rect 7920 8188 7984 8192
rect 7920 8132 7924 8188
rect 7924 8132 7980 8188
rect 7980 8132 7984 8188
rect 7920 8128 7984 8132
rect 8000 8188 8064 8192
rect 8000 8132 8004 8188
rect 8004 8132 8060 8188
rect 8060 8132 8064 8188
rect 8000 8128 8064 8132
rect 8080 8188 8144 8192
rect 8080 8132 8084 8188
rect 8084 8132 8140 8188
rect 8140 8132 8144 8188
rect 8080 8128 8144 8132
rect 11819 8188 11883 8192
rect 11819 8132 11823 8188
rect 11823 8132 11879 8188
rect 11879 8132 11883 8188
rect 11819 8128 11883 8132
rect 11899 8188 11963 8192
rect 11899 8132 11903 8188
rect 11903 8132 11959 8188
rect 11959 8132 11963 8188
rect 11899 8128 11963 8132
rect 11979 8188 12043 8192
rect 11979 8132 11983 8188
rect 11983 8132 12039 8188
rect 12039 8132 12043 8188
rect 11979 8128 12043 8132
rect 12059 8188 12123 8192
rect 12059 8132 12063 8188
rect 12063 8132 12119 8188
rect 12119 8132 12123 8188
rect 12059 8128 12123 8132
rect 15798 8188 15862 8192
rect 15798 8132 15802 8188
rect 15802 8132 15858 8188
rect 15858 8132 15862 8188
rect 15798 8128 15862 8132
rect 15878 8188 15942 8192
rect 15878 8132 15882 8188
rect 15882 8132 15938 8188
rect 15938 8132 15942 8188
rect 15878 8128 15942 8132
rect 15958 8188 16022 8192
rect 15958 8132 15962 8188
rect 15962 8132 16018 8188
rect 16018 8132 16022 8188
rect 15958 8128 16022 8132
rect 16038 8188 16102 8192
rect 16038 8132 16042 8188
rect 16042 8132 16098 8188
rect 16098 8132 16102 8188
rect 16038 8128 16102 8132
rect 4521 7644 4585 7648
rect 4521 7588 4525 7644
rect 4525 7588 4581 7644
rect 4581 7588 4585 7644
rect 4521 7584 4585 7588
rect 4601 7644 4665 7648
rect 4601 7588 4605 7644
rect 4605 7588 4661 7644
rect 4661 7588 4665 7644
rect 4601 7584 4665 7588
rect 4681 7644 4745 7648
rect 4681 7588 4685 7644
rect 4685 7588 4741 7644
rect 4741 7588 4745 7644
rect 4681 7584 4745 7588
rect 4761 7644 4825 7648
rect 4761 7588 4765 7644
rect 4765 7588 4821 7644
rect 4821 7588 4825 7644
rect 4761 7584 4825 7588
rect 8500 7644 8564 7648
rect 8500 7588 8504 7644
rect 8504 7588 8560 7644
rect 8560 7588 8564 7644
rect 8500 7584 8564 7588
rect 8580 7644 8644 7648
rect 8580 7588 8584 7644
rect 8584 7588 8640 7644
rect 8640 7588 8644 7644
rect 8580 7584 8644 7588
rect 8660 7644 8724 7648
rect 8660 7588 8664 7644
rect 8664 7588 8720 7644
rect 8720 7588 8724 7644
rect 8660 7584 8724 7588
rect 8740 7644 8804 7648
rect 8740 7588 8744 7644
rect 8744 7588 8800 7644
rect 8800 7588 8804 7644
rect 8740 7584 8804 7588
rect 12479 7644 12543 7648
rect 12479 7588 12483 7644
rect 12483 7588 12539 7644
rect 12539 7588 12543 7644
rect 12479 7584 12543 7588
rect 12559 7644 12623 7648
rect 12559 7588 12563 7644
rect 12563 7588 12619 7644
rect 12619 7588 12623 7644
rect 12559 7584 12623 7588
rect 12639 7644 12703 7648
rect 12639 7588 12643 7644
rect 12643 7588 12699 7644
rect 12699 7588 12703 7644
rect 12639 7584 12703 7588
rect 12719 7644 12783 7648
rect 12719 7588 12723 7644
rect 12723 7588 12779 7644
rect 12779 7588 12783 7644
rect 12719 7584 12783 7588
rect 16458 7644 16522 7648
rect 16458 7588 16462 7644
rect 16462 7588 16518 7644
rect 16518 7588 16522 7644
rect 16458 7584 16522 7588
rect 16538 7644 16602 7648
rect 16538 7588 16542 7644
rect 16542 7588 16598 7644
rect 16598 7588 16602 7644
rect 16538 7584 16602 7588
rect 16618 7644 16682 7648
rect 16618 7588 16622 7644
rect 16622 7588 16678 7644
rect 16678 7588 16682 7644
rect 16618 7584 16682 7588
rect 16698 7644 16762 7648
rect 16698 7588 16702 7644
rect 16702 7588 16758 7644
rect 16758 7588 16762 7644
rect 16698 7584 16762 7588
rect 3861 7100 3925 7104
rect 3861 7044 3865 7100
rect 3865 7044 3921 7100
rect 3921 7044 3925 7100
rect 3861 7040 3925 7044
rect 3941 7100 4005 7104
rect 3941 7044 3945 7100
rect 3945 7044 4001 7100
rect 4001 7044 4005 7100
rect 3941 7040 4005 7044
rect 4021 7100 4085 7104
rect 4021 7044 4025 7100
rect 4025 7044 4081 7100
rect 4081 7044 4085 7100
rect 4021 7040 4085 7044
rect 4101 7100 4165 7104
rect 4101 7044 4105 7100
rect 4105 7044 4161 7100
rect 4161 7044 4165 7100
rect 4101 7040 4165 7044
rect 7840 7100 7904 7104
rect 7840 7044 7844 7100
rect 7844 7044 7900 7100
rect 7900 7044 7904 7100
rect 7840 7040 7904 7044
rect 7920 7100 7984 7104
rect 7920 7044 7924 7100
rect 7924 7044 7980 7100
rect 7980 7044 7984 7100
rect 7920 7040 7984 7044
rect 8000 7100 8064 7104
rect 8000 7044 8004 7100
rect 8004 7044 8060 7100
rect 8060 7044 8064 7100
rect 8000 7040 8064 7044
rect 8080 7100 8144 7104
rect 8080 7044 8084 7100
rect 8084 7044 8140 7100
rect 8140 7044 8144 7100
rect 8080 7040 8144 7044
rect 11819 7100 11883 7104
rect 11819 7044 11823 7100
rect 11823 7044 11879 7100
rect 11879 7044 11883 7100
rect 11819 7040 11883 7044
rect 11899 7100 11963 7104
rect 11899 7044 11903 7100
rect 11903 7044 11959 7100
rect 11959 7044 11963 7100
rect 11899 7040 11963 7044
rect 11979 7100 12043 7104
rect 11979 7044 11983 7100
rect 11983 7044 12039 7100
rect 12039 7044 12043 7100
rect 11979 7040 12043 7044
rect 12059 7100 12123 7104
rect 12059 7044 12063 7100
rect 12063 7044 12119 7100
rect 12119 7044 12123 7100
rect 12059 7040 12123 7044
rect 15798 7100 15862 7104
rect 15798 7044 15802 7100
rect 15802 7044 15858 7100
rect 15858 7044 15862 7100
rect 15798 7040 15862 7044
rect 15878 7100 15942 7104
rect 15878 7044 15882 7100
rect 15882 7044 15938 7100
rect 15938 7044 15942 7100
rect 15878 7040 15942 7044
rect 15958 7100 16022 7104
rect 15958 7044 15962 7100
rect 15962 7044 16018 7100
rect 16018 7044 16022 7100
rect 15958 7040 16022 7044
rect 16038 7100 16102 7104
rect 16038 7044 16042 7100
rect 16042 7044 16098 7100
rect 16098 7044 16102 7100
rect 16038 7040 16102 7044
rect 4521 6556 4585 6560
rect 4521 6500 4525 6556
rect 4525 6500 4581 6556
rect 4581 6500 4585 6556
rect 4521 6496 4585 6500
rect 4601 6556 4665 6560
rect 4601 6500 4605 6556
rect 4605 6500 4661 6556
rect 4661 6500 4665 6556
rect 4601 6496 4665 6500
rect 4681 6556 4745 6560
rect 4681 6500 4685 6556
rect 4685 6500 4741 6556
rect 4741 6500 4745 6556
rect 4681 6496 4745 6500
rect 4761 6556 4825 6560
rect 4761 6500 4765 6556
rect 4765 6500 4821 6556
rect 4821 6500 4825 6556
rect 4761 6496 4825 6500
rect 8500 6556 8564 6560
rect 8500 6500 8504 6556
rect 8504 6500 8560 6556
rect 8560 6500 8564 6556
rect 8500 6496 8564 6500
rect 8580 6556 8644 6560
rect 8580 6500 8584 6556
rect 8584 6500 8640 6556
rect 8640 6500 8644 6556
rect 8580 6496 8644 6500
rect 8660 6556 8724 6560
rect 8660 6500 8664 6556
rect 8664 6500 8720 6556
rect 8720 6500 8724 6556
rect 8660 6496 8724 6500
rect 8740 6556 8804 6560
rect 8740 6500 8744 6556
rect 8744 6500 8800 6556
rect 8800 6500 8804 6556
rect 8740 6496 8804 6500
rect 12479 6556 12543 6560
rect 12479 6500 12483 6556
rect 12483 6500 12539 6556
rect 12539 6500 12543 6556
rect 12479 6496 12543 6500
rect 12559 6556 12623 6560
rect 12559 6500 12563 6556
rect 12563 6500 12619 6556
rect 12619 6500 12623 6556
rect 12559 6496 12623 6500
rect 12639 6556 12703 6560
rect 12639 6500 12643 6556
rect 12643 6500 12699 6556
rect 12699 6500 12703 6556
rect 12639 6496 12703 6500
rect 12719 6556 12783 6560
rect 12719 6500 12723 6556
rect 12723 6500 12779 6556
rect 12779 6500 12783 6556
rect 12719 6496 12783 6500
rect 16458 6556 16522 6560
rect 16458 6500 16462 6556
rect 16462 6500 16518 6556
rect 16518 6500 16522 6556
rect 16458 6496 16522 6500
rect 16538 6556 16602 6560
rect 16538 6500 16542 6556
rect 16542 6500 16598 6556
rect 16598 6500 16602 6556
rect 16538 6496 16602 6500
rect 16618 6556 16682 6560
rect 16618 6500 16622 6556
rect 16622 6500 16678 6556
rect 16678 6500 16682 6556
rect 16618 6496 16682 6500
rect 16698 6556 16762 6560
rect 16698 6500 16702 6556
rect 16702 6500 16758 6556
rect 16758 6500 16762 6556
rect 16698 6496 16762 6500
rect 3861 6012 3925 6016
rect 3861 5956 3865 6012
rect 3865 5956 3921 6012
rect 3921 5956 3925 6012
rect 3861 5952 3925 5956
rect 3941 6012 4005 6016
rect 3941 5956 3945 6012
rect 3945 5956 4001 6012
rect 4001 5956 4005 6012
rect 3941 5952 4005 5956
rect 4021 6012 4085 6016
rect 4021 5956 4025 6012
rect 4025 5956 4081 6012
rect 4081 5956 4085 6012
rect 4021 5952 4085 5956
rect 4101 6012 4165 6016
rect 4101 5956 4105 6012
rect 4105 5956 4161 6012
rect 4161 5956 4165 6012
rect 4101 5952 4165 5956
rect 7840 6012 7904 6016
rect 7840 5956 7844 6012
rect 7844 5956 7900 6012
rect 7900 5956 7904 6012
rect 7840 5952 7904 5956
rect 7920 6012 7984 6016
rect 7920 5956 7924 6012
rect 7924 5956 7980 6012
rect 7980 5956 7984 6012
rect 7920 5952 7984 5956
rect 8000 6012 8064 6016
rect 8000 5956 8004 6012
rect 8004 5956 8060 6012
rect 8060 5956 8064 6012
rect 8000 5952 8064 5956
rect 8080 6012 8144 6016
rect 8080 5956 8084 6012
rect 8084 5956 8140 6012
rect 8140 5956 8144 6012
rect 8080 5952 8144 5956
rect 11819 6012 11883 6016
rect 11819 5956 11823 6012
rect 11823 5956 11879 6012
rect 11879 5956 11883 6012
rect 11819 5952 11883 5956
rect 11899 6012 11963 6016
rect 11899 5956 11903 6012
rect 11903 5956 11959 6012
rect 11959 5956 11963 6012
rect 11899 5952 11963 5956
rect 11979 6012 12043 6016
rect 11979 5956 11983 6012
rect 11983 5956 12039 6012
rect 12039 5956 12043 6012
rect 11979 5952 12043 5956
rect 12059 6012 12123 6016
rect 12059 5956 12063 6012
rect 12063 5956 12119 6012
rect 12119 5956 12123 6012
rect 12059 5952 12123 5956
rect 15798 6012 15862 6016
rect 15798 5956 15802 6012
rect 15802 5956 15858 6012
rect 15858 5956 15862 6012
rect 15798 5952 15862 5956
rect 15878 6012 15942 6016
rect 15878 5956 15882 6012
rect 15882 5956 15938 6012
rect 15938 5956 15942 6012
rect 15878 5952 15942 5956
rect 15958 6012 16022 6016
rect 15958 5956 15962 6012
rect 15962 5956 16018 6012
rect 16018 5956 16022 6012
rect 15958 5952 16022 5956
rect 16038 6012 16102 6016
rect 16038 5956 16042 6012
rect 16042 5956 16098 6012
rect 16098 5956 16102 6012
rect 16038 5952 16102 5956
rect 4521 5468 4585 5472
rect 4521 5412 4525 5468
rect 4525 5412 4581 5468
rect 4581 5412 4585 5468
rect 4521 5408 4585 5412
rect 4601 5468 4665 5472
rect 4601 5412 4605 5468
rect 4605 5412 4661 5468
rect 4661 5412 4665 5468
rect 4601 5408 4665 5412
rect 4681 5468 4745 5472
rect 4681 5412 4685 5468
rect 4685 5412 4741 5468
rect 4741 5412 4745 5468
rect 4681 5408 4745 5412
rect 4761 5468 4825 5472
rect 4761 5412 4765 5468
rect 4765 5412 4821 5468
rect 4821 5412 4825 5468
rect 4761 5408 4825 5412
rect 8500 5468 8564 5472
rect 8500 5412 8504 5468
rect 8504 5412 8560 5468
rect 8560 5412 8564 5468
rect 8500 5408 8564 5412
rect 8580 5468 8644 5472
rect 8580 5412 8584 5468
rect 8584 5412 8640 5468
rect 8640 5412 8644 5468
rect 8580 5408 8644 5412
rect 8660 5468 8724 5472
rect 8660 5412 8664 5468
rect 8664 5412 8720 5468
rect 8720 5412 8724 5468
rect 8660 5408 8724 5412
rect 8740 5468 8804 5472
rect 8740 5412 8744 5468
rect 8744 5412 8800 5468
rect 8800 5412 8804 5468
rect 8740 5408 8804 5412
rect 12479 5468 12543 5472
rect 12479 5412 12483 5468
rect 12483 5412 12539 5468
rect 12539 5412 12543 5468
rect 12479 5408 12543 5412
rect 12559 5468 12623 5472
rect 12559 5412 12563 5468
rect 12563 5412 12619 5468
rect 12619 5412 12623 5468
rect 12559 5408 12623 5412
rect 12639 5468 12703 5472
rect 12639 5412 12643 5468
rect 12643 5412 12699 5468
rect 12699 5412 12703 5468
rect 12639 5408 12703 5412
rect 12719 5468 12783 5472
rect 12719 5412 12723 5468
rect 12723 5412 12779 5468
rect 12779 5412 12783 5468
rect 12719 5408 12783 5412
rect 16458 5468 16522 5472
rect 16458 5412 16462 5468
rect 16462 5412 16518 5468
rect 16518 5412 16522 5468
rect 16458 5408 16522 5412
rect 16538 5468 16602 5472
rect 16538 5412 16542 5468
rect 16542 5412 16598 5468
rect 16598 5412 16602 5468
rect 16538 5408 16602 5412
rect 16618 5468 16682 5472
rect 16618 5412 16622 5468
rect 16622 5412 16678 5468
rect 16678 5412 16682 5468
rect 16618 5408 16682 5412
rect 16698 5468 16762 5472
rect 16698 5412 16702 5468
rect 16702 5412 16758 5468
rect 16758 5412 16762 5468
rect 16698 5408 16762 5412
rect 3861 4924 3925 4928
rect 3861 4868 3865 4924
rect 3865 4868 3921 4924
rect 3921 4868 3925 4924
rect 3861 4864 3925 4868
rect 3941 4924 4005 4928
rect 3941 4868 3945 4924
rect 3945 4868 4001 4924
rect 4001 4868 4005 4924
rect 3941 4864 4005 4868
rect 4021 4924 4085 4928
rect 4021 4868 4025 4924
rect 4025 4868 4081 4924
rect 4081 4868 4085 4924
rect 4021 4864 4085 4868
rect 4101 4924 4165 4928
rect 4101 4868 4105 4924
rect 4105 4868 4161 4924
rect 4161 4868 4165 4924
rect 4101 4864 4165 4868
rect 7840 4924 7904 4928
rect 7840 4868 7844 4924
rect 7844 4868 7900 4924
rect 7900 4868 7904 4924
rect 7840 4864 7904 4868
rect 7920 4924 7984 4928
rect 7920 4868 7924 4924
rect 7924 4868 7980 4924
rect 7980 4868 7984 4924
rect 7920 4864 7984 4868
rect 8000 4924 8064 4928
rect 8000 4868 8004 4924
rect 8004 4868 8060 4924
rect 8060 4868 8064 4924
rect 8000 4864 8064 4868
rect 8080 4924 8144 4928
rect 8080 4868 8084 4924
rect 8084 4868 8140 4924
rect 8140 4868 8144 4924
rect 8080 4864 8144 4868
rect 11819 4924 11883 4928
rect 11819 4868 11823 4924
rect 11823 4868 11879 4924
rect 11879 4868 11883 4924
rect 11819 4864 11883 4868
rect 11899 4924 11963 4928
rect 11899 4868 11903 4924
rect 11903 4868 11959 4924
rect 11959 4868 11963 4924
rect 11899 4864 11963 4868
rect 11979 4924 12043 4928
rect 11979 4868 11983 4924
rect 11983 4868 12039 4924
rect 12039 4868 12043 4924
rect 11979 4864 12043 4868
rect 12059 4924 12123 4928
rect 12059 4868 12063 4924
rect 12063 4868 12119 4924
rect 12119 4868 12123 4924
rect 12059 4864 12123 4868
rect 15798 4924 15862 4928
rect 15798 4868 15802 4924
rect 15802 4868 15858 4924
rect 15858 4868 15862 4924
rect 15798 4864 15862 4868
rect 15878 4924 15942 4928
rect 15878 4868 15882 4924
rect 15882 4868 15938 4924
rect 15938 4868 15942 4924
rect 15878 4864 15942 4868
rect 15958 4924 16022 4928
rect 15958 4868 15962 4924
rect 15962 4868 16018 4924
rect 16018 4868 16022 4924
rect 15958 4864 16022 4868
rect 16038 4924 16102 4928
rect 16038 4868 16042 4924
rect 16042 4868 16098 4924
rect 16098 4868 16102 4924
rect 16038 4864 16102 4868
rect 4521 4380 4585 4384
rect 4521 4324 4525 4380
rect 4525 4324 4581 4380
rect 4581 4324 4585 4380
rect 4521 4320 4585 4324
rect 4601 4380 4665 4384
rect 4601 4324 4605 4380
rect 4605 4324 4661 4380
rect 4661 4324 4665 4380
rect 4601 4320 4665 4324
rect 4681 4380 4745 4384
rect 4681 4324 4685 4380
rect 4685 4324 4741 4380
rect 4741 4324 4745 4380
rect 4681 4320 4745 4324
rect 4761 4380 4825 4384
rect 4761 4324 4765 4380
rect 4765 4324 4821 4380
rect 4821 4324 4825 4380
rect 4761 4320 4825 4324
rect 8500 4380 8564 4384
rect 8500 4324 8504 4380
rect 8504 4324 8560 4380
rect 8560 4324 8564 4380
rect 8500 4320 8564 4324
rect 8580 4380 8644 4384
rect 8580 4324 8584 4380
rect 8584 4324 8640 4380
rect 8640 4324 8644 4380
rect 8580 4320 8644 4324
rect 8660 4380 8724 4384
rect 8660 4324 8664 4380
rect 8664 4324 8720 4380
rect 8720 4324 8724 4380
rect 8660 4320 8724 4324
rect 8740 4380 8804 4384
rect 8740 4324 8744 4380
rect 8744 4324 8800 4380
rect 8800 4324 8804 4380
rect 8740 4320 8804 4324
rect 12479 4380 12543 4384
rect 12479 4324 12483 4380
rect 12483 4324 12539 4380
rect 12539 4324 12543 4380
rect 12479 4320 12543 4324
rect 12559 4380 12623 4384
rect 12559 4324 12563 4380
rect 12563 4324 12619 4380
rect 12619 4324 12623 4380
rect 12559 4320 12623 4324
rect 12639 4380 12703 4384
rect 12639 4324 12643 4380
rect 12643 4324 12699 4380
rect 12699 4324 12703 4380
rect 12639 4320 12703 4324
rect 12719 4380 12783 4384
rect 12719 4324 12723 4380
rect 12723 4324 12779 4380
rect 12779 4324 12783 4380
rect 12719 4320 12783 4324
rect 16458 4380 16522 4384
rect 16458 4324 16462 4380
rect 16462 4324 16518 4380
rect 16518 4324 16522 4380
rect 16458 4320 16522 4324
rect 16538 4380 16602 4384
rect 16538 4324 16542 4380
rect 16542 4324 16598 4380
rect 16598 4324 16602 4380
rect 16538 4320 16602 4324
rect 16618 4380 16682 4384
rect 16618 4324 16622 4380
rect 16622 4324 16678 4380
rect 16678 4324 16682 4380
rect 16618 4320 16682 4324
rect 16698 4380 16762 4384
rect 16698 4324 16702 4380
rect 16702 4324 16758 4380
rect 16758 4324 16762 4380
rect 16698 4320 16762 4324
rect 3861 3836 3925 3840
rect 3861 3780 3865 3836
rect 3865 3780 3921 3836
rect 3921 3780 3925 3836
rect 3861 3776 3925 3780
rect 3941 3836 4005 3840
rect 3941 3780 3945 3836
rect 3945 3780 4001 3836
rect 4001 3780 4005 3836
rect 3941 3776 4005 3780
rect 4021 3836 4085 3840
rect 4021 3780 4025 3836
rect 4025 3780 4081 3836
rect 4081 3780 4085 3836
rect 4021 3776 4085 3780
rect 4101 3836 4165 3840
rect 4101 3780 4105 3836
rect 4105 3780 4161 3836
rect 4161 3780 4165 3836
rect 4101 3776 4165 3780
rect 7840 3836 7904 3840
rect 7840 3780 7844 3836
rect 7844 3780 7900 3836
rect 7900 3780 7904 3836
rect 7840 3776 7904 3780
rect 7920 3836 7984 3840
rect 7920 3780 7924 3836
rect 7924 3780 7980 3836
rect 7980 3780 7984 3836
rect 7920 3776 7984 3780
rect 8000 3836 8064 3840
rect 8000 3780 8004 3836
rect 8004 3780 8060 3836
rect 8060 3780 8064 3836
rect 8000 3776 8064 3780
rect 8080 3836 8144 3840
rect 8080 3780 8084 3836
rect 8084 3780 8140 3836
rect 8140 3780 8144 3836
rect 8080 3776 8144 3780
rect 11819 3836 11883 3840
rect 11819 3780 11823 3836
rect 11823 3780 11879 3836
rect 11879 3780 11883 3836
rect 11819 3776 11883 3780
rect 11899 3836 11963 3840
rect 11899 3780 11903 3836
rect 11903 3780 11959 3836
rect 11959 3780 11963 3836
rect 11899 3776 11963 3780
rect 11979 3836 12043 3840
rect 11979 3780 11983 3836
rect 11983 3780 12039 3836
rect 12039 3780 12043 3836
rect 11979 3776 12043 3780
rect 12059 3836 12123 3840
rect 12059 3780 12063 3836
rect 12063 3780 12119 3836
rect 12119 3780 12123 3836
rect 12059 3776 12123 3780
rect 15798 3836 15862 3840
rect 15798 3780 15802 3836
rect 15802 3780 15858 3836
rect 15858 3780 15862 3836
rect 15798 3776 15862 3780
rect 15878 3836 15942 3840
rect 15878 3780 15882 3836
rect 15882 3780 15938 3836
rect 15938 3780 15942 3836
rect 15878 3776 15942 3780
rect 15958 3836 16022 3840
rect 15958 3780 15962 3836
rect 15962 3780 16018 3836
rect 16018 3780 16022 3836
rect 15958 3776 16022 3780
rect 16038 3836 16102 3840
rect 16038 3780 16042 3836
rect 16042 3780 16098 3836
rect 16098 3780 16102 3836
rect 16038 3776 16102 3780
rect 4521 3292 4585 3296
rect 4521 3236 4525 3292
rect 4525 3236 4581 3292
rect 4581 3236 4585 3292
rect 4521 3232 4585 3236
rect 4601 3292 4665 3296
rect 4601 3236 4605 3292
rect 4605 3236 4661 3292
rect 4661 3236 4665 3292
rect 4601 3232 4665 3236
rect 4681 3292 4745 3296
rect 4681 3236 4685 3292
rect 4685 3236 4741 3292
rect 4741 3236 4745 3292
rect 4681 3232 4745 3236
rect 4761 3292 4825 3296
rect 4761 3236 4765 3292
rect 4765 3236 4821 3292
rect 4821 3236 4825 3292
rect 4761 3232 4825 3236
rect 8500 3292 8564 3296
rect 8500 3236 8504 3292
rect 8504 3236 8560 3292
rect 8560 3236 8564 3292
rect 8500 3232 8564 3236
rect 8580 3292 8644 3296
rect 8580 3236 8584 3292
rect 8584 3236 8640 3292
rect 8640 3236 8644 3292
rect 8580 3232 8644 3236
rect 8660 3292 8724 3296
rect 8660 3236 8664 3292
rect 8664 3236 8720 3292
rect 8720 3236 8724 3292
rect 8660 3232 8724 3236
rect 8740 3292 8804 3296
rect 8740 3236 8744 3292
rect 8744 3236 8800 3292
rect 8800 3236 8804 3292
rect 8740 3232 8804 3236
rect 12479 3292 12543 3296
rect 12479 3236 12483 3292
rect 12483 3236 12539 3292
rect 12539 3236 12543 3292
rect 12479 3232 12543 3236
rect 12559 3292 12623 3296
rect 12559 3236 12563 3292
rect 12563 3236 12619 3292
rect 12619 3236 12623 3292
rect 12559 3232 12623 3236
rect 12639 3292 12703 3296
rect 12639 3236 12643 3292
rect 12643 3236 12699 3292
rect 12699 3236 12703 3292
rect 12639 3232 12703 3236
rect 12719 3292 12783 3296
rect 12719 3236 12723 3292
rect 12723 3236 12779 3292
rect 12779 3236 12783 3292
rect 12719 3232 12783 3236
rect 16458 3292 16522 3296
rect 16458 3236 16462 3292
rect 16462 3236 16518 3292
rect 16518 3236 16522 3292
rect 16458 3232 16522 3236
rect 16538 3292 16602 3296
rect 16538 3236 16542 3292
rect 16542 3236 16598 3292
rect 16598 3236 16602 3292
rect 16538 3232 16602 3236
rect 16618 3292 16682 3296
rect 16618 3236 16622 3292
rect 16622 3236 16678 3292
rect 16678 3236 16682 3292
rect 16618 3232 16682 3236
rect 16698 3292 16762 3296
rect 16698 3236 16702 3292
rect 16702 3236 16758 3292
rect 16758 3236 16762 3292
rect 16698 3232 16762 3236
rect 3861 2748 3925 2752
rect 3861 2692 3865 2748
rect 3865 2692 3921 2748
rect 3921 2692 3925 2748
rect 3861 2688 3925 2692
rect 3941 2748 4005 2752
rect 3941 2692 3945 2748
rect 3945 2692 4001 2748
rect 4001 2692 4005 2748
rect 3941 2688 4005 2692
rect 4021 2748 4085 2752
rect 4021 2692 4025 2748
rect 4025 2692 4081 2748
rect 4081 2692 4085 2748
rect 4021 2688 4085 2692
rect 4101 2748 4165 2752
rect 4101 2692 4105 2748
rect 4105 2692 4161 2748
rect 4161 2692 4165 2748
rect 4101 2688 4165 2692
rect 7840 2748 7904 2752
rect 7840 2692 7844 2748
rect 7844 2692 7900 2748
rect 7900 2692 7904 2748
rect 7840 2688 7904 2692
rect 7920 2748 7984 2752
rect 7920 2692 7924 2748
rect 7924 2692 7980 2748
rect 7980 2692 7984 2748
rect 7920 2688 7984 2692
rect 8000 2748 8064 2752
rect 8000 2692 8004 2748
rect 8004 2692 8060 2748
rect 8060 2692 8064 2748
rect 8000 2688 8064 2692
rect 8080 2748 8144 2752
rect 8080 2692 8084 2748
rect 8084 2692 8140 2748
rect 8140 2692 8144 2748
rect 8080 2688 8144 2692
rect 11819 2748 11883 2752
rect 11819 2692 11823 2748
rect 11823 2692 11879 2748
rect 11879 2692 11883 2748
rect 11819 2688 11883 2692
rect 11899 2748 11963 2752
rect 11899 2692 11903 2748
rect 11903 2692 11959 2748
rect 11959 2692 11963 2748
rect 11899 2688 11963 2692
rect 11979 2748 12043 2752
rect 11979 2692 11983 2748
rect 11983 2692 12039 2748
rect 12039 2692 12043 2748
rect 11979 2688 12043 2692
rect 12059 2748 12123 2752
rect 12059 2692 12063 2748
rect 12063 2692 12119 2748
rect 12119 2692 12123 2748
rect 12059 2688 12123 2692
rect 15798 2748 15862 2752
rect 15798 2692 15802 2748
rect 15802 2692 15858 2748
rect 15858 2692 15862 2748
rect 15798 2688 15862 2692
rect 15878 2748 15942 2752
rect 15878 2692 15882 2748
rect 15882 2692 15938 2748
rect 15938 2692 15942 2748
rect 15878 2688 15942 2692
rect 15958 2748 16022 2752
rect 15958 2692 15962 2748
rect 15962 2692 16018 2748
rect 16018 2692 16022 2748
rect 15958 2688 16022 2692
rect 16038 2748 16102 2752
rect 16038 2692 16042 2748
rect 16042 2692 16098 2748
rect 16098 2692 16102 2748
rect 16038 2688 16102 2692
rect 4521 2204 4585 2208
rect 4521 2148 4525 2204
rect 4525 2148 4581 2204
rect 4581 2148 4585 2204
rect 4521 2144 4585 2148
rect 4601 2204 4665 2208
rect 4601 2148 4605 2204
rect 4605 2148 4661 2204
rect 4661 2148 4665 2204
rect 4601 2144 4665 2148
rect 4681 2204 4745 2208
rect 4681 2148 4685 2204
rect 4685 2148 4741 2204
rect 4741 2148 4745 2204
rect 4681 2144 4745 2148
rect 4761 2204 4825 2208
rect 4761 2148 4765 2204
rect 4765 2148 4821 2204
rect 4821 2148 4825 2204
rect 4761 2144 4825 2148
rect 8500 2204 8564 2208
rect 8500 2148 8504 2204
rect 8504 2148 8560 2204
rect 8560 2148 8564 2204
rect 8500 2144 8564 2148
rect 8580 2204 8644 2208
rect 8580 2148 8584 2204
rect 8584 2148 8640 2204
rect 8640 2148 8644 2204
rect 8580 2144 8644 2148
rect 8660 2204 8724 2208
rect 8660 2148 8664 2204
rect 8664 2148 8720 2204
rect 8720 2148 8724 2204
rect 8660 2144 8724 2148
rect 8740 2204 8804 2208
rect 8740 2148 8744 2204
rect 8744 2148 8800 2204
rect 8800 2148 8804 2204
rect 8740 2144 8804 2148
rect 12479 2204 12543 2208
rect 12479 2148 12483 2204
rect 12483 2148 12539 2204
rect 12539 2148 12543 2204
rect 12479 2144 12543 2148
rect 12559 2204 12623 2208
rect 12559 2148 12563 2204
rect 12563 2148 12619 2204
rect 12619 2148 12623 2204
rect 12559 2144 12623 2148
rect 12639 2204 12703 2208
rect 12639 2148 12643 2204
rect 12643 2148 12699 2204
rect 12699 2148 12703 2204
rect 12639 2144 12703 2148
rect 12719 2204 12783 2208
rect 12719 2148 12723 2204
rect 12723 2148 12779 2204
rect 12779 2148 12783 2204
rect 12719 2144 12783 2148
rect 16458 2204 16522 2208
rect 16458 2148 16462 2204
rect 16462 2148 16518 2204
rect 16518 2148 16522 2204
rect 16458 2144 16522 2148
rect 16538 2204 16602 2208
rect 16538 2148 16542 2204
rect 16542 2148 16598 2204
rect 16598 2148 16602 2204
rect 16538 2144 16602 2148
rect 16618 2204 16682 2208
rect 16618 2148 16622 2204
rect 16622 2148 16678 2204
rect 16678 2148 16682 2204
rect 16618 2144 16682 2148
rect 16698 2204 16762 2208
rect 16698 2148 16702 2204
rect 16702 2148 16758 2204
rect 16758 2148 16762 2204
rect 16698 2144 16762 2148
<< metal4 >>
rect 3853 17984 4173 18000
rect 3853 17920 3861 17984
rect 3925 17920 3941 17984
rect 4005 17920 4021 17984
rect 4085 17920 4101 17984
rect 4165 17920 4173 17984
rect 3853 16896 4173 17920
rect 3853 16832 3861 16896
rect 3925 16832 3941 16896
rect 4005 16832 4021 16896
rect 4085 16832 4101 16896
rect 4165 16832 4173 16896
rect 3853 16098 4173 16832
rect 3853 15862 3895 16098
rect 4131 15862 4173 16098
rect 3853 15808 4173 15862
rect 3853 15744 3861 15808
rect 3925 15744 3941 15808
rect 4005 15744 4021 15808
rect 4085 15744 4101 15808
rect 4165 15744 4173 15808
rect 3853 14720 4173 15744
rect 3853 14656 3861 14720
rect 3925 14656 3941 14720
rect 4005 14656 4021 14720
rect 4085 14656 4101 14720
rect 4165 14656 4173 14720
rect 3853 13632 4173 14656
rect 3853 13568 3861 13632
rect 3925 13568 3941 13632
rect 4005 13568 4021 13632
rect 4085 13568 4101 13632
rect 4165 13568 4173 13632
rect 3853 12544 4173 13568
rect 3853 12480 3861 12544
rect 3925 12480 3941 12544
rect 4005 12480 4021 12544
rect 4085 12480 4101 12544
rect 4165 12480 4173 12544
rect 3853 12154 4173 12480
rect 3853 11918 3895 12154
rect 4131 11918 4173 12154
rect 3853 11456 4173 11918
rect 3853 11392 3861 11456
rect 3925 11392 3941 11456
rect 4005 11392 4021 11456
rect 4085 11392 4101 11456
rect 4165 11392 4173 11456
rect 3853 10368 4173 11392
rect 3853 10304 3861 10368
rect 3925 10304 3941 10368
rect 4005 10304 4021 10368
rect 4085 10304 4101 10368
rect 4165 10304 4173 10368
rect 3853 9280 4173 10304
rect 3853 9216 3861 9280
rect 3925 9216 3941 9280
rect 4005 9216 4021 9280
rect 4085 9216 4101 9280
rect 4165 9216 4173 9280
rect 3853 8210 4173 9216
rect 3853 8192 3895 8210
rect 4131 8192 4173 8210
rect 3853 8128 3861 8192
rect 4165 8128 4173 8192
rect 3853 7974 3895 8128
rect 4131 7974 4173 8128
rect 3853 7104 4173 7974
rect 3853 7040 3861 7104
rect 3925 7040 3941 7104
rect 4005 7040 4021 7104
rect 4085 7040 4101 7104
rect 4165 7040 4173 7104
rect 3853 6016 4173 7040
rect 3853 5952 3861 6016
rect 3925 5952 3941 6016
rect 4005 5952 4021 6016
rect 4085 5952 4101 6016
rect 4165 5952 4173 6016
rect 3853 4928 4173 5952
rect 3853 4864 3861 4928
rect 3925 4864 3941 4928
rect 4005 4864 4021 4928
rect 4085 4864 4101 4928
rect 4165 4864 4173 4928
rect 3853 4266 4173 4864
rect 3853 4030 3895 4266
rect 4131 4030 4173 4266
rect 3853 3840 4173 4030
rect 3853 3776 3861 3840
rect 3925 3776 3941 3840
rect 4005 3776 4021 3840
rect 4085 3776 4101 3840
rect 4165 3776 4173 3840
rect 3853 2752 4173 3776
rect 3853 2688 3861 2752
rect 3925 2688 3941 2752
rect 4005 2688 4021 2752
rect 4085 2688 4101 2752
rect 4165 2688 4173 2752
rect 3853 2128 4173 2688
rect 4513 17440 4833 18000
rect 4513 17376 4521 17440
rect 4585 17376 4601 17440
rect 4665 17376 4681 17440
rect 4745 17376 4761 17440
rect 4825 17376 4833 17440
rect 4513 16758 4833 17376
rect 4513 16522 4555 16758
rect 4791 16522 4833 16758
rect 4513 16352 4833 16522
rect 4513 16288 4521 16352
rect 4585 16288 4601 16352
rect 4665 16288 4681 16352
rect 4745 16288 4761 16352
rect 4825 16288 4833 16352
rect 4513 15264 4833 16288
rect 4513 15200 4521 15264
rect 4585 15200 4601 15264
rect 4665 15200 4681 15264
rect 4745 15200 4761 15264
rect 4825 15200 4833 15264
rect 4513 14176 4833 15200
rect 4513 14112 4521 14176
rect 4585 14112 4601 14176
rect 4665 14112 4681 14176
rect 4745 14112 4761 14176
rect 4825 14112 4833 14176
rect 4513 13088 4833 14112
rect 4513 13024 4521 13088
rect 4585 13024 4601 13088
rect 4665 13024 4681 13088
rect 4745 13024 4761 13088
rect 4825 13024 4833 13088
rect 4513 12814 4833 13024
rect 4513 12578 4555 12814
rect 4791 12578 4833 12814
rect 4513 12000 4833 12578
rect 4513 11936 4521 12000
rect 4585 11936 4601 12000
rect 4665 11936 4681 12000
rect 4745 11936 4761 12000
rect 4825 11936 4833 12000
rect 4513 10912 4833 11936
rect 4513 10848 4521 10912
rect 4585 10848 4601 10912
rect 4665 10848 4681 10912
rect 4745 10848 4761 10912
rect 4825 10848 4833 10912
rect 4513 9824 4833 10848
rect 4513 9760 4521 9824
rect 4585 9760 4601 9824
rect 4665 9760 4681 9824
rect 4745 9760 4761 9824
rect 4825 9760 4833 9824
rect 4513 8870 4833 9760
rect 4513 8736 4555 8870
rect 4791 8736 4833 8870
rect 4513 8672 4521 8736
rect 4825 8672 4833 8736
rect 4513 8634 4555 8672
rect 4791 8634 4833 8672
rect 4513 7648 4833 8634
rect 4513 7584 4521 7648
rect 4585 7584 4601 7648
rect 4665 7584 4681 7648
rect 4745 7584 4761 7648
rect 4825 7584 4833 7648
rect 4513 6560 4833 7584
rect 4513 6496 4521 6560
rect 4585 6496 4601 6560
rect 4665 6496 4681 6560
rect 4745 6496 4761 6560
rect 4825 6496 4833 6560
rect 4513 5472 4833 6496
rect 4513 5408 4521 5472
rect 4585 5408 4601 5472
rect 4665 5408 4681 5472
rect 4745 5408 4761 5472
rect 4825 5408 4833 5472
rect 4513 4926 4833 5408
rect 4513 4690 4555 4926
rect 4791 4690 4833 4926
rect 4513 4384 4833 4690
rect 4513 4320 4521 4384
rect 4585 4320 4601 4384
rect 4665 4320 4681 4384
rect 4745 4320 4761 4384
rect 4825 4320 4833 4384
rect 4513 3296 4833 4320
rect 4513 3232 4521 3296
rect 4585 3232 4601 3296
rect 4665 3232 4681 3296
rect 4745 3232 4761 3296
rect 4825 3232 4833 3296
rect 4513 2208 4833 3232
rect 4513 2144 4521 2208
rect 4585 2144 4601 2208
rect 4665 2144 4681 2208
rect 4745 2144 4761 2208
rect 4825 2144 4833 2208
rect 4513 2128 4833 2144
rect 7832 17984 8152 18000
rect 7832 17920 7840 17984
rect 7904 17920 7920 17984
rect 7984 17920 8000 17984
rect 8064 17920 8080 17984
rect 8144 17920 8152 17984
rect 7832 16896 8152 17920
rect 7832 16832 7840 16896
rect 7904 16832 7920 16896
rect 7984 16832 8000 16896
rect 8064 16832 8080 16896
rect 8144 16832 8152 16896
rect 7832 16098 8152 16832
rect 7832 15862 7874 16098
rect 8110 15862 8152 16098
rect 7832 15808 8152 15862
rect 7832 15744 7840 15808
rect 7904 15744 7920 15808
rect 7984 15744 8000 15808
rect 8064 15744 8080 15808
rect 8144 15744 8152 15808
rect 7832 14720 8152 15744
rect 7832 14656 7840 14720
rect 7904 14656 7920 14720
rect 7984 14656 8000 14720
rect 8064 14656 8080 14720
rect 8144 14656 8152 14720
rect 7832 13632 8152 14656
rect 7832 13568 7840 13632
rect 7904 13568 7920 13632
rect 7984 13568 8000 13632
rect 8064 13568 8080 13632
rect 8144 13568 8152 13632
rect 7832 12544 8152 13568
rect 7832 12480 7840 12544
rect 7904 12480 7920 12544
rect 7984 12480 8000 12544
rect 8064 12480 8080 12544
rect 8144 12480 8152 12544
rect 7832 12154 8152 12480
rect 7832 11918 7874 12154
rect 8110 11918 8152 12154
rect 7832 11456 8152 11918
rect 7832 11392 7840 11456
rect 7904 11392 7920 11456
rect 7984 11392 8000 11456
rect 8064 11392 8080 11456
rect 8144 11392 8152 11456
rect 7832 10368 8152 11392
rect 7832 10304 7840 10368
rect 7904 10304 7920 10368
rect 7984 10304 8000 10368
rect 8064 10304 8080 10368
rect 8144 10304 8152 10368
rect 7832 9280 8152 10304
rect 7832 9216 7840 9280
rect 7904 9216 7920 9280
rect 7984 9216 8000 9280
rect 8064 9216 8080 9280
rect 8144 9216 8152 9280
rect 7832 8210 8152 9216
rect 7832 8192 7874 8210
rect 8110 8192 8152 8210
rect 7832 8128 7840 8192
rect 8144 8128 8152 8192
rect 7832 7974 7874 8128
rect 8110 7974 8152 8128
rect 7832 7104 8152 7974
rect 7832 7040 7840 7104
rect 7904 7040 7920 7104
rect 7984 7040 8000 7104
rect 8064 7040 8080 7104
rect 8144 7040 8152 7104
rect 7832 6016 8152 7040
rect 7832 5952 7840 6016
rect 7904 5952 7920 6016
rect 7984 5952 8000 6016
rect 8064 5952 8080 6016
rect 8144 5952 8152 6016
rect 7832 4928 8152 5952
rect 7832 4864 7840 4928
rect 7904 4864 7920 4928
rect 7984 4864 8000 4928
rect 8064 4864 8080 4928
rect 8144 4864 8152 4928
rect 7832 4266 8152 4864
rect 7832 4030 7874 4266
rect 8110 4030 8152 4266
rect 7832 3840 8152 4030
rect 7832 3776 7840 3840
rect 7904 3776 7920 3840
rect 7984 3776 8000 3840
rect 8064 3776 8080 3840
rect 8144 3776 8152 3840
rect 7832 2752 8152 3776
rect 7832 2688 7840 2752
rect 7904 2688 7920 2752
rect 7984 2688 8000 2752
rect 8064 2688 8080 2752
rect 8144 2688 8152 2752
rect 7832 2128 8152 2688
rect 8492 17440 8812 18000
rect 8492 17376 8500 17440
rect 8564 17376 8580 17440
rect 8644 17376 8660 17440
rect 8724 17376 8740 17440
rect 8804 17376 8812 17440
rect 8492 16758 8812 17376
rect 8492 16522 8534 16758
rect 8770 16522 8812 16758
rect 8492 16352 8812 16522
rect 8492 16288 8500 16352
rect 8564 16288 8580 16352
rect 8644 16288 8660 16352
rect 8724 16288 8740 16352
rect 8804 16288 8812 16352
rect 8492 15264 8812 16288
rect 8492 15200 8500 15264
rect 8564 15200 8580 15264
rect 8644 15200 8660 15264
rect 8724 15200 8740 15264
rect 8804 15200 8812 15264
rect 8492 14176 8812 15200
rect 8492 14112 8500 14176
rect 8564 14112 8580 14176
rect 8644 14112 8660 14176
rect 8724 14112 8740 14176
rect 8804 14112 8812 14176
rect 8492 13088 8812 14112
rect 8492 13024 8500 13088
rect 8564 13024 8580 13088
rect 8644 13024 8660 13088
rect 8724 13024 8740 13088
rect 8804 13024 8812 13088
rect 8492 12814 8812 13024
rect 8492 12578 8534 12814
rect 8770 12578 8812 12814
rect 8492 12000 8812 12578
rect 8492 11936 8500 12000
rect 8564 11936 8580 12000
rect 8644 11936 8660 12000
rect 8724 11936 8740 12000
rect 8804 11936 8812 12000
rect 8492 10912 8812 11936
rect 8492 10848 8500 10912
rect 8564 10848 8580 10912
rect 8644 10848 8660 10912
rect 8724 10848 8740 10912
rect 8804 10848 8812 10912
rect 8492 9824 8812 10848
rect 8492 9760 8500 9824
rect 8564 9760 8580 9824
rect 8644 9760 8660 9824
rect 8724 9760 8740 9824
rect 8804 9760 8812 9824
rect 8492 8870 8812 9760
rect 8492 8736 8534 8870
rect 8770 8736 8812 8870
rect 8492 8672 8500 8736
rect 8804 8672 8812 8736
rect 8492 8634 8534 8672
rect 8770 8634 8812 8672
rect 8492 7648 8812 8634
rect 8492 7584 8500 7648
rect 8564 7584 8580 7648
rect 8644 7584 8660 7648
rect 8724 7584 8740 7648
rect 8804 7584 8812 7648
rect 8492 6560 8812 7584
rect 8492 6496 8500 6560
rect 8564 6496 8580 6560
rect 8644 6496 8660 6560
rect 8724 6496 8740 6560
rect 8804 6496 8812 6560
rect 8492 5472 8812 6496
rect 8492 5408 8500 5472
rect 8564 5408 8580 5472
rect 8644 5408 8660 5472
rect 8724 5408 8740 5472
rect 8804 5408 8812 5472
rect 8492 4926 8812 5408
rect 8492 4690 8534 4926
rect 8770 4690 8812 4926
rect 8492 4384 8812 4690
rect 8492 4320 8500 4384
rect 8564 4320 8580 4384
rect 8644 4320 8660 4384
rect 8724 4320 8740 4384
rect 8804 4320 8812 4384
rect 8492 3296 8812 4320
rect 8492 3232 8500 3296
rect 8564 3232 8580 3296
rect 8644 3232 8660 3296
rect 8724 3232 8740 3296
rect 8804 3232 8812 3296
rect 8492 2208 8812 3232
rect 8492 2144 8500 2208
rect 8564 2144 8580 2208
rect 8644 2144 8660 2208
rect 8724 2144 8740 2208
rect 8804 2144 8812 2208
rect 8492 2128 8812 2144
rect 11811 17984 12131 18000
rect 11811 17920 11819 17984
rect 11883 17920 11899 17984
rect 11963 17920 11979 17984
rect 12043 17920 12059 17984
rect 12123 17920 12131 17984
rect 11811 16896 12131 17920
rect 11811 16832 11819 16896
rect 11883 16832 11899 16896
rect 11963 16832 11979 16896
rect 12043 16832 12059 16896
rect 12123 16832 12131 16896
rect 11811 16098 12131 16832
rect 11811 15862 11853 16098
rect 12089 15862 12131 16098
rect 11811 15808 12131 15862
rect 11811 15744 11819 15808
rect 11883 15744 11899 15808
rect 11963 15744 11979 15808
rect 12043 15744 12059 15808
rect 12123 15744 12131 15808
rect 11811 14720 12131 15744
rect 11811 14656 11819 14720
rect 11883 14656 11899 14720
rect 11963 14656 11979 14720
rect 12043 14656 12059 14720
rect 12123 14656 12131 14720
rect 11811 13632 12131 14656
rect 11811 13568 11819 13632
rect 11883 13568 11899 13632
rect 11963 13568 11979 13632
rect 12043 13568 12059 13632
rect 12123 13568 12131 13632
rect 11811 12544 12131 13568
rect 11811 12480 11819 12544
rect 11883 12480 11899 12544
rect 11963 12480 11979 12544
rect 12043 12480 12059 12544
rect 12123 12480 12131 12544
rect 11811 12154 12131 12480
rect 11811 11918 11853 12154
rect 12089 11918 12131 12154
rect 11811 11456 12131 11918
rect 11811 11392 11819 11456
rect 11883 11392 11899 11456
rect 11963 11392 11979 11456
rect 12043 11392 12059 11456
rect 12123 11392 12131 11456
rect 11811 10368 12131 11392
rect 11811 10304 11819 10368
rect 11883 10304 11899 10368
rect 11963 10304 11979 10368
rect 12043 10304 12059 10368
rect 12123 10304 12131 10368
rect 11811 9280 12131 10304
rect 11811 9216 11819 9280
rect 11883 9216 11899 9280
rect 11963 9216 11979 9280
rect 12043 9216 12059 9280
rect 12123 9216 12131 9280
rect 11811 8210 12131 9216
rect 11811 8192 11853 8210
rect 12089 8192 12131 8210
rect 11811 8128 11819 8192
rect 12123 8128 12131 8192
rect 11811 7974 11853 8128
rect 12089 7974 12131 8128
rect 11811 7104 12131 7974
rect 11811 7040 11819 7104
rect 11883 7040 11899 7104
rect 11963 7040 11979 7104
rect 12043 7040 12059 7104
rect 12123 7040 12131 7104
rect 11811 6016 12131 7040
rect 11811 5952 11819 6016
rect 11883 5952 11899 6016
rect 11963 5952 11979 6016
rect 12043 5952 12059 6016
rect 12123 5952 12131 6016
rect 11811 4928 12131 5952
rect 11811 4864 11819 4928
rect 11883 4864 11899 4928
rect 11963 4864 11979 4928
rect 12043 4864 12059 4928
rect 12123 4864 12131 4928
rect 11811 4266 12131 4864
rect 11811 4030 11853 4266
rect 12089 4030 12131 4266
rect 11811 3840 12131 4030
rect 11811 3776 11819 3840
rect 11883 3776 11899 3840
rect 11963 3776 11979 3840
rect 12043 3776 12059 3840
rect 12123 3776 12131 3840
rect 11811 2752 12131 3776
rect 11811 2688 11819 2752
rect 11883 2688 11899 2752
rect 11963 2688 11979 2752
rect 12043 2688 12059 2752
rect 12123 2688 12131 2752
rect 11811 2128 12131 2688
rect 12471 17440 12791 18000
rect 12471 17376 12479 17440
rect 12543 17376 12559 17440
rect 12623 17376 12639 17440
rect 12703 17376 12719 17440
rect 12783 17376 12791 17440
rect 12471 16758 12791 17376
rect 12471 16522 12513 16758
rect 12749 16522 12791 16758
rect 12471 16352 12791 16522
rect 12471 16288 12479 16352
rect 12543 16288 12559 16352
rect 12623 16288 12639 16352
rect 12703 16288 12719 16352
rect 12783 16288 12791 16352
rect 12471 15264 12791 16288
rect 12471 15200 12479 15264
rect 12543 15200 12559 15264
rect 12623 15200 12639 15264
rect 12703 15200 12719 15264
rect 12783 15200 12791 15264
rect 12471 14176 12791 15200
rect 12471 14112 12479 14176
rect 12543 14112 12559 14176
rect 12623 14112 12639 14176
rect 12703 14112 12719 14176
rect 12783 14112 12791 14176
rect 12471 13088 12791 14112
rect 12471 13024 12479 13088
rect 12543 13024 12559 13088
rect 12623 13024 12639 13088
rect 12703 13024 12719 13088
rect 12783 13024 12791 13088
rect 12471 12814 12791 13024
rect 12471 12578 12513 12814
rect 12749 12578 12791 12814
rect 12471 12000 12791 12578
rect 12471 11936 12479 12000
rect 12543 11936 12559 12000
rect 12623 11936 12639 12000
rect 12703 11936 12719 12000
rect 12783 11936 12791 12000
rect 12471 10912 12791 11936
rect 12471 10848 12479 10912
rect 12543 10848 12559 10912
rect 12623 10848 12639 10912
rect 12703 10848 12719 10912
rect 12783 10848 12791 10912
rect 12471 9824 12791 10848
rect 12471 9760 12479 9824
rect 12543 9760 12559 9824
rect 12623 9760 12639 9824
rect 12703 9760 12719 9824
rect 12783 9760 12791 9824
rect 12471 8870 12791 9760
rect 12471 8736 12513 8870
rect 12749 8736 12791 8870
rect 12471 8672 12479 8736
rect 12783 8672 12791 8736
rect 12471 8634 12513 8672
rect 12749 8634 12791 8672
rect 12471 7648 12791 8634
rect 12471 7584 12479 7648
rect 12543 7584 12559 7648
rect 12623 7584 12639 7648
rect 12703 7584 12719 7648
rect 12783 7584 12791 7648
rect 12471 6560 12791 7584
rect 12471 6496 12479 6560
rect 12543 6496 12559 6560
rect 12623 6496 12639 6560
rect 12703 6496 12719 6560
rect 12783 6496 12791 6560
rect 12471 5472 12791 6496
rect 12471 5408 12479 5472
rect 12543 5408 12559 5472
rect 12623 5408 12639 5472
rect 12703 5408 12719 5472
rect 12783 5408 12791 5472
rect 12471 4926 12791 5408
rect 12471 4690 12513 4926
rect 12749 4690 12791 4926
rect 12471 4384 12791 4690
rect 12471 4320 12479 4384
rect 12543 4320 12559 4384
rect 12623 4320 12639 4384
rect 12703 4320 12719 4384
rect 12783 4320 12791 4384
rect 12471 3296 12791 4320
rect 12471 3232 12479 3296
rect 12543 3232 12559 3296
rect 12623 3232 12639 3296
rect 12703 3232 12719 3296
rect 12783 3232 12791 3296
rect 12471 2208 12791 3232
rect 12471 2144 12479 2208
rect 12543 2144 12559 2208
rect 12623 2144 12639 2208
rect 12703 2144 12719 2208
rect 12783 2144 12791 2208
rect 12471 2128 12791 2144
rect 15790 17984 16110 18000
rect 15790 17920 15798 17984
rect 15862 17920 15878 17984
rect 15942 17920 15958 17984
rect 16022 17920 16038 17984
rect 16102 17920 16110 17984
rect 15790 16896 16110 17920
rect 15790 16832 15798 16896
rect 15862 16832 15878 16896
rect 15942 16832 15958 16896
rect 16022 16832 16038 16896
rect 16102 16832 16110 16896
rect 15790 16098 16110 16832
rect 15790 15862 15832 16098
rect 16068 15862 16110 16098
rect 15790 15808 16110 15862
rect 15790 15744 15798 15808
rect 15862 15744 15878 15808
rect 15942 15744 15958 15808
rect 16022 15744 16038 15808
rect 16102 15744 16110 15808
rect 15790 14720 16110 15744
rect 15790 14656 15798 14720
rect 15862 14656 15878 14720
rect 15942 14656 15958 14720
rect 16022 14656 16038 14720
rect 16102 14656 16110 14720
rect 15790 13632 16110 14656
rect 15790 13568 15798 13632
rect 15862 13568 15878 13632
rect 15942 13568 15958 13632
rect 16022 13568 16038 13632
rect 16102 13568 16110 13632
rect 15790 12544 16110 13568
rect 15790 12480 15798 12544
rect 15862 12480 15878 12544
rect 15942 12480 15958 12544
rect 16022 12480 16038 12544
rect 16102 12480 16110 12544
rect 15790 12154 16110 12480
rect 15790 11918 15832 12154
rect 16068 11918 16110 12154
rect 15790 11456 16110 11918
rect 15790 11392 15798 11456
rect 15862 11392 15878 11456
rect 15942 11392 15958 11456
rect 16022 11392 16038 11456
rect 16102 11392 16110 11456
rect 15790 10368 16110 11392
rect 15790 10304 15798 10368
rect 15862 10304 15878 10368
rect 15942 10304 15958 10368
rect 16022 10304 16038 10368
rect 16102 10304 16110 10368
rect 15790 9280 16110 10304
rect 15790 9216 15798 9280
rect 15862 9216 15878 9280
rect 15942 9216 15958 9280
rect 16022 9216 16038 9280
rect 16102 9216 16110 9280
rect 15790 8210 16110 9216
rect 15790 8192 15832 8210
rect 16068 8192 16110 8210
rect 15790 8128 15798 8192
rect 16102 8128 16110 8192
rect 15790 7974 15832 8128
rect 16068 7974 16110 8128
rect 15790 7104 16110 7974
rect 15790 7040 15798 7104
rect 15862 7040 15878 7104
rect 15942 7040 15958 7104
rect 16022 7040 16038 7104
rect 16102 7040 16110 7104
rect 15790 6016 16110 7040
rect 15790 5952 15798 6016
rect 15862 5952 15878 6016
rect 15942 5952 15958 6016
rect 16022 5952 16038 6016
rect 16102 5952 16110 6016
rect 15790 4928 16110 5952
rect 15790 4864 15798 4928
rect 15862 4864 15878 4928
rect 15942 4864 15958 4928
rect 16022 4864 16038 4928
rect 16102 4864 16110 4928
rect 15790 4266 16110 4864
rect 15790 4030 15832 4266
rect 16068 4030 16110 4266
rect 15790 3840 16110 4030
rect 15790 3776 15798 3840
rect 15862 3776 15878 3840
rect 15942 3776 15958 3840
rect 16022 3776 16038 3840
rect 16102 3776 16110 3840
rect 15790 2752 16110 3776
rect 15790 2688 15798 2752
rect 15862 2688 15878 2752
rect 15942 2688 15958 2752
rect 16022 2688 16038 2752
rect 16102 2688 16110 2752
rect 15790 2128 16110 2688
rect 16450 17440 16770 18000
rect 16450 17376 16458 17440
rect 16522 17376 16538 17440
rect 16602 17376 16618 17440
rect 16682 17376 16698 17440
rect 16762 17376 16770 17440
rect 16450 16758 16770 17376
rect 16450 16522 16492 16758
rect 16728 16522 16770 16758
rect 16450 16352 16770 16522
rect 16450 16288 16458 16352
rect 16522 16288 16538 16352
rect 16602 16288 16618 16352
rect 16682 16288 16698 16352
rect 16762 16288 16770 16352
rect 16450 15264 16770 16288
rect 16450 15200 16458 15264
rect 16522 15200 16538 15264
rect 16602 15200 16618 15264
rect 16682 15200 16698 15264
rect 16762 15200 16770 15264
rect 16450 14176 16770 15200
rect 16450 14112 16458 14176
rect 16522 14112 16538 14176
rect 16602 14112 16618 14176
rect 16682 14112 16698 14176
rect 16762 14112 16770 14176
rect 16450 13088 16770 14112
rect 16450 13024 16458 13088
rect 16522 13024 16538 13088
rect 16602 13024 16618 13088
rect 16682 13024 16698 13088
rect 16762 13024 16770 13088
rect 16450 12814 16770 13024
rect 16450 12578 16492 12814
rect 16728 12578 16770 12814
rect 16450 12000 16770 12578
rect 16450 11936 16458 12000
rect 16522 11936 16538 12000
rect 16602 11936 16618 12000
rect 16682 11936 16698 12000
rect 16762 11936 16770 12000
rect 16450 10912 16770 11936
rect 16450 10848 16458 10912
rect 16522 10848 16538 10912
rect 16602 10848 16618 10912
rect 16682 10848 16698 10912
rect 16762 10848 16770 10912
rect 16450 9824 16770 10848
rect 16450 9760 16458 9824
rect 16522 9760 16538 9824
rect 16602 9760 16618 9824
rect 16682 9760 16698 9824
rect 16762 9760 16770 9824
rect 16450 8870 16770 9760
rect 16450 8736 16492 8870
rect 16728 8736 16770 8870
rect 16450 8672 16458 8736
rect 16762 8672 16770 8736
rect 16450 8634 16492 8672
rect 16728 8634 16770 8672
rect 16450 7648 16770 8634
rect 16450 7584 16458 7648
rect 16522 7584 16538 7648
rect 16602 7584 16618 7648
rect 16682 7584 16698 7648
rect 16762 7584 16770 7648
rect 16450 6560 16770 7584
rect 16450 6496 16458 6560
rect 16522 6496 16538 6560
rect 16602 6496 16618 6560
rect 16682 6496 16698 6560
rect 16762 6496 16770 6560
rect 16450 5472 16770 6496
rect 16450 5408 16458 5472
rect 16522 5408 16538 5472
rect 16602 5408 16618 5472
rect 16682 5408 16698 5472
rect 16762 5408 16770 5472
rect 16450 4926 16770 5408
rect 16450 4690 16492 4926
rect 16728 4690 16770 4926
rect 16450 4384 16770 4690
rect 16450 4320 16458 4384
rect 16522 4320 16538 4384
rect 16602 4320 16618 4384
rect 16682 4320 16698 4384
rect 16762 4320 16770 4384
rect 16450 3296 16770 4320
rect 16450 3232 16458 3296
rect 16522 3232 16538 3296
rect 16602 3232 16618 3296
rect 16682 3232 16698 3296
rect 16762 3232 16770 3296
rect 16450 2208 16770 3232
rect 16450 2144 16458 2208
rect 16522 2144 16538 2208
rect 16602 2144 16618 2208
rect 16682 2144 16698 2208
rect 16762 2144 16770 2208
rect 16450 2128 16770 2144
<< via4 >>
rect 3895 15862 4131 16098
rect 3895 11918 4131 12154
rect 3895 8192 4131 8210
rect 3895 8128 3925 8192
rect 3925 8128 3941 8192
rect 3941 8128 4005 8192
rect 4005 8128 4021 8192
rect 4021 8128 4085 8192
rect 4085 8128 4101 8192
rect 4101 8128 4131 8192
rect 3895 7974 4131 8128
rect 3895 4030 4131 4266
rect 4555 16522 4791 16758
rect 4555 12578 4791 12814
rect 4555 8736 4791 8870
rect 4555 8672 4585 8736
rect 4585 8672 4601 8736
rect 4601 8672 4665 8736
rect 4665 8672 4681 8736
rect 4681 8672 4745 8736
rect 4745 8672 4761 8736
rect 4761 8672 4791 8736
rect 4555 8634 4791 8672
rect 4555 4690 4791 4926
rect 7874 15862 8110 16098
rect 7874 11918 8110 12154
rect 7874 8192 8110 8210
rect 7874 8128 7904 8192
rect 7904 8128 7920 8192
rect 7920 8128 7984 8192
rect 7984 8128 8000 8192
rect 8000 8128 8064 8192
rect 8064 8128 8080 8192
rect 8080 8128 8110 8192
rect 7874 7974 8110 8128
rect 7874 4030 8110 4266
rect 8534 16522 8770 16758
rect 8534 12578 8770 12814
rect 8534 8736 8770 8870
rect 8534 8672 8564 8736
rect 8564 8672 8580 8736
rect 8580 8672 8644 8736
rect 8644 8672 8660 8736
rect 8660 8672 8724 8736
rect 8724 8672 8740 8736
rect 8740 8672 8770 8736
rect 8534 8634 8770 8672
rect 8534 4690 8770 4926
rect 11853 15862 12089 16098
rect 11853 11918 12089 12154
rect 11853 8192 12089 8210
rect 11853 8128 11883 8192
rect 11883 8128 11899 8192
rect 11899 8128 11963 8192
rect 11963 8128 11979 8192
rect 11979 8128 12043 8192
rect 12043 8128 12059 8192
rect 12059 8128 12089 8192
rect 11853 7974 12089 8128
rect 11853 4030 12089 4266
rect 12513 16522 12749 16758
rect 12513 12578 12749 12814
rect 12513 8736 12749 8870
rect 12513 8672 12543 8736
rect 12543 8672 12559 8736
rect 12559 8672 12623 8736
rect 12623 8672 12639 8736
rect 12639 8672 12703 8736
rect 12703 8672 12719 8736
rect 12719 8672 12749 8736
rect 12513 8634 12749 8672
rect 12513 4690 12749 4926
rect 15832 15862 16068 16098
rect 15832 11918 16068 12154
rect 15832 8192 16068 8210
rect 15832 8128 15862 8192
rect 15862 8128 15878 8192
rect 15878 8128 15942 8192
rect 15942 8128 15958 8192
rect 15958 8128 16022 8192
rect 16022 8128 16038 8192
rect 16038 8128 16068 8192
rect 15832 7974 16068 8128
rect 15832 4030 16068 4266
rect 16492 16522 16728 16758
rect 16492 12578 16728 12814
rect 16492 8736 16728 8870
rect 16492 8672 16522 8736
rect 16522 8672 16538 8736
rect 16538 8672 16602 8736
rect 16602 8672 16618 8736
rect 16618 8672 16682 8736
rect 16682 8672 16698 8736
rect 16698 8672 16728 8736
rect 16492 8634 16728 8672
rect 16492 4690 16728 4926
<< metal5 >>
rect 1976 16758 17988 16800
rect 1976 16522 4555 16758
rect 4791 16522 8534 16758
rect 8770 16522 12513 16758
rect 12749 16522 16492 16758
rect 16728 16522 17988 16758
rect 1976 16480 17988 16522
rect 1976 16098 17988 16140
rect 1976 15862 3895 16098
rect 4131 15862 7874 16098
rect 8110 15862 11853 16098
rect 12089 15862 15832 16098
rect 16068 15862 17988 16098
rect 1976 15820 17988 15862
rect 1976 12814 17988 12856
rect 1976 12578 4555 12814
rect 4791 12578 8534 12814
rect 8770 12578 12513 12814
rect 12749 12578 16492 12814
rect 16728 12578 17988 12814
rect 1976 12536 17988 12578
rect 1976 12154 17988 12196
rect 1976 11918 3895 12154
rect 4131 11918 7874 12154
rect 8110 11918 11853 12154
rect 12089 11918 15832 12154
rect 16068 11918 17988 12154
rect 1976 11876 17988 11918
rect 1976 8870 17988 8912
rect 1976 8634 4555 8870
rect 4791 8634 8534 8870
rect 8770 8634 12513 8870
rect 12749 8634 16492 8870
rect 16728 8634 17988 8870
rect 1976 8592 17988 8634
rect 1976 8210 17988 8252
rect 1976 7974 3895 8210
rect 4131 7974 7874 8210
rect 8110 7974 11853 8210
rect 12089 7974 15832 8210
rect 16068 7974 17988 8210
rect 1976 7932 17988 7974
rect 1976 4926 17988 4968
rect 1976 4690 4555 4926
rect 4791 4690 8534 4926
rect 8770 4690 12513 4926
rect 12749 4690 16492 4926
rect 16728 4690 17988 4926
rect 1976 4648 17988 4690
rect 1976 4266 17988 4308
rect 1976 4030 3895 4266
rect 4131 4030 7874 4266
rect 8110 4030 11853 4266
rect 12089 4030 15832 4266
rect 16068 4030 17988 4266
rect 1976 3988 17988 4030
use sky130_fd_sc_hd__inv_2  _113_
timestamp 0
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 0
transform 1 0 8648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _115_
timestamp 0
transform -1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 0
transform -1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _117_
timestamp 0
transform -1 0 10304 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _118_
timestamp 0
transform -1 0 8924 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 0
transform 1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _120_
timestamp 0
transform 1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _121_
timestamp 0
transform -1 0 8464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _122_
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _123_
timestamp 0
transform -1 0 9660 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _124_
timestamp 0
transform -1 0 8188 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 0
transform -1 0 7820 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _126_
timestamp 0
transform 1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _127_
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 0
transform 1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _129_
timestamp 0
transform -1 0 8188 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 0
transform 1 0 6808 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _131_
timestamp 0
transform 1 0 8280 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 0
transform 1 0 9108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _133_
timestamp 0
transform 1 0 12052 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _134_
timestamp 0
transform -1 0 11868 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _135_
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _136_
timestamp 0
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _137_
timestamp 0
transform 1 0 10488 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _138_
timestamp 0
transform 1 0 9844 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _139_
timestamp 0
transform 1 0 8648 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _140_
timestamp 0
transform 1 0 7268 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 0
transform -1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _142_
timestamp 0
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _143_
timestamp 0
transform -1 0 11316 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _144_
timestamp 0
transform -1 0 10304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _145_
timestamp 0
transform 1 0 7360 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _146_
timestamp 0
transform 1 0 7176 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _147_
timestamp 0
transform 1 0 10120 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _148_
timestamp 0
transform -1 0 10948 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _149_
timestamp 0
transform 1 0 10948 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _150_
timestamp 0
transform -1 0 10672 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _151_
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _152_
timestamp 0
transform -1 0 13892 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _153_
timestamp 0
transform -1 0 13248 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _154_
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _155_
timestamp 0
transform 1 0 12420 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _156_
timestamp 0
transform 1 0 11960 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _157_
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _158_
timestamp 0
transform 1 0 13064 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _159_
timestamp 0
transform -1 0 14168 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _160_
timestamp 0
transform 1 0 14168 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _162_
timestamp 0
transform -1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _163_
timestamp 0
transform 1 0 14352 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _164_
timestamp 0
transform 1 0 14996 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _165_
timestamp 0
transform -1 0 15088 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _166_
timestamp 0
transform -1 0 13892 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _167_
timestamp 0
transform 1 0 12972 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _168_
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _169_
timestamp 0
transform -1 0 14904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _170_
timestamp 0
transform -1 0 15088 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _171_
timestamp 0
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 0
transform -1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _173_
timestamp 0
transform -1 0 15548 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _174_
timestamp 0
transform -1 0 15456 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _175_
timestamp 0
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _176_
timestamp 0
transform 1 0 12880 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _177_
timestamp 0
transform 1 0 12144 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _178_
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _179_
timestamp 0
transform -1 0 12052 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _180_
timestamp 0
transform -1 0 13248 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _181_
timestamp 0
transform 1 0 13524 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _182_
timestamp 0
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _183_
timestamp 0
transform 1 0 13064 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _184_
timestamp 0
transform 1 0 13432 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _185_
timestamp 0
transform -1 0 13432 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _186_
timestamp 0
transform -1 0 13524 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _187_
timestamp 0
transform -1 0 15732 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _188_
timestamp 0
transform 1 0 14168 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _189_
timestamp 0
transform -1 0 13064 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _190_
timestamp 0
transform 1 0 12512 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _191_
timestamp 0
transform 1 0 13156 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _192_
timestamp 0
transform -1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _193_
timestamp 0
transform 1 0 11224 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _194_
timestamp 0
transform 1 0 12420 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _195_
timestamp 0
transform -1 0 12604 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _196_
timestamp 0
transform 1 0 13800 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _197_
timestamp 0
transform -1 0 10672 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _198_
timestamp 0
transform 1 0 10028 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _199_
timestamp 0
transform 1 0 10396 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _200_
timestamp 0
transform 1 0 11040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _201_
timestamp 0
transform -1 0 11868 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _202_
timestamp 0
transform 1 0 10396 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _203_
timestamp 0
transform -1 0 11040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _204_
timestamp 0
transform -1 0 11224 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _205_
timestamp 0
transform -1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _206_
timestamp 0
transform 1 0 10212 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _207_
timestamp 0
transform 1 0 10304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _208_
timestamp 0
transform -1 0 11868 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _209_
timestamp 0
transform 1 0 9752 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _210_
timestamp 0
transform 1 0 8280 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _211_
timestamp 0
transform -1 0 9476 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _212_
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _213_
timestamp 0
transform -1 0 9016 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _214_
timestamp 0
transform -1 0 10028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _215_
timestamp 0
transform -1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _216_
timestamp 0
transform 1 0 10672 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _217_
timestamp 0
transform 1 0 8372 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _218_
timestamp 0
transform 1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _219_
timestamp 0
transform 1 0 8740 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _220_
timestamp 0
transform -1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _221_
timestamp 0
transform -1 0 8740 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _222_
timestamp 0
transform 1 0 8556 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _223_
timestamp 0
transform 1 0 8648 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _224_
timestamp 0
transform 1 0 9016 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _225_
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _226_
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _227_
timestamp 0
transform 1 0 6348 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _228_
timestamp 0
transform 1 0 6532 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _229_
timestamp 0
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _230_
timestamp 0
transform 1 0 7268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _231_
timestamp 0
transform -1 0 7176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _232_
timestamp 0
transform -1 0 7728 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _233_
timestamp 0
transform 1 0 7176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 0
transform -1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 3404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 4692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 5796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_57
timestamp 0
transform 1 0 7268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_76
timestamp 0
transform 1 0 9016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_95
timestamp 0
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_102
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_123
timestamp 0
transform 1 0 13340 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 0
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 0
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14996 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 16100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 0
transform 1 0 17572 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 2300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 3404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 4508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 5612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 7268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 8372 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_81
timestamp 0
transform 1 0 9476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_89
timestamp 0
transform 1 0 10212 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_95
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_107
timestamp 0
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 12420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 15732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 0
transform 1 0 17572 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 3404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 8004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 9108 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 9844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 12052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 13156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 14260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 16100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_165
timestamp 0
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_169
timestamp 0
transform 1 0 17572 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 2300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 3404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 5612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 7268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 10580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 11684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 12420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 13524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 15732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 0
transform 1 0 16836 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp 0
transform 1 0 17572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 3404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 4692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 5796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 8004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 9108 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 9660 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 9844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 13156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 0
transform 1 0 14260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 14812 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 0
transform 1 0 16100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_165
timestamp 0
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_169
timestamp 0
transform 1 0 17572 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 5612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 7268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 8372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 10580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 11684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 12420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 14628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 15732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 16836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 0
transform 1 0 17572 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 2300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 3404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 8004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 9108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 9844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_97
timestamp 0
transform 1 0 10948 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_105
timestamp 0
transform 1 0 11684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_117
timestamp 0
transform 1 0 12788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 0
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 0
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_165
timestamp 0
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_169
timestamp 0
transform 1 0 17572 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 5612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 0
transform 1 0 7268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_74
timestamp 0
transform 1 0 8832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_82
timestamp 0
transform 1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 12420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 13524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 14628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 15732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 16836 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 17388 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 0
transform 1 0 17572 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 3404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 4692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_53
timestamp 0
transform 1 0 6900 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_90
timestamp 0
transform 1 0 10304 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_107
timestamp 0
transform 1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_113
timestamp 0
transform 1 0 12420 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_119
timestamp 0
transform 1 0 12972 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_125
timestamp 0
transform 1 0 13524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_136
timestamp 0
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_165
timestamp 0
transform 1 0 17204 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_169
timestamp 0
transform 1 0 17572 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 5612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_51
timestamp 0
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_67
timestamp 0
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_78
timestamp 0
transform 1 0 9200 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_90
timestamp 0
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_102
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 0
transform 1 0 12144 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_113
timestamp 0
transform 1 0 12420 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_124
timestamp 0
transform 1 0 13432 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_132
timestamp 0
transform 1 0 14168 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_143
timestamp 0
transform 1 0 15180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_155
timestamp 0
transform 1 0 16284 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 17388 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 0
transform 1 0 17572 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 3404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 5796 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_53
timestamp 0
transform 1 0 6900 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_63
timestamp 0
transform 1 0 7820 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_75
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_85
timestamp 0
transform 1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_105
timestamp 0
transform 1 0 11684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_132
timestamp 0
transform 1 0 14168 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_144
timestamp 0
transform 1 0 15272 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_156
timestamp 0
transform 1 0 16376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 5612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_51
timestamp 0
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 0
transform 1 0 7268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_70
timestamp 0
transform 1 0 8464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_83
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_106
timestamp 0
transform 1 0 11776 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_129
timestamp 0
transform 1 0 13892 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_142
timestamp 0
transform 1 0 15088 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_154
timestamp 0
transform 1 0 16192 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_162
timestamp 0
transform 1 0 16928 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_169
timestamp 0
transform 1 0 17572 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_7
timestamp 0
transform 1 0 2668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_19
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_41
timestamp 0
transform 1 0 5796 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_49
timestamp 0
transform 1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_67
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 0
transform 1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 0
transform 1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_95
timestamp 0
transform 1 0 10764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_107
timestamp 0
transform 1 0 11868 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_119
timestamp 0
transform 1 0 12972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_131
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_147
timestamp 0
transform 1 0 15548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_159
timestamp 0
transform 1 0 16652 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_165
timestamp 0
transform 1 0 17204 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 3404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 5612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_69
timestamp 0
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_81
timestamp 0
transform 1 0 9476 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_89
timestamp 0
transform 1 0 10212 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_95
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_107
timestamp 0
transform 1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 0
transform 1 0 12420 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_122
timestamp 0
transform 1 0 13248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_130
timestamp 0
transform 1 0 13984 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_146
timestamp 0
transform 1 0 15456 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_158
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 0
transform 1 0 17296 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 0
transform 1 0 17572 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 3404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 4692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_41
timestamp 0
transform 1 0 5796 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_49
timestamp 0
transform 1 0 6532 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_56
timestamp 0
transform 1 0 7176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_68
timestamp 0
transform 1 0 8280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_79
timestamp 0
transform 1 0 9292 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 0
transform 1 0 9844 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_109
timestamp 0
transform 1 0 12052 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_129
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_149
timestamp 0
transform 1 0 15732 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_161
timestamp 0
transform 1 0 16836 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_165
timestamp 0
transform 1 0 17204 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_13
timestamp 0
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_25
timestamp 0
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_37
timestamp 0
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 0
transform 1 0 8004 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_88
timestamp 0
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_98
timestamp 0
transform 1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_108
timestamp 0
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 12420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_125
timestamp 0
transform 1 0 13524 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_133
timestamp 0
transform 1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_146
timestamp 0
transform 1 0 15456 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_158
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 0
transform 1 0 17572 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_6
timestamp 0
transform 1 0 2576 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 0
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_53
timestamp 0
transform 1 0 6900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_62
timestamp 0
transform 1 0 7728 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_70
timestamp 0
transform 1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_79
timestamp 0
transform 1 0 9292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 0
transform 1 0 9844 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_93
timestamp 0
transform 1 0 10580 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_98
timestamp 0
transform 1 0 11040 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_110
timestamp 0
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_118
timestamp 0
transform 1 0 12880 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_124
timestamp 0
transform 1 0 13432 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14996 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 0
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_165
timestamp 0
transform 1 0 17204 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_7
timestamp 0
transform 1 0 2668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_19
timestamp 0
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_31
timestamp 0
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_43
timestamp 0
transform 1 0 5980 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 7268 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_81
timestamp 0
transform 1 0 9476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_90
timestamp 0
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_107
timestamp 0
transform 1 0 11868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_135
timestamp 0
transform 1 0 14444 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_147
timestamp 0
transform 1 0 15548 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_159
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_163
timestamp 0
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 0
transform 1 0 17572 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 3404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 4692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_41
timestamp 0
transform 1 0 5796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_54
timestamp 0
transform 1 0 6992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_60
timestamp 0
transform 1 0 7544 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 0
transform 1 0 9476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 0
transform 1 0 9844 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_94
timestamp 0
transform 1 0 10672 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_106
timestamp 0
transform 1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_115
timestamp 0
transform 1 0 12604 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_127
timestamp 0
transform 1 0 13708 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_165
timestamp 0
transform 1 0 17204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_169
timestamp 0
transform 1 0 17572 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_7
timestamp 0
transform 1 0 2668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_19
timestamp 0
transform 1 0 3772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_31
timestamp 0
transform 1 0 4876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_43
timestamp 0
transform 1 0 5980 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 7268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_69
timestamp 0
transform 1 0 8372 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 10580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 11684 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 0
transform 1 0 12420 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_119
timestamp 0
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_128
timestamp 0
transform 1 0 13800 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_140
timestamp 0
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_152
timestamp 0
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_156
timestamp 0
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 0
transform 1 0 17572 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 3404 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 4692 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 5796 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 0
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_65
timestamp 0
transform 1 0 8004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_69
timestamp 0
transform 1 0 8372 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 0
transform 1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 0
transform 1 0 9844 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_101
timestamp 0
transform 1 0 11316 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_113
timestamp 0
transform 1 0 12420 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_128
timestamp 0
transform 1 0 13800 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 0
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_165
timestamp 0
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_169
timestamp 0
transform 1 0 17572 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 0
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 0
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 0
transform 1 0 5612 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_76
timestamp 0
transform 1 0 9016 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_92
timestamp 0
transform 1 0 10488 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 0
transform 1 0 11868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 13524 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 0
transform 1 0 14628 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 0
transform 1 0 15732 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 0
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 0
transform 1 0 17572 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 3404 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 4692 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 8004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 9108 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_85
timestamp 0
transform 1 0 9844 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_98
timestamp 0
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_110
timestamp 0
transform 1 0 12144 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_122
timestamp 0
transform 1 0 13248 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 0
transform 1 0 14352 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 0
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_165
timestamp 0
transform 1 0 17204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_169
timestamp 0
transform 1 0 17572 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 2300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 3404 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 5612 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 7268 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 8372 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 9476 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 10580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 11684 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 12420 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 15732 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 16836 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 0
transform 1 0 17572 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 3404 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 4692 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 5796 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 0
transform 1 0 6900 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 0
transform 1 0 8004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 0
transform 1 0 9108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 9844 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 13156 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 14260 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_165
timestamp 0
transform 1 0 17204 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_169
timestamp 0
transform 1 0 17572 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 0
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 0
transform 1 0 5612 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 6716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 7268 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 8372 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 9476 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 10580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 11684 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 0
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 0
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 0
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 15732 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 16836 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_169
timestamp 0
transform 1 0 17572 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 2300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 3404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 4692 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 5796 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 0
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 0
transform 1 0 8004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 0
transform 1 0 9108 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 9844 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 0
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 0
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 13156 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 14260 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14996 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 0
transform 1 0 16100 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_165
timestamp 0
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_169
timestamp 0
transform 1 0 17572 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 0
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 0
transform 1 0 5612 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 0
transform 1 0 6716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 7084 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 7268 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 0
transform 1 0 8372 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 0
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 0
transform 1 0 10580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 0
transform 1 0 11684 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 12420 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 13524 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 0
transform 1 0 14628 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 0
transform 1 0 15732 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 0
transform 1 0 16836 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_169
timestamp 0
transform 1 0 17572 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 2300 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 3404 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 4692 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 0
transform 1 0 5796 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_53
timestamp 0
transform 1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_57
timestamp 0
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_69
timestamp 0
transform 1 0 8372 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 0
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_89
timestamp 0
transform 1 0 10212 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_95
timestamp 0
transform 1 0 10764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_102
timestamp 0
transform 1 0 11408 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_109
timestamp 0
transform 1 0 12052 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_117
timestamp 0
transform 1 0 12788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_129
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 0
transform 1 0 14628 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 14996 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 0
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_165
timestamp 0
transform 1 0 17204 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_169
timestamp 0
transform 1 0 17572 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 0
transform 1 0 9844 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 0
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 0
transform -1 0 17664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 0
transform -1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 0
transform -1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 0
transform 1 0 11684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 0
transform 1 0 9844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 0
transform 1 0 2300 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 0
transform 1 0 12420 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 0
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 0
transform -1 0 17664 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 0
transform -1 0 17480 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 0
transform -1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 0
transform 1 0 9108 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 0
transform 1 0 2300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 0
transform 1 0 7820 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 0
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 0
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 0
transform -1 0 10764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 0
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 0
transform 1 0 17296 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 0
transform -1 0 12788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 0
transform -1 0 10764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 0
transform -1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 0
transform -1 0 2668 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_29
timestamp 0
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 17940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_30
timestamp 0
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 17940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_31
timestamp 0
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_32
timestamp 0
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 17940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_33
timestamp 0
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_34
timestamp 0
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 17940 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_35
timestamp 0
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_36
timestamp 0
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_37
timestamp 0
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_38
timestamp 0
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 17940 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_39
timestamp 0
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_40
timestamp 0
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_41
timestamp 0
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_42
timestamp 0
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 17940 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_43
timestamp 0
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 17940 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_44
timestamp 0
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 17940 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_45
timestamp 0
transform 1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 17940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_46
timestamp 0
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 17940 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_47
timestamp 0
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_48
timestamp 0
transform 1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 17940 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_49
timestamp 0
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 17940 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_50
timestamp 0
transform 1 0 2024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 17940 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_51
timestamp 0
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 17940 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_52
timestamp 0
transform 1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 17940 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_53
timestamp 0
transform 1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 17940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_54
timestamp 0
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 17940 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_55
timestamp 0
transform 1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 17940 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_56
timestamp 0
transform 1 0 2024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 17940 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_57
timestamp 0
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 17940 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 0
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 0
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 0
transform 1 0 9752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 0
transform 1 0 12328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 0
transform 1 0 14904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 0
transform 1 0 17480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 0
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_65
timestamp 0
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_66
timestamp 0
transform 1 0 17480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 0
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_68
timestamp 0
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_69
timestamp 0
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 0
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_71
timestamp 0
transform 1 0 12328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_72
timestamp 0
transform 1 0 17480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 0
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_74
timestamp 0
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp 0
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 0
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp 0
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp 0
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 0
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp 0
transform 1 0 9752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp 0
transform 1 0 14904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 0
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp 0
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp 0
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 0
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_86
timestamp 0
transform 1 0 9752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp 0
transform 1 0 14904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 0
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp 0
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_90
timestamp 0
transform 1 0 17480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 0
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp 0
transform 1 0 9752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp 0
transform 1 0 14904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 0
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_95
timestamp 0
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp 0
transform 1 0 17480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 0
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_98
timestamp 0
transform 1 0 9752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_99
timestamp 0
transform 1 0 14904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 0
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_101
timestamp 0
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_102
timestamp 0
transform 1 0 17480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 0
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_104
timestamp 0
transform 1 0 9752 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_105
timestamp 0
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 0
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_107
timestamp 0
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_108
timestamp 0
transform 1 0 17480 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 0
transform 1 0 4600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_110
timestamp 0
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_111
timestamp 0
transform 1 0 14904 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 0
transform 1 0 7176 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_113
timestamp 0
transform 1 0 12328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_114
timestamp 0
transform 1 0 17480 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 0
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_116
timestamp 0
transform 1 0 9752 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_117
timestamp 0
transform 1 0 14904 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 0
transform 1 0 7176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_119
timestamp 0
transform 1 0 12328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_120
timestamp 0
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 0
transform 1 0 4600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_122
timestamp 0
transform 1 0 9752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_123
timestamp 0
transform 1 0 14904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 0
transform 1 0 7176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_125
timestamp 0
transform 1 0 12328 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_126
timestamp 0
transform 1 0 17480 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 0
transform 1 0 4600 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_128
timestamp 0
transform 1 0 9752 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_129
timestamp 0
transform 1 0 14904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 0
transform 1 0 7176 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_131
timestamp 0
transform 1 0 12328 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_132
timestamp 0
transform 1 0 17480 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 0
transform 1 0 4600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_134
timestamp 0
transform 1 0 9752 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_135
timestamp 0
transform 1 0 14904 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 0
transform 1 0 7176 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_137
timestamp 0
transform 1 0 12328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_138
timestamp 0
transform 1 0 17480 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 0
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_140
timestamp 0
transform 1 0 9752 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_141
timestamp 0
transform 1 0 14904 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 0
transform 1 0 7176 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 0
transform 1 0 12328 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 0
transform 1 0 17480 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_145
timestamp 0
transform 1 0 4600 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_146
timestamp 0
transform 1 0 7176 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_147
timestamp 0
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_148
timestamp 0
transform 1 0 12328 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 0
transform 1 0 14904 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 0
transform 1 0 17480 0 1 17408
box -38 -48 130 592
<< labels >>
rlabel metal1 s 9982 17408 9982 17408 4 VGND
rlabel metal1 s 9982 17952 9982 17952 4 VPWR
rlabel metal2 s 9062 1622 9062 1622 4 A[0]
rlabel metal2 s 10994 1588 10994 1588 4 A[1]
rlabel metal3 s 17526 8891 17526 8891 4 A[2]
rlabel metal2 s 17434 10455 17434 10455 4 A[3]
rlabel metal2 s 17526 10999 17526 10999 4 A[4]
rlabel metal1 s 11684 17646 11684 17646 4 A[5]
rlabel metal1 s 9844 17646 9844 17646 4 A[6]
rlabel metal3 s 912 10268 912 10268 4 A[7]
rlabel metal2 s 12282 1588 12282 1588 4 B[0]
rlabel metal2 s 11638 1554 11638 1554 4 B[1]
rlabel metal2 s 17618 7701 17618 7701 4 B[2]
rlabel metal2 s 17342 11679 17342 11679 4 B[3]
rlabel metal1 s 16468 12750 16468 12750 4 B[4]
rlabel metal1 s 11132 17646 11132 17646 4 B[5]
rlabel metal1 s 9154 17646 9154 17646 4 B[6]
rlabel metal3 s 1510 10948 1510 10948 4 B[7]
rlabel metal2 s 13018 13702 13018 13702 4 _000_
rlabel metal1 s 11086 13804 11086 13804 4 _001_
rlabel metal1 s 14674 9588 14674 9588 4 _002_
rlabel metal1 s 11362 13940 11362 13940 4 _003_
rlabel metal1 s 12328 13838 12328 13838 4 _004_
rlabel metal2 s 13478 11526 13478 11526 4 _005_
rlabel metal2 s 13202 12036 13202 12036 4 _006_
rlabel metal2 s 11086 10438 11086 10438 4 _007_
rlabel metal2 s 13110 11254 13110 11254 4 _008_
rlabel metal2 s 12282 12036 12282 12036 4 _009_
rlabel metal2 s 13846 12070 13846 12070 4 _010_
rlabel metal1 s 10304 13294 10304 13294 4 _011_
rlabel metal2 s 11270 13668 11270 13668 4 _012_
rlabel metal1 s 10764 13226 10764 13226 4 _013_
rlabel metal1 s 10902 13770 10902 13770 4 _014_
rlabel metal2 s 11546 14246 11546 14246 4 _015_
rlabel metal1 s 11316 14246 11316 14246 4 _016_
rlabel metal2 s 10902 11526 10902 11526 4 _017_
rlabel metal1 s 11362 11764 11362 11764 4 _018_
rlabel metal1 s 10672 9690 10672 9690 4 _019_
rlabel metal2 s 10258 10438 10258 10438 4 _020_
rlabel metal1 s 11132 10778 11132 10778 4 _021_
rlabel metal2 s 9338 12036 9338 12036 4 _022_
rlabel metal1 s 9246 12784 9246 12784 4 _023_
rlabel metal1 s 9246 13328 9246 13328 4 _024_
rlabel metal1 s 9062 13294 9062 13294 4 _025_
rlabel metal1 s 8556 13498 8556 13498 4 _026_
rlabel metal1 s 10718 13328 10718 13328 4 _027_
rlabel metal2 s 11178 13668 11178 13668 4 _028_
rlabel metal2 s 9522 13668 9522 13668 4 _029_
rlabel metal1 s 9062 13770 9062 13770 4 _030_
rlabel metal1 s 9430 10676 9430 10676 4 _031_
rlabel metal2 s 8786 10540 8786 10540 4 _032_
rlabel metal1 s 8326 10574 8326 10574 4 _033_
rlabel metal2 s 8602 10234 8602 10234 4 _034_
rlabel metal1 s 9108 10234 9108 10234 4 _035_
rlabel metal2 s 6762 12988 6762 12988 4 _036_
rlabel metal1 s 7314 11084 7314 11084 4 _037_
rlabel metal1 s 7820 12342 7820 12342 4 _038_
rlabel metal1 s 6900 12750 6900 12750 4 _039_
rlabel metal1 s 7222 12410 7222 12410 4 _040_
rlabel metal1 s 7130 10234 7130 10234 4 _041_
rlabel metal1 s 7130 10642 7130 10642 4 _042_
rlabel metal1 s 7084 10778 7084 10778 4 _043_
rlabel metal2 s 7682 11798 7682 11798 4 _044_
rlabel metal2 s 8418 6477 8418 6477 4 _045_
rlabel metal1 s 9108 9146 9108 9146 4 _046_
rlabel metal1 s 9246 6732 9246 6732 4 _047_
rlabel metal1 s 8188 7378 8188 7378 4 _048_
rlabel metal1 s 10074 6222 10074 6222 4 _049_
rlabel metal2 s 8326 6732 8326 6732 4 _050_
rlabel metal2 s 8050 6460 8050 6460 4 _051_
rlabel metal1 s 8832 6426 8832 6426 4 _052_
rlabel metal2 s 13156 10030 13156 10030 4 _053_
rlabel metal1 s 12903 9962 12903 9962 4 _054_
rlabel metal2 s 9062 7582 9062 7582 4 _055_
rlabel metal2 s 7774 7650 7774 7650 4 _056_
rlabel metal2 s 9890 10812 9890 10812 4 _057_
rlabel metal2 s 8970 6970 8970 6970 4 _058_
rlabel metal1 s 9568 6766 9568 6766 4 _059_
rlabel metal1 s 7360 8942 7360 8942 4 _060_
rlabel metal2 s 13386 8602 13386 8602 4 _061_
rlabel metal1 s 8924 9146 8924 9146 4 _062_
rlabel metal1 s 14398 6664 14398 6664 4 _063_
rlabel metal2 s 12006 6460 12006 6460 4 _064_
rlabel metal2 s 11178 6460 11178 6460 4 _065_
rlabel metal1 s 10764 6290 10764 6290 4 _066_
rlabel metal1 s 11546 6358 11546 6358 4 _067_
rlabel metal1 s 10396 6222 10396 6222 4 _068_
rlabel metal1 s 10350 6426 10350 6426 4 _069_
rlabel metal1 s 12926 9520 12926 9520 4 _070_
rlabel metal2 s 7682 6970 7682 6970 4 _071_
rlabel metal1 s 13064 11050 13064 11050 4 _072_
rlabel metal1 s 10994 7888 10994 7888 4 _073_
rlabel metal2 s 11270 8160 11270 8160 4 _074_
rlabel metal1 s 11086 8364 11086 8364 4 _075_
rlabel metal2 s 12466 11407 12466 11407 4 _076_
rlabel metal1 s 12052 10030 12052 10030 4 _077_
rlabel metal1 s 10442 8500 10442 8500 4 _078_
rlabel metal1 s 10994 8432 10994 8432 4 _079_
rlabel metal1 s 10442 7922 10442 7922 4 _080_
rlabel metal1 s 13524 7854 13524 7854 4 _081_
rlabel metal2 s 13846 8262 13846 8262 4 _082_
rlabel metal1 s 13386 8058 13386 8058 4 _083_
rlabel metal1 s 12466 8432 12466 8432 4 _084_
rlabel metal1 s 13478 8364 13478 8364 4 _085_
rlabel metal1 s 12098 6358 12098 6358 4 _086_
rlabel metal1 s 14766 8466 14766 8466 4 _087_
rlabel metal1 s 13570 6766 13570 6766 4 _088_
rlabel metal1 s 14352 7174 14352 7174 4 _089_
rlabel metal2 s 14858 7174 14858 7174 4 _090_
rlabel metal2 s 14398 7582 14398 7582 4 _091_
rlabel metal1 s 15272 8942 15272 8942 4 _092_
rlabel metal2 s 14766 7684 14766 7684 4 _093_
rlabel metal2 s 14766 8942 14766 8942 4 _094_
rlabel metal1 s 14030 8398 14030 8398 4 _095_
rlabel metal2 s 13938 9316 13938 9316 4 _096_
rlabel metal1 s 14536 10642 14536 10642 4 _097_
rlabel metal1 s 15042 10642 15042 10642 4 _098_
rlabel metal2 s 15042 10234 15042 10234 4 _099_
rlabel metal1 s 14858 10064 14858 10064 4 _100_
rlabel metal1 s 14996 9554 14996 9554 4 _101_
rlabel metal2 s 15502 9316 15502 9316 4 _102_
rlabel metal1 s 14398 9350 14398 9350 4 _103_
rlabel metal1 s 13202 9962 13202 9962 4 _104_
rlabel metal1 s 12788 9554 12788 9554 4 _105_
rlabel metal1 s 11546 9996 11546 9996 4 _106_
rlabel metal1 s 11454 9996 11454 9996 4 _107_
rlabel metal1 s 12650 9622 12650 9622 4 _108_
rlabel metal1 s 13432 12818 13432 12818 4 _109_
rlabel metal1 s 13570 13294 13570 13294 4 _110_
rlabel metal1 s 13386 13328 13386 13328 4 _111_
rlabel metal1 s 11776 13838 11776 13838 4 _112_
rlabel metal1 s 10120 6766 10120 6766 4 net1
rlabel metal1 s 12098 2550 12098 2550 4 net10
rlabel metal1 s 15916 6766 15916 6766 4 net11
rlabel metal2 s 14858 11356 14858 11356 4 net12
rlabel metal1 s 13202 12852 13202 12852 4 net13
rlabel metal1 s 11270 17510 11270 17510 4 net14
rlabel metal2 s 9430 14926 9430 14926 4 net15
rlabel metal2 s 5934 10914 5934 10914 4 net16
rlabel metal1 s 8050 6902 8050 6902 4 net17
rlabel metal1 s 8970 2618 8970 2618 4 net18
rlabel metal1 s 4922 8874 4922 8874 4 net19
rlabel metal1 s 12558 8398 12558 8398 4 net2
rlabel metal1 s 9476 2414 9476 2414 4 net20
rlabel metal2 s 10718 5372 10718 5372 4 net21
rlabel metal1 s 17158 8398 17158 8398 4 net22
rlabel metal1 s 13892 9622 13892 9622 4 net23
rlabel metal1 s 12788 17646 12788 17646 4 net24
rlabel metal1 s 11086 17578 11086 17578 4 net25
rlabel metal2 s 8694 11526 8694 11526 4 net26
rlabel metal1 s 2622 12852 2622 12852 4 net27
rlabel metal1 s 13984 7854 13984 7854 4 net3
rlabel metal1 s 15410 10540 15410 10540 4 net4
rlabel metal1 s 13754 13294 13754 13294 4 net5
rlabel metal1 s 11270 17782 11270 17782 4 net6
rlabel metal1 s 9752 12818 9752 12818 4 net7
rlabel metal1 s 6256 10642 6256 10642 4 net8
rlabel metal1 s 12788 2482 12788 2482 4 net9
rlabel metal2 s 7774 1588 7774 1588 4 opcode[0]
rlabel metal2 s 8418 1588 8418 1588 4 opcode[1]
rlabel metal3 s 958 8908 958 8908 4 opcode[2]
rlabel metal2 s 9706 1520 9706 1520 4 out[0]
rlabel metal1 s 10442 2822 10442 2822 4 out[1]
rlabel metal2 s 17342 8279 17342 8279 4 out[2]
rlabel metal2 s 17526 9741 17526 9741 4 out[3]
rlabel metal2 s 12282 18540 12282 18540 4 out[4]
rlabel metal1 s 10442 17850 10442 17850 4 out[5]
rlabel metal3 s 958 11628 958 11628 4 out[6]
rlabel metal3 s 1556 12308 1556 12308 4 out[7]
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 A[0]
port 1 nsew
flabel metal2 s 10966 0 11022 800 0 FreeSans 280 90 0 0 A[1]
port 2 nsew
flabel metal3 s 19200 8848 20000 8968 0 FreeSans 600 0 0 0 A[2]
port 3 nsew
flabel metal3 s 19200 10208 20000 10328 0 FreeSans 600 0 0 0 A[3]
port 4 nsew
flabel metal3 s 19200 10888 20000 11008 0 FreeSans 600 0 0 0 A[4]
port 5 nsew
flabel metal2 s 11610 19200 11666 20000 0 FreeSans 280 90 0 0 A[5]
port 6 nsew
flabel metal2 s 9678 19200 9734 20000 0 FreeSans 280 90 0 0 A[6]
port 7 nsew
flabel metal3 s 0 10208 800 10328 0 FreeSans 600 0 0 0 A[7]
port 8 nsew
flabel metal2 s 12254 0 12310 800 0 FreeSans 280 90 0 0 B[0]
port 9 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 B[1]
port 10 nsew
flabel metal3 s 19200 7488 20000 7608 0 FreeSans 600 0 0 0 B[2]
port 11 nsew
flabel metal3 s 19200 11568 20000 11688 0 FreeSans 600 0 0 0 B[3]
port 12 nsew
flabel metal3 s 19200 12248 20000 12368 0 FreeSans 600 0 0 0 B[4]
port 13 nsew
flabel metal2 s 10966 19200 11022 20000 0 FreeSans 280 90 0 0 B[5]
port 14 nsew
flabel metal2 s 9034 19200 9090 20000 0 FreeSans 280 90 0 0 B[6]
port 15 nsew
flabel metal3 s 0 10888 800 11008 0 FreeSans 600 0 0 0 B[7]
port 16 nsew
flabel metal5 s 1976 16480 17988 16800 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal5 s 1976 12536 17988 12856 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal5 s 1976 8592 17988 8912 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal5 s 1976 4648 17988 4968 0 FreeSans 3200 0 0 0 VGND
port 17 nsew
flabel metal4 s 16450 2128 16770 18000 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 12471 2128 12791 18000 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 8492 2128 8812 18000 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal4 s 4513 2128 4833 18000 0 FreeSans 2400 90 0 0 VGND
port 17 nsew
flabel metal5 s 1976 15820 17988 16140 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal5 s 1976 11876 17988 12196 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal5 s 1976 7932 17988 8252 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal5 s 1976 3988 17988 4308 0 FreeSans 3200 0 0 0 VPWR
port 18 nsew
flabel metal4 s 15790 2128 16110 18000 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 11811 2128 12131 18000 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 7832 2128 8152 18000 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal4 s 3853 2128 4173 18000 0 FreeSans 2400 90 0 0 VPWR
port 18 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 opcode[0]
port 19 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 opcode[1]
port 20 nsew
flabel metal3 s 0 8848 800 8968 0 FreeSans 600 0 0 0 opcode[2]
port 21 nsew
flabel metal2 s 9678 0 9734 800 0 FreeSans 280 90 0 0 out[0]
port 22 nsew
flabel metal2 s 10322 0 10378 800 0 FreeSans 280 90 0 0 out[1]
port 23 nsew
flabel metal3 s 19200 8168 20000 8288 0 FreeSans 600 0 0 0 out[2]
port 24 nsew
flabel metal3 s 19200 9528 20000 9648 0 FreeSans 600 0 0 0 out[3]
port 25 nsew
flabel metal2 s 12254 19200 12310 20000 0 FreeSans 280 90 0 0 out[4]
port 26 nsew
flabel metal2 s 10322 19200 10378 20000 0 FreeSans 280 90 0 0 out[5]
port 27 nsew
flabel metal3 s 0 11568 800 11688 0 FreeSans 600 0 0 0 out[6]
port 28 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 out[7]
port 29 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
