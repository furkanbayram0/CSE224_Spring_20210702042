magic
tech sky130A
magscale 1 2
timestamp 1747874834
<< nwell >>
rect 1066 2159 78882 77830
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 842 2128 78844 77840
<< metal2 >>
rect 28354 79200 28410 80000
rect 30930 79200 30986 80000
rect 31574 79200 31630 80000
rect 32218 79200 32274 80000
rect 34794 79200 34850 80000
rect 38014 79200 38070 80000
rect 44454 79200 44510 80000
rect 45098 79200 45154 80000
rect 45742 79200 45798 80000
rect 46386 79200 46442 80000
rect 7746 0 7802 800
rect 18050 0 18106 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 35438 0 35494 800
rect 37370 0 37426 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 45098 0 45154 800
rect 48318 0 48374 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 53470 0 53526 800
rect 55402 0 55458 800
rect 61842 0 61898 800
rect 62486 0 62542 800
rect 63130 0 63186 800
rect 63774 0 63830 800
<< obsm2 >>
rect 846 79144 28298 79200
rect 28466 79144 30874 79200
rect 31042 79144 31518 79200
rect 31686 79144 32162 79200
rect 32330 79144 34738 79200
rect 34906 79144 37958 79200
rect 38126 79144 44398 79200
rect 44566 79144 45042 79200
rect 45210 79144 45686 79200
rect 45854 79144 46330 79200
rect 46498 79144 78550 79200
rect 846 856 78550 79144
rect 846 734 7690 856
rect 7858 734 17994 856
rect 18162 734 27654 856
rect 27822 734 28942 856
rect 29110 734 29586 856
rect 29754 734 30230 856
rect 30398 734 31518 856
rect 31686 734 32162 856
rect 32330 734 32806 856
rect 32974 734 33450 856
rect 33618 734 35382 856
rect 35550 734 37314 856
rect 37482 734 42466 856
rect 42634 734 43754 856
rect 43922 734 45042 856
rect 45210 734 48262 856
rect 48430 734 48906 856
rect 49074 734 50194 856
rect 50362 734 53414 856
rect 53582 734 55346 856
rect 55514 734 61786 856
rect 61954 734 62430 856
rect 62598 734 63074 856
rect 63242 734 63718 856
rect 63886 734 78550 856
<< metal3 >>
rect 79200 53728 80000 53848
rect 79200 53048 80000 53168
rect 79200 52368 80000 52488
rect 79200 51688 80000 51808
rect 0 51008 800 51128
rect 79200 51008 80000 51128
rect 79200 50328 80000 50448
rect 79200 49648 80000 49768
rect 79200 48968 80000 49088
rect 79200 48288 80000 48408
rect 79200 47608 80000 47728
rect 0 46928 800 47048
rect 79200 46928 80000 47048
rect 79200 46248 80000 46368
rect 0 45568 800 45688
rect 79200 45568 80000 45688
rect 0 44888 800 45008
rect 79200 44888 80000 45008
rect 0 44208 800 44328
rect 79200 44208 80000 44328
rect 0 43528 800 43648
rect 79200 43528 80000 43648
rect 0 42848 800 42968
rect 79200 42848 80000 42968
rect 0 42168 800 42288
rect 79200 42168 80000 42288
rect 0 41488 800 41608
rect 79200 41488 80000 41608
rect 0 40808 800 40928
rect 79200 40808 80000 40928
rect 79200 40128 80000 40248
rect 79200 39448 80000 39568
rect 79200 38768 80000 38888
rect 0 38088 800 38208
rect 79200 38088 80000 38208
rect 79200 37408 80000 37528
rect 79200 36728 80000 36848
rect 79200 36048 80000 36168
rect 0 35368 800 35488
rect 79200 35368 80000 35488
rect 79200 34688 80000 34808
rect 79200 34008 80000 34128
rect 0 33328 800 33448
rect 79200 33328 80000 33448
rect 79200 32648 80000 32768
rect 79200 31968 80000 32088
rect 79200 31288 80000 31408
rect 0 29928 800 30048
rect 79200 28568 80000 28688
<< obsm3 >>
rect 798 53928 79200 77825
rect 798 53648 79120 53928
rect 798 53248 79200 53648
rect 798 52968 79120 53248
rect 798 52568 79200 52968
rect 798 52288 79120 52568
rect 798 51888 79200 52288
rect 798 51608 79120 51888
rect 798 51208 79200 51608
rect 880 50928 79120 51208
rect 798 50528 79200 50928
rect 798 50248 79120 50528
rect 798 49848 79200 50248
rect 798 49568 79120 49848
rect 798 49168 79200 49568
rect 798 48888 79120 49168
rect 798 48488 79200 48888
rect 798 48208 79120 48488
rect 798 47808 79200 48208
rect 798 47528 79120 47808
rect 798 47128 79200 47528
rect 880 46848 79120 47128
rect 798 46448 79200 46848
rect 798 46168 79120 46448
rect 798 45768 79200 46168
rect 880 45488 79120 45768
rect 798 45088 79200 45488
rect 880 44808 79120 45088
rect 798 44408 79200 44808
rect 880 44128 79120 44408
rect 798 43728 79200 44128
rect 880 43448 79120 43728
rect 798 43048 79200 43448
rect 880 42768 79120 43048
rect 798 42368 79200 42768
rect 880 42088 79120 42368
rect 798 41688 79200 42088
rect 880 41408 79120 41688
rect 798 41008 79200 41408
rect 880 40728 79120 41008
rect 798 40328 79200 40728
rect 798 40048 79120 40328
rect 798 39648 79200 40048
rect 798 39368 79120 39648
rect 798 38968 79200 39368
rect 798 38688 79120 38968
rect 798 38288 79200 38688
rect 880 38008 79120 38288
rect 798 37608 79200 38008
rect 798 37328 79120 37608
rect 798 36928 79200 37328
rect 798 36648 79120 36928
rect 798 36248 79200 36648
rect 798 35968 79120 36248
rect 798 35568 79200 35968
rect 880 35288 79120 35568
rect 798 34888 79200 35288
rect 798 34608 79120 34888
rect 798 34208 79200 34608
rect 798 33928 79120 34208
rect 798 33528 79200 33928
rect 880 33248 79120 33528
rect 798 32848 79200 33248
rect 798 32568 79120 32848
rect 798 32168 79200 32568
rect 798 31888 79120 32168
rect 798 31488 79200 31888
rect 798 31208 79120 31488
rect 798 30128 79200 31208
rect 880 29848 79200 30128
rect 798 28768 79200 29848
rect 798 28488 79120 28768
rect 798 2143 79200 28488
<< metal4 >>
rect 1944 2128 2264 77840
rect 2604 2128 2924 77840
rect 6944 2128 7264 77840
rect 7604 2128 7924 77840
rect 11944 2128 12264 77840
rect 12604 2128 12924 77840
rect 16944 2128 17264 77840
rect 17604 2128 17924 77840
rect 21944 2128 22264 77840
rect 22604 2128 22924 77840
rect 26944 2128 27264 77840
rect 27604 2128 27924 77840
rect 31944 2128 32264 77840
rect 32604 2128 32924 77840
rect 36944 2128 37264 77840
rect 37604 2128 37924 77840
rect 41944 2128 42264 77840
rect 42604 2128 42924 77840
rect 46944 2128 47264 77840
rect 47604 2128 47924 77840
rect 51944 2128 52264 77840
rect 52604 2128 52924 77840
rect 56944 2128 57264 77840
rect 57604 2128 57924 77840
rect 61944 2128 62264 77840
rect 62604 2128 62924 77840
rect 66944 2128 67264 77840
rect 67604 2128 67924 77840
rect 71944 2128 72264 77840
rect 72604 2128 72924 77840
rect 76944 2128 77264 77840
rect 77604 2128 77924 77840
<< obsm4 >>
rect 11283 2619 11864 77349
rect 12344 2619 12524 77349
rect 13004 2619 16864 77349
rect 17344 2619 17524 77349
rect 18004 2619 21864 77349
rect 22344 2619 22524 77349
rect 23004 2619 26864 77349
rect 27344 2619 27524 77349
rect 28004 2619 31864 77349
rect 32344 2619 32524 77349
rect 33004 2619 36864 77349
rect 37344 2619 37524 77349
rect 38004 2619 41864 77349
rect 42344 2619 42524 77349
rect 43004 2619 46864 77349
rect 47344 2619 47524 77349
rect 48004 2619 51864 77349
rect 52344 2619 52524 77349
rect 53004 2619 56864 77349
rect 57344 2619 57524 77349
rect 58004 2619 61864 77349
rect 62344 2619 62524 77349
rect 63004 2619 66864 77349
rect 67344 2619 67524 77349
rect 68004 2619 71864 77349
rect 72344 2619 72437 77349
<< metal5 >>
rect 1056 73676 78892 73996
rect 1056 73016 78892 73336
rect 1056 68676 78892 68996
rect 1056 68016 78892 68336
rect 1056 63676 78892 63996
rect 1056 63016 78892 63336
rect 1056 58676 78892 58996
rect 1056 58016 78892 58336
rect 1056 53676 78892 53996
rect 1056 53016 78892 53336
rect 1056 48676 78892 48996
rect 1056 48016 78892 48336
rect 1056 43676 78892 43996
rect 1056 43016 78892 43336
rect 1056 38676 78892 38996
rect 1056 38016 78892 38336
rect 1056 33676 78892 33996
rect 1056 33016 78892 33336
rect 1056 28676 78892 28996
rect 1056 28016 78892 28336
rect 1056 23676 78892 23996
rect 1056 23016 78892 23336
rect 1056 18676 78892 18996
rect 1056 18016 78892 18336
rect 1056 13676 78892 13996
rect 1056 13016 78892 13336
rect 1056 8676 78892 8996
rect 1056 8016 78892 8336
rect 1056 3676 78892 3996
rect 1056 3016 78892 3336
<< obsm5 >>
rect 29372 16500 48276 16820
<< labels >>
rlabel metal2 s 62486 0 62542 800 6 A1[0]
port 1 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 A1[1]
port 2 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 A1[2]
port 3 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 A1[3]
port 4 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 A1[4]
port 5 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 A2[0]
port 6 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 A2[1]
port 7 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 A2[2]
port 8 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 A2[3]
port 9 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 A2[4]
port 10 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 A3[0]
port 11 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 A3[1]
port 12 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 A3[2]
port 13 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 A3[3]
port 14 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 A3[4]
port 15 nsew signal input
rlabel metal3 s 79200 31288 80000 31408 6 ALU_result[0]
port 16 nsew signal output
rlabel metal3 s 79200 32648 80000 32768 6 ALU_result[10]
port 17 nsew signal output
rlabel metal3 s 79200 53728 80000 53848 6 ALU_result[11]
port 18 nsew signal output
rlabel metal3 s 79200 40128 80000 40248 6 ALU_result[12]
port 19 nsew signal output
rlabel metal3 s 79200 40808 80000 40928 6 ALU_result[13]
port 20 nsew signal output
rlabel metal3 s 79200 39448 80000 39568 6 ALU_result[14]
port 21 nsew signal output
rlabel metal3 s 79200 46248 80000 46368 6 ALU_result[15]
port 22 nsew signal output
rlabel metal3 s 79200 42168 80000 42288 6 ALU_result[16]
port 23 nsew signal output
rlabel metal3 s 79200 42848 80000 42968 6 ALU_result[17]
port 24 nsew signal output
rlabel metal3 s 79200 43528 80000 43648 6 ALU_result[18]
port 25 nsew signal output
rlabel metal3 s 79200 47608 80000 47728 6 ALU_result[19]
port 26 nsew signal output
rlabel metal3 s 79200 37408 80000 37528 6 ALU_result[1]
port 27 nsew signal output
rlabel metal3 s 79200 44888 80000 45008 6 ALU_result[20]
port 28 nsew signal output
rlabel metal3 s 79200 46928 80000 47048 6 ALU_result[21]
port 29 nsew signal output
rlabel metal3 s 79200 44208 80000 44328 6 ALU_result[22]
port 30 nsew signal output
rlabel metal3 s 79200 53048 80000 53168 6 ALU_result[23]
port 31 nsew signal output
rlabel metal3 s 79200 45568 80000 45688 6 ALU_result[24]
port 32 nsew signal output
rlabel metal3 s 79200 48968 80000 49088 6 ALU_result[25]
port 33 nsew signal output
rlabel metal3 s 79200 48288 80000 48408 6 ALU_result[26]
port 34 nsew signal output
rlabel metal3 s 79200 52368 80000 52488 6 ALU_result[27]
port 35 nsew signal output
rlabel metal3 s 79200 51008 80000 51128 6 ALU_result[28]
port 36 nsew signal output
rlabel metal3 s 79200 50328 80000 50448 6 ALU_result[29]
port 37 nsew signal output
rlabel metal3 s 79200 36048 80000 36168 6 ALU_result[2]
port 38 nsew signal output
rlabel metal3 s 79200 51688 80000 51808 6 ALU_result[30]
port 39 nsew signal output
rlabel metal3 s 79200 49648 80000 49768 6 ALU_result[31]
port 40 nsew signal output
rlabel metal3 s 79200 38088 80000 38208 6 ALU_result[3]
port 41 nsew signal output
rlabel metal3 s 79200 33328 80000 33448 6 ALU_result[4]
port 42 nsew signal output
rlabel metal3 s 79200 38768 80000 38888 6 ALU_result[5]
port 43 nsew signal output
rlabel metal3 s 79200 34008 80000 34128 6 ALU_result[6]
port 44 nsew signal output
rlabel metal3 s 79200 35368 80000 35488 6 ALU_result[7]
port 45 nsew signal output
rlabel metal3 s 79200 41488 80000 41608 6 ALU_result[8]
port 46 nsew signal output
rlabel metal3 s 79200 31968 80000 32088 6 ALU_result[9]
port 47 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 CLK
port 48 nsew signal input
rlabel metal4 s 2604 2128 2924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 22604 2128 22924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 27604 2128 27924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 32604 2128 32924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 37604 2128 37924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 42604 2128 42924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 47604 2128 47924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 52604 2128 52924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 57604 2128 57924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 62604 2128 62924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 67604 2128 67924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 72604 2128 72924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 77604 2128 77924 77840 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 3676 78892 3996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 8676 78892 8996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 13676 78892 13996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 18676 78892 18996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 23676 78892 23996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 28676 78892 28996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 33676 78892 33996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 38676 78892 38996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 43676 78892 43996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 48676 78892 48996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 53676 78892 53996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 58676 78892 58996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 63676 78892 63996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 68676 78892 68996 6 VGND
port 49 nsew ground bidirectional
rlabel metal5 s 1056 73676 78892 73996 6 VGND
port 49 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 21944 2128 22264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 26944 2128 27264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 31944 2128 32264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 36944 2128 37264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 41944 2128 42264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 46944 2128 47264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 51944 2128 52264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 56944 2128 57264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 61944 2128 62264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 66944 2128 67264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 71944 2128 72264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal4 s 76944 2128 77264 77840 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 3016 78892 3336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 8016 78892 8336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 13016 78892 13336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 18016 78892 18336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 23016 78892 23336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 28016 78892 28336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 33016 78892 33336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 38016 78892 38336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 43016 78892 43336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 48016 78892 48336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 53016 78892 53336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 58016 78892 58336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 63016 78892 63336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 68016 78892 68336 6 VPWR
port 50 nsew power bidirectional
rlabel metal5 s 1056 73016 78892 73336 6 VPWR
port 50 nsew power bidirectional
rlabel metal2 s 63774 0 63830 800 6 WD3[0]
port 51 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 WD3[10]
port 52 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 WD3[11]
port 53 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 WD3[12]
port 54 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 WD3[13]
port 55 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 WD3[14]
port 56 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 WD3[15]
port 57 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 WD3[16]
port 58 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 WD3[17]
port 59 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 WD3[18]
port 60 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 WD3[19]
port 61 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 WD3[1]
port 62 nsew signal input
rlabel metal2 s 45742 79200 45798 80000 6 WD3[20]
port 63 nsew signal input
rlabel metal2 s 28354 79200 28410 80000 6 WD3[21]
port 64 nsew signal input
rlabel metal2 s 45098 79200 45154 80000 6 WD3[22]
port 65 nsew signal input
rlabel metal2 s 32218 79200 32274 80000 6 WD3[23]
port 66 nsew signal input
rlabel metal2 s 38014 79200 38070 80000 6 WD3[24]
port 67 nsew signal input
rlabel metal2 s 44454 79200 44510 80000 6 WD3[25]
port 68 nsew signal input
rlabel metal2 s 34794 79200 34850 80000 6 WD3[26]
port 69 nsew signal input
rlabel metal2 s 31574 79200 31630 80000 6 WD3[27]
port 70 nsew signal input
rlabel metal2 s 30930 79200 30986 80000 6 WD3[28]
port 71 nsew signal input
rlabel metal2 s 46386 79200 46442 80000 6 WD3[29]
port 72 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 WD3[2]
port 73 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 WD3[30]
port 74 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 WD3[31]
port 75 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 WD3[3]
port 76 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 WD3[4]
port 77 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 WD3[5]
port 78 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 WD3[6]
port 79 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 WD3[7]
port 80 nsew signal input
rlabel metal3 s 79200 28568 80000 28688 6 WD3[8]
port 81 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 WD3[9]
port 82 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 WE3
port 83 nsew signal input
rlabel metal3 s 79200 36728 80000 36848 6 opcode[0]
port 84 nsew signal input
rlabel metal3 s 79200 34688 80000 34808 6 opcode[1]
port 85 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17878966
string GDS_FILE /openlane/designs/project4/runs/RUN_2025.05.22_00.40.45/results/signoff/project4.magic.gds
string GDS_START 778696
<< end >>

