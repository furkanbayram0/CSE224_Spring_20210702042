magic
tech sky130A
magscale 1 2
timestamp 1745718354
<< nwell >>
rect 1066 2159 6846 9809
<< obsli1 >>
rect 1104 2159 6808 9809
<< obsm1 >>
rect 842 2128 6808 9840
<< obsm2 >>
rect 846 711 6512 10985
<< metal3 >>
rect 0 10888 800 11008
rect 0 10208 800 10328
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
rect 0 7488 800 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 0 5448 800 5568
rect 0 4768 800 4888
rect 0 4088 800 4208
rect 0 3408 800 3528
rect 0 2728 800 2848
rect 0 2048 800 2168
rect 0 1368 800 1488
rect 0 688 800 808
<< obsm3 >>
rect 880 10808 2922 10981
rect 798 10408 2922 10808
rect 880 10128 2922 10408
rect 798 9728 2922 10128
rect 880 9448 2922 9728
rect 798 9048 2922 9448
rect 880 8768 2922 9048
rect 798 8368 2922 8768
rect 880 8088 2922 8368
rect 798 7688 2922 8088
rect 880 7408 2922 7688
rect 798 7008 2922 7408
rect 880 6728 2922 7008
rect 798 6328 2922 6728
rect 880 6048 2922 6328
rect 798 5648 2922 6048
rect 880 5368 2922 5648
rect 798 4968 2922 5368
rect 880 4688 2922 4968
rect 798 4288 2922 4688
rect 880 4008 2922 4288
rect 798 3608 2922 4008
rect 880 3328 2922 3608
rect 798 2928 2922 3328
rect 880 2648 2922 2928
rect 798 2248 2922 2648
rect 880 1968 2922 2248
rect 798 1568 2922 1968
rect 880 1288 2922 1568
rect 798 888 2922 1288
rect 880 715 2922 888
<< metal4 >>
rect 1944 2128 2264 9840
rect 2604 2128 2924 9840
<< labels >>
rlabel metal4 s 2604 2128 2924 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 688 800 808 6 in[0]
port 3 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 in[1]
port 4 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 in[2]
port 5 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 in[3]
port 6 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 in[4]
port 7 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 in[5]
port 8 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 in[6]
port 9 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 in[7]
port 10 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 out[0]
port 11 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 out[1]
port 12 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 out[2]
port 13 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 out[3]
port 14 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 out[4]
port 15 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 out[5]
port 16 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 out[6]
port 17 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 out[7]
port 18 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 8000 12000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 186224
string GDS_FILE /openlane/designs/project1/runs/RUN_2025.04.27_01.45.23/results/signoff/project1.magic.gds
string GDS_START 96222
<< end >>

