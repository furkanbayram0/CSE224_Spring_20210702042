VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO project3
  CLASS BLOCK ;
  FOREIGN project3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 90.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.020 10.640 39.620 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.020 10.640 64.620 79.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.380 74.300 19.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.380 74.300 44.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 68.380 74.300 69.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 10.640 36.320 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.720 10.640 61.320 79.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.080 74.300 16.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.080 74.300 41.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 65.080 74.300 66.680 ;
    END
  END VPWR
  PIN an0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 43.560 80.000 44.160 ;
    END
  END an0
  PIN an1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 49.000 80.000 49.600 ;
    END
  END an1
  PIN an2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 54.440 80.000 55.040 ;
    END
  END an2
  PIN an3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 59.880 80.000 60.480 ;
    END
  END an3
  PIN an4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 65.320 80.000 65.920 ;
    END
  END an4
  PIN an5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 70.760 80.000 71.360 ;
    END
  END an5
  PIN an6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 76.200 80.000 76.800 ;
    END
  END an6
  PIN an7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 81.640 80.000 82.240 ;
    END
  END an7
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END rst
  PIN seg0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 76.000 5.480 80.000 6.080 ;
    END
  END seg0
  PIN seg1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 76.000 10.920 80.000 11.520 ;
    END
  END seg1
  PIN seg2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 76.000 16.360 80.000 16.960 ;
    END
  END seg2
  PIN seg3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 76.000 21.800 80.000 22.400 ;
    END
  END seg3
  PIN seg4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 76.000 27.240 80.000 27.840 ;
    END
  END seg4
  PIN seg5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 76.000 32.680 80.000 33.280 ;
    END
  END seg5
  PIN seg6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 76.000 38.120 80.000 38.720 ;
    END
  END seg6
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 74.250 79.070 ;
      LAYER li1 ;
        RECT 5.520 10.795 74.060 78.965 ;
      LAYER met1 ;
        RECT 3.290 8.200 78.590 79.860 ;
      LAYER met2 ;
        RECT 3.320 5.595 78.560 82.125 ;
      LAYER met3 ;
        RECT 3.030 81.240 75.600 82.105 ;
        RECT 3.030 77.200 76.000 81.240 ;
        RECT 3.030 75.800 75.600 77.200 ;
        RECT 3.030 71.760 76.000 75.800 ;
        RECT 3.030 70.360 75.600 71.760 ;
        RECT 3.030 67.680 76.000 70.360 ;
        RECT 4.400 66.320 76.000 67.680 ;
        RECT 4.400 66.280 75.600 66.320 ;
        RECT 3.030 64.920 75.600 66.280 ;
        RECT 3.030 60.880 76.000 64.920 ;
        RECT 3.030 59.480 75.600 60.880 ;
        RECT 3.030 55.440 76.000 59.480 ;
        RECT 3.030 54.040 75.600 55.440 ;
        RECT 3.030 50.000 76.000 54.040 ;
        RECT 3.030 48.600 75.600 50.000 ;
        RECT 3.030 44.560 76.000 48.600 ;
        RECT 3.030 43.160 75.600 44.560 ;
        RECT 3.030 39.120 76.000 43.160 ;
        RECT 3.030 37.720 75.600 39.120 ;
        RECT 3.030 33.680 76.000 37.720 ;
        RECT 3.030 32.280 75.600 33.680 ;
        RECT 3.030 28.240 76.000 32.280 ;
        RECT 3.030 26.840 75.600 28.240 ;
        RECT 3.030 22.800 76.000 26.840 ;
        RECT 4.400 21.400 75.600 22.800 ;
        RECT 3.030 17.360 76.000 21.400 ;
        RECT 3.030 15.960 75.600 17.360 ;
        RECT 3.030 11.920 76.000 15.960 ;
        RECT 3.030 10.520 75.600 11.920 ;
        RECT 3.030 6.480 76.000 10.520 ;
        RECT 3.030 5.615 75.600 6.480 ;
      LAYER met4 ;
        RECT 3.055 10.240 9.320 77.345 ;
        RECT 11.720 10.240 12.620 77.345 ;
        RECT 15.020 10.240 34.320 77.345 ;
        RECT 36.720 10.240 37.620 77.345 ;
        RECT 40.020 10.240 59.320 77.345 ;
        RECT 61.720 10.240 62.620 77.345 ;
        RECT 65.020 10.240 70.545 77.345 ;
        RECT 3.055 7.655 70.545 10.240 ;
  END
END project3
END LIBRARY

