VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO project2
  CLASS BLOCK ;
  FOREIGN project2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 44.240 100.000 44.840 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 51.040 100.000 51.640 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 54.440 100.000 55.040 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 96.000 58.330 100.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END A[7]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 37.440 100.000 38.040 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 57.840 100.000 58.440 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 96.000 61.240 100.000 61.840 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 96.000 55.110 100.000 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 96.000 45.450 100.000 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END B[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 22.565 10.640 24.165 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.460 10.640 44.060 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.355 10.640 63.955 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.250 10.640 83.850 90.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 23.240 89.940 24.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 42.960 89.940 44.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 62.680 89.940 64.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 82.400 89.940 84.000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.265 10.640 20.865 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.160 10.640 40.760 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.055 10.640 60.655 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.950 10.640 80.550 90.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 19.940 89.940 21.540 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 39.660 89.940 41.260 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 59.380 89.940 60.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 79.100 89.940 80.700 ;
    END
  END VPWR
  PIN opcode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END opcode[0]
  PIN opcode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END opcode[1]
  PIN opcode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END opcode[2]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 40.840 100.000 41.440 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 96.000 61.550 100.000 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 96.000 51.890 100.000 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END out[7]
  OBS
      LAYER nwell ;
        RECT 9.930 10.795 89.890 89.950 ;
      LAYER li1 ;
        RECT 10.120 10.795 89.700 89.845 ;
      LAYER met1 ;
        RECT 5.590 10.640 89.700 90.000 ;
      LAYER met2 ;
        RECT 5.610 95.720 44.890 96.000 ;
        RECT 45.730 95.720 48.110 96.000 ;
        RECT 48.950 95.720 51.330 96.000 ;
        RECT 52.170 95.720 54.550 96.000 ;
        RECT 55.390 95.720 57.770 96.000 ;
        RECT 58.610 95.720 60.990 96.000 ;
        RECT 61.830 95.720 88.230 96.000 ;
        RECT 5.610 4.280 88.230 95.720 ;
        RECT 5.610 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 88.230 4.280 ;
      LAYER met3 ;
        RECT 4.000 62.240 96.000 89.925 ;
        RECT 4.400 60.840 95.600 62.240 ;
        RECT 4.000 58.840 96.000 60.840 ;
        RECT 4.400 57.440 95.600 58.840 ;
        RECT 4.000 55.440 96.000 57.440 ;
        RECT 4.400 54.040 95.600 55.440 ;
        RECT 4.000 52.040 96.000 54.040 ;
        RECT 4.400 50.640 95.600 52.040 ;
        RECT 4.000 48.640 96.000 50.640 ;
        RECT 4.000 47.240 95.600 48.640 ;
        RECT 4.000 45.240 96.000 47.240 ;
        RECT 4.400 43.840 95.600 45.240 ;
        RECT 4.000 41.840 96.000 43.840 ;
        RECT 4.000 40.440 95.600 41.840 ;
        RECT 4.000 38.440 96.000 40.440 ;
        RECT 4.000 37.040 95.600 38.440 ;
        RECT 4.000 10.715 96.000 37.040 ;
  END
END project2
END LIBRARY

