magic
tech sky130A
magscale 1 2
timestamp 1748900824
<< nwell >>
rect 1066 2159 58918 57681
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 1104 2128 58880 57712
<< obsm2 >>
rect 1950 2139 58586 57701
<< metal3 >>
rect 59200 55224 60000 55344
rect 59200 53592 60000 53712
rect 59200 51960 60000 52080
rect 59200 50328 60000 50448
rect 0 49784 800 49904
rect 59200 48696 60000 48816
rect 59200 47064 60000 47184
rect 59200 45432 60000 45552
rect 59200 43800 60000 43920
rect 59200 42168 60000 42288
rect 59200 40536 60000 40656
rect 59200 38904 60000 39024
rect 59200 37272 60000 37392
rect 59200 35640 60000 35760
rect 59200 34008 60000 34128
rect 59200 32376 60000 32496
rect 59200 30744 60000 30864
rect 0 29928 800 30048
rect 59200 29112 60000 29232
rect 59200 27480 60000 27600
rect 59200 25848 60000 25968
rect 59200 24216 60000 24336
rect 59200 22584 60000 22704
rect 59200 20952 60000 21072
rect 59200 19320 60000 19440
rect 59200 17688 60000 17808
rect 59200 16056 60000 16176
rect 59200 14424 60000 14544
rect 59200 12792 60000 12912
rect 59200 11160 60000 11280
rect 0 10072 800 10192
rect 59200 9528 60000 9648
rect 59200 7896 60000 8016
rect 59200 6264 60000 6384
rect 59200 4632 60000 4752
<< obsm3 >>
rect 1946 55424 59200 57697
rect 1946 55144 59120 55424
rect 1946 53792 59200 55144
rect 1946 53512 59120 53792
rect 1946 52160 59200 53512
rect 1946 51880 59120 52160
rect 1946 50528 59200 51880
rect 1946 50248 59120 50528
rect 1946 48896 59200 50248
rect 1946 48616 59120 48896
rect 1946 47264 59200 48616
rect 1946 46984 59120 47264
rect 1946 45632 59200 46984
rect 1946 45352 59120 45632
rect 1946 44000 59200 45352
rect 1946 43720 59120 44000
rect 1946 42368 59200 43720
rect 1946 42088 59120 42368
rect 1946 40736 59200 42088
rect 1946 40456 59120 40736
rect 1946 39104 59200 40456
rect 1946 38824 59120 39104
rect 1946 37472 59200 38824
rect 1946 37192 59120 37472
rect 1946 35840 59200 37192
rect 1946 35560 59120 35840
rect 1946 34208 59200 35560
rect 1946 33928 59120 34208
rect 1946 32576 59200 33928
rect 1946 32296 59120 32576
rect 1946 30944 59200 32296
rect 1946 30664 59120 30944
rect 1946 29312 59200 30664
rect 1946 29032 59120 29312
rect 1946 27680 59200 29032
rect 1946 27400 59120 27680
rect 1946 26048 59200 27400
rect 1946 25768 59120 26048
rect 1946 24416 59200 25768
rect 1946 24136 59120 24416
rect 1946 22784 59200 24136
rect 1946 22504 59120 22784
rect 1946 21152 59200 22504
rect 1946 20872 59120 21152
rect 1946 19520 59200 20872
rect 1946 19240 59120 19520
rect 1946 17888 59200 19240
rect 1946 17608 59120 17888
rect 1946 16256 59200 17608
rect 1946 15976 59120 16256
rect 1946 14624 59200 15976
rect 1946 14344 59120 14624
rect 1946 12992 59200 14344
rect 1946 12712 59120 12992
rect 1946 11360 59200 12712
rect 1946 11080 59120 11360
rect 1946 9728 59200 11080
rect 1946 9448 59120 9728
rect 1946 8096 59200 9448
rect 1946 7816 59120 8096
rect 1946 6464 59200 7816
rect 1946 6184 59120 6464
rect 1946 4832 59200 6184
rect 1946 4552 59120 4832
rect 1946 2143 59200 4552
<< metal4 >>
rect 1944 2128 2264 57712
rect 2604 2128 2924 57712
rect 6944 2128 7264 57712
rect 7604 2128 7924 57712
rect 11944 2128 12264 57712
rect 12604 2128 12924 57712
rect 16944 2128 17264 57712
rect 17604 2128 17924 57712
rect 21944 2128 22264 57712
rect 22604 2128 22924 57712
rect 26944 2128 27264 57712
rect 27604 2128 27924 57712
rect 31944 2128 32264 57712
rect 32604 2128 32924 57712
rect 36944 2128 37264 57712
rect 37604 2128 37924 57712
rect 41944 2128 42264 57712
rect 42604 2128 42924 57712
rect 46944 2128 47264 57712
rect 47604 2128 47924 57712
rect 51944 2128 52264 57712
rect 52604 2128 52924 57712
rect 56944 2128 57264 57712
rect 57604 2128 57924 57712
<< metal5 >>
rect 1056 53676 58928 53996
rect 1056 53016 58928 53336
rect 1056 48676 58928 48996
rect 1056 48016 58928 48336
rect 1056 43676 58928 43996
rect 1056 43016 58928 43336
rect 1056 38676 58928 38996
rect 1056 38016 58928 38336
rect 1056 33676 58928 33996
rect 1056 33016 58928 33336
rect 1056 28676 58928 28996
rect 1056 28016 58928 28336
rect 1056 23676 58928 23996
rect 1056 23016 58928 23336
rect 1056 18676 58928 18996
rect 1056 18016 58928 18336
rect 1056 13676 58928 13996
rect 1056 13016 58928 13336
rect 1056 8676 58928 8996
rect 1056 8016 58928 8336
rect 1056 3676 58928 3996
rect 1056 3016 58928 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 22604 2128 22924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27604 2128 27924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 32604 2128 32924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37604 2128 37924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42604 2128 42924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47604 2128 47924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 52604 2128 52924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 57604 2128 57924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 58928 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8676 58928 8996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13676 58928 13996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18676 58928 18996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 23676 58928 23996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 28676 58928 28996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 33676 58928 33996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 38676 58928 38996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 43676 58928 43996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 48676 58928 48996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 53676 58928 53996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 21944 2128 22264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26944 2128 27264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 31944 2128 32264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 36944 2128 37264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 41944 2128 42264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46944 2128 47264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 51944 2128 52264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 56944 2128 57264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 58928 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8016 58928 8336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13016 58928 13336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 18016 58928 18336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 23016 58928 23336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 28016 58928 28336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 33016 58928 33336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 38016 58928 38336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 43016 58928 43336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 48016 58928 48336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 53016 58928 53336 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 10072 800 10192 6 clk
port 3 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 control
port 4 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 reset
port 5 nsew signal input
rlabel metal3 s 59200 55224 60000 55344 6 result[0]
port 6 nsew signal output
rlabel metal3 s 59200 38904 60000 39024 6 result[10]
port 7 nsew signal output
rlabel metal3 s 59200 37272 60000 37392 6 result[11]
port 8 nsew signal output
rlabel metal3 s 59200 35640 60000 35760 6 result[12]
port 9 nsew signal output
rlabel metal3 s 59200 34008 60000 34128 6 result[13]
port 10 nsew signal output
rlabel metal3 s 59200 32376 60000 32496 6 result[14]
port 11 nsew signal output
rlabel metal3 s 59200 30744 60000 30864 6 result[15]
port 12 nsew signal output
rlabel metal3 s 59200 29112 60000 29232 6 result[16]
port 13 nsew signal output
rlabel metal3 s 59200 27480 60000 27600 6 result[17]
port 14 nsew signal output
rlabel metal3 s 59200 25848 60000 25968 6 result[18]
port 15 nsew signal output
rlabel metal3 s 59200 24216 60000 24336 6 result[19]
port 16 nsew signal output
rlabel metal3 s 59200 53592 60000 53712 6 result[1]
port 17 nsew signal output
rlabel metal3 s 59200 22584 60000 22704 6 result[20]
port 18 nsew signal output
rlabel metal3 s 59200 20952 60000 21072 6 result[21]
port 19 nsew signal output
rlabel metal3 s 59200 19320 60000 19440 6 result[22]
port 20 nsew signal output
rlabel metal3 s 59200 17688 60000 17808 6 result[23]
port 21 nsew signal output
rlabel metal3 s 59200 16056 60000 16176 6 result[24]
port 22 nsew signal output
rlabel metal3 s 59200 14424 60000 14544 6 result[25]
port 23 nsew signal output
rlabel metal3 s 59200 12792 60000 12912 6 result[26]
port 24 nsew signal output
rlabel metal3 s 59200 11160 60000 11280 6 result[27]
port 25 nsew signal output
rlabel metal3 s 59200 9528 60000 9648 6 result[28]
port 26 nsew signal output
rlabel metal3 s 59200 7896 60000 8016 6 result[29]
port 27 nsew signal output
rlabel metal3 s 59200 51960 60000 52080 6 result[2]
port 28 nsew signal output
rlabel metal3 s 59200 6264 60000 6384 6 result[30]
port 29 nsew signal output
rlabel metal3 s 59200 4632 60000 4752 6 result[31]
port 30 nsew signal output
rlabel metal3 s 59200 50328 60000 50448 6 result[3]
port 31 nsew signal output
rlabel metal3 s 59200 48696 60000 48816 6 result[4]
port 32 nsew signal output
rlabel metal3 s 59200 47064 60000 47184 6 result[5]
port 33 nsew signal output
rlabel metal3 s 59200 45432 60000 45552 6 result[6]
port 34 nsew signal output
rlabel metal3 s 59200 43800 60000 43920 6 result[7]
port 35 nsew signal output
rlabel metal3 s 59200 42168 60000 42288 6 result[8]
port 36 nsew signal output
rlabel metal3 s 59200 40536 60000 40656 6 result[9]
port 37 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1954416
string GDS_FILE /openlane/designs/project5/runs/RUN_2025.06.02_21.46.29/results/signoff/top_module.magic.gds
string GDS_START 22340
<< end >>

