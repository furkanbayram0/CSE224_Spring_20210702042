* NGSPICE file created from project3.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

.subckt project3 VGND VPWR an7 clk rst seg0 seg1 seg2 seg3 seg4 seg5 seg6 an6 an5
+ an4 an3 an2 an1 an0
XANTENNA__203__B _075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_294_ decoder.digit\[1\] _155_ _067_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__a21boi_1
XANTENNA__304__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_346_ clknet_2_0__leaf_clk _007_ _044_ VGND VGND VPWR VPWR one_second_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_277_ one_second_counter\[24\] _127_ _148_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__and3_1
X_200_ _075_ _085_ _093_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__and3b_1
XFILLER_0_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__171__A2 decoder.digit\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_329_ net1 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__211__B _100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__312__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__307__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__217__A one_second_counter\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput7 net7 VGND VGND VPWR VPWR seg5 sky130_fd_sc_hd__buf_1
XFILLER_0_2_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_293_ _158_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__320__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__230__A one_second_counter\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_276_ _127_ _148_ one_second_counter\[24\] VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__a21oi_1
X_345_ clknet_2_2__leaf_clk _006_ _043_ VGND VGND VPWR VPWR one_second_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__315__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__225__A _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_328_ net1 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__inv_2
X_259_ _136_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xproject3_10 VGND VGND VPWR VPWR an0 project3_10/LO sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_12_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__323__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__217__B _077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput8 net8 VGND VGND VPWR VPWR seg6 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_2_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__318__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_361_ clknet_2_2__leaf_clk _063_ _059_ VGND VGND VPWR VPWR decoder.digit\[3\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_15_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_292_ decoder.digit\[3\] decoder.digit\[1\] _156_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__230__B _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_275_ _147_ _145_ _148_ _127_ _027_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a221oi_2
X_344_ clknet_2_1__leaf_clk _005_ _042_ VGND VGND VPWR VPWR one_second_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__174__A1 one_second_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__241__A _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__209__C _100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_327_ _161_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_189_ _086_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__buf_2
XANTENNA__326__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_258_ _127_ _135_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__236__A _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xproject3_11 VGND VGND VPWR VPWR an1 project3_11/LO sky130_fd_sc_hd__conb_1
XFILLER_0_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_291_ _157_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_360_ clknet_2_2__leaf_clk _062_ _058_ VGND VGND VPWR VPWR decoder.digit\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__228__B one_second_counter\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__186__C1 one_second_counter\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__329__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_274_ _083_ _135_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__and2_1
X_343_ clknet_2_0__leaf_clk _004_ _041_ VGND VGND VPWR VPWR one_second_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__174__A2 decoder.digit\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_257_ one_second_counter\[19\] one_second_counter\[18\] one_second_counter\[17\]
+ one_second_counter\[16\] VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__and4_1
X_188_ _085_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__inv_2
X_326_ _161_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xproject3_12 VGND VGND VPWR VPWR an2 project3_12/LO sky130_fd_sc_hd__conb_1
X_309_ _160_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__162__A one_second_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__260__A _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_290_ decoder.digit\[3\] decoder.digit\[2\] decoder.digit\[0\] VGND VGND VPWR VPWR
+ _157_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__244__B one_second_counter\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__256__A4 _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_342_ clknet_2_1__leaf_clk _003_ _040_ VGND VGND VPWR VPWR one_second_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_273_ one_second_counter\[23\] VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__inv_2
XANTENNA__165__A decoder.digit\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_187_ _073_ _084_ one_second_counter\[26\] VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__a21bo_2
X_256_ one_second_counter\[18\] one_second_counter\[17\] one_second_counter\[16\]
+ _127_ one_second_counter\[19\] VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__a41o_1
X_325_ _161_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__inv_2
Xproject3_13 VGND VGND VPWR VPWR an3 project3_13/LO sky130_fd_sc_hd__conb_1
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__162__B decoder.digit\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_308_ _160_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__inv_2
X_239_ _121_ _119_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__nand2_1
XANTENNA__247__B _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__258__A _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__244__C _078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_272_ _146_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__clkbuf_1
X_341_ clknet_2_1__leaf_clk _002_ _039_ VGND VGND VPWR VPWR one_second_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__165__B decoder.digit\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__271__A _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_324_ _161_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__inv_2
X_186_ _074_ _082_ _083_ one_second_counter\[24\] VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__o211ai_2
X_255_ _132_ _129_ _133_ _095_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xproject3_14 VGND VGND VPWR VPWR an4 project3_14/LO sky130_fd_sc_hd__conb_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload1 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_307_ _160_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__inv_2
X_238_ one_second_counter\[14\] VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__inv_2
X_169_ _065_ _069_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__and2_1
XANTENNA__162__C decoder.digit\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__179__A _075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__186__A2 _082_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ clknet_2_3__leaf_clk _001_ _038_ VGND VGND VPWR VPWR one_second_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_20_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_271_ _085_ _144_ _145_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__and3_1
XANTENNA__181__B one_second_counter\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_254_ one_second_counter\[17\] one_second_counter\[16\] _127_ one_second_counter\[18\]
+ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__a31o_1
X_323_ _161_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__inv_2
X_185_ one_second_counter\[23\] one_second_counter\[22\] one_second_counter\[20\]
+ one_second_counter\[21\] VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__192__A one_second_counter\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xproject3_15 VGND VGND VPWR VPWR an5 project3_15/LO sky130_fd_sc_hd__conb_1
Xclkload2 clknet_2_3__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__277__A one_second_counter\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_168_ one_second_enable _068_ _064_ decoder.digit\[2\] VGND VGND VPWR VPWR _069_
+ sky130_fd_sc_hd__o2bb2a_1
X_306_ net1 VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__buf_4
X_237_ _120_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__289__A1 decoder.digit\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__290__A decoder.digit\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__285__A decoder.digit\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_270_ one_second_counter\[22\] _143_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_322_ _161_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__inv_2
X_184_ one_second_counter\[8\] _077_ _079_ _081_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__o31a_1
XFILLER_0_19_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_253_ one_second_counter\[18\] one_second_counter\[17\] VGND VGND VPWR VPWR _132_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__192__B one_second_counter\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xproject3_16 VGND VGND VPWR VPWR an6 project3_16/LO sky130_fd_sc_hd__conb_1
XFILLER_0_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_305_ _159_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__277__B _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_236_ _095_ _118_ _119_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__and3_1
X_167_ decoder.digit\[0\] _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__nor2_1
XANTENNA__289__A2 _155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__288__A _068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_219_ _107_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__buf_1
XFILLER_0_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__195__B one_second_counter\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__181__D _078_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__296__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__234__B1 one_second_counter\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_321_ _161_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ one_second_counter\[17\] one_second_counter\[16\] _080_ one_second_counter\[18\]
+ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__and4b_1
X_252_ _027_ _131_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_235_ one_second_counter\[12\] one_second_counter\[13\] _114_ VGND VGND VPWR VPWR
+ _119_ sky130_fd_sc_hd__nand3_2
X_304_ _159_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_166_ decoder.digit\[2\] _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_218_ _105_ _085_ _106_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__288__B _155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__290__C decoder.digit\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__299__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__195__C one_second_counter\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_182_ one_second_counter\[19\] one_second_counter\[13\] one_second_counter\[14\]
+ one_second_counter\[15\] VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__and4b_1
X_320_ _161_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__inv_2
X_251_ one_second_counter\[17\] _129_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__234__A1 one_second_counter\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_234_ one_second_counter\[12\] _114_ one_second_counter\[13\] VGND VGND VPWR VPWR
+ _118_ sky130_fd_sc_hd__a21o_1
X_165_ decoder.digit\[3\] decoder.digit\[1\] VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_303_ _159_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__inv_2
X_217_ one_second_counter\[8\] _077_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__255__C1 _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_181_ one_second_counter\[11\] one_second_counter\[10\] one_second_counter\[9\] _078_
+ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_13_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_250_ _130_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__234__A2 _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _159_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__inv_2
X_233_ _117_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__207__A2 _075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_164_ decoder.digit\[3\] _065_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ one_second_counter\[8\] _077_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__246__B1 _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ one_second_counter\[15\] one_second_counter\[14\] one_second_counter\[12\]
+ one_second_counter\[13\] VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_13_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_301_ _159_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__inv_2
X_232_ _095_ _115_ _116_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__and3_1
X_163_ decoder.digit\[2\] _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nand2_1
XANTENNA__302__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__212__A _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_215_ _104_ _102_ _086_ _077_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__310__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__204__B _075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__305__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__173__B1 decoder.digit\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_162_ one_second_enable decoder.digit\[1\] decoder.digit\[0\] VGND VGND VPWR VPWR
+ _064_ sky130_fd_sc_hd__and3_1
X_231_ one_second_counter\[12\] _114_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__nand2_1
X_300_ _159_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
Xinput1 rst VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_10_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_214_ one_second_counter\[7\] VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__313__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__223__A one_second_counter\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__308__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__321__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__173__A1 one_second_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__231__A one_second_counter\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__316__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__226__A _112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_230_ one_second_counter\[12\] _114_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_359_ clknet_2_2__leaf_clk _061_ _057_ VGND VGND VPWR VPWR decoder.digit\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_213_ _103_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__276__B1 one_second_counter\[24\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__218__B _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__324__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xproject3_9 VGND VGND VPWR VPWR project3_9/HI an7 sky130_fd_sc_hd__conb_1
XANTENNA__319__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__231__B _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_358_ clknet_2_1__leaf_clk _060_ _056_ VGND VGND VPWR VPWR decoder.digit\[0\] sky130_fd_sc_hd__dfrtp_4
X_289_ decoder.digit\[0\] _155_ _066_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__a21oi_1
XANTENNA__327__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_212_ _095_ _101_ _102_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_6_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__294__A1 decoder.digit\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__276__A1 _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_288_ _068_ _155_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__nor2_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_357_ clknet_2_0__leaf_clk _027_ _055_ VGND VGND VPWR VPWR one_second_enable sky130_fd_sc_hd__dfrtp_2
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_211_ one_second_counter\[6\] _100_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__294__A2 _155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__229__C _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_356_ clknet_2_2__leaf_clk _018_ _054_ VGND VGND VPWR VPWR one_second_counter\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_287_ decoder.digit\[2\] decoder.digit\[1\] _068_ _156_ decoder.digit\[3\] VGND VGND
+ VPWR VPWR net2 sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_210_ one_second_counter\[6\] _100_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_339_ clknet_2_0__leaf_clk _026_ _037_ VGND VGND VPWR VPWR one_second_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__248__B _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__264__A _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_286_ decoder.digit\[1\] decoder.digit\[0\] _155_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__and3b_1
X_355_ clknet_2_1__leaf_clk _017_ _053_ VGND VGND VPWR VPWR one_second_counter\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ clknet_2_2__leaf_clk _025_ _036_ VGND VGND VPWR VPWR one_second_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_269_ one_second_counter\[22\] _143_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__370__A net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__280__A one_second_counter\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__190__A one_second_counter\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__168__A1_N one_second_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__182__B one_second_counter\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_354_ clknet_2_3__leaf_clk _016_ _052_ VGND VGND VPWR VPWR one_second_counter\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_285_ decoder.digit\[3\] decoder.digit\[2\] VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__nor2_2
XANTENNA__215__C1 _077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_337_ clknet_2_3__leaf_clk _024_ _035_ VGND VGND VPWR VPWR one_second_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_199_ one_second_counter\[2\] one_second_counter\[1\] one_second_counter\[0\] one_second_counter\[3\]
+ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__a31o_1
XANTENNA__188__A _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_268_ _142_ _140_ _143_ _027_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_370_ net2 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_353_ clknet_2_3__leaf_clk _015_ _051_ VGND VGND VPWR VPWR one_second_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__267__C _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_284_ one_second_counter\[26\] one_second_counter\[25\] _095_ _154_ VGND VGND VPWR
+ VPWR _018_ sky130_fd_sc_hd__o211a_1
XANTENNA__193__B _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__177__C one_second_counter\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_198_ _092_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__clkbuf_1
X_336_ clknet_2_3__leaf_clk _023_ _034_ VGND VGND VPWR VPWR one_second_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_267_ one_second_counter\[20\] one_second_counter\[21\] _127_ _135_ VGND VGND VPWR
+ VPWR _143_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_319_ _161_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__286__B decoder.digit\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__297__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_283_ _073_ _084_ _150_ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__a21o_1
XANTENNA__177__D one_second_counter\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_352_ clknet_2_0__leaf_clk _014_ _050_ VGND VGND VPWR VPWR one_second_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_197_ _090_ _085_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__and3_1
X_335_ clknet_2_1__leaf_clk _022_ _033_ VGND VGND VPWR VPWR one_second_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_266_ one_second_counter\[21\] VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_318_ _161_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_249_ _095_ _128_ _129_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_14_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__286__C _155_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_282_ _153_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__clkbuf_1
X_351_ clknet_2_0__leaf_clk _013_ _049_ VGND VGND VPWR VPWR one_second_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ clknet_2_0__leaf_clk _021_ _032_ VGND VGND VPWR VPWR one_second_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_265_ _141_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_196_ one_second_counter\[1\] one_second_counter\[0\] one_second_counter\[2\] VGND
+ VGND VPWR VPWR _091_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_179_ _075_ _076_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__and2_2
X_248_ one_second_counter\[16\] _127_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__nand2_1
X_317_ net1 VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__buf_4
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_350_ clknet_2_3__leaf_clk _012_ _048_ VGND VGND VPWR VPWR one_second_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_281_ _085_ _151_ _152_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__202__A _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_264_ _085_ _139_ _140_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_333_ clknet_2_1__leaf_clk _020_ _031_ VGND VGND VPWR VPWR one_second_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_195_ one_second_counter\[2\] one_second_counter\[1\] one_second_counter\[0\] VGND
+ VGND VPWR VPWR _090_ sky130_fd_sc_hd__nand3_1
X_316_ _160_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__inv_2
X_247_ one_second_counter\[16\] _127_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_178_ one_second_counter\[7\] one_second_counter\[6\] one_second_counter\[5\] one_second_counter\[4\]
+ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__300__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__227__A1 one_second_counter\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__205__A _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_280_ one_second_counter\[25\] _150_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_263_ one_second_counter\[20\] _136_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__nand2_1
X_194_ _089_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__clkbuf_1
X_332_ clknet_2_1__leaf_clk _019_ _030_ VGND VGND VPWR VPWR one_second_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__303__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__213__A _103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_315_ _160_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__inv_2
X_177_ one_second_counter\[3\] one_second_counter\[2\] one_second_counter\[1\] one_second_counter\[0\]
+ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__and4_2
X_246_ _125_ _123_ _127_ _027_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a211oi_1
X_229_ _027_ _113_ _114_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nor3_1
XANTENNA__210__B _100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__311__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__306__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__216__A one_second_counter\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_262_ one_second_counter\[20\] _136_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__or2_1
X_193_ _087_ _085_ _088_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_331_ clknet_2_1__leaf_clk _011_ _029_ VGND VGND VPWR VPWR one_second_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__284__B1 _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_245_ _126_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__clkbuf_4
X_176_ one_second_counter\[18\] one_second_counter\[17\] one_second_counter\[19\]
+ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__a21o_1
X_314_ _160_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__314__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__224__A one_second_counter\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__309__A _160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__254__A3 _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_228_ one_second_counter\[11\] one_second_counter\[10\] _109_ VGND VGND VPWR VPWR
+ _114_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_9_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__221__B one_second_counter\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__322__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__232__A _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__216__B _077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__317__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_330_ clknet_2_3__leaf_clk _000_ _028_ VGND VGND VPWR VPWR one_second_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__287__D1 decoder.digit\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_261_ _138_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__buf_1
X_192_ one_second_counter\[1\] one_second_counter\[0\] VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_22_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_175_ one_second_counter\[25\] VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__inv_2
X_313_ _160_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__inv_2
X_244_ one_second_counter\[11\] one_second_counter\[10\] _078_ _109_ VGND VGND VPWR
+ VPWR _126_ sky130_fd_sc_hd__and4_1
XANTENNA__275__B2 _127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__208__C _075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_227_ one_second_counter\[10\] _109_ one_second_counter\[11\] VGND VGND VPWR VPWR
+ _113_ sky130_fd_sc_hd__a21oi_1
XANTENNA__235__A one_second_counter\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__325__A _161_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__221__C _075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ _095_ _134_ _137_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__and3_1
X_191_ one_second_counter\[1\] one_second_counter\[0\] VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__284__A2 one_second_counter\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__328__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_312_ _160_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__inv_2
X_174_ one_second_enable decoder.digit\[0\] _072_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__a21oi_1
X_243_ one_second_counter\[15\] VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output4_A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__184__A1 one_second_counter\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_226_ _112_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__235__B one_second_counter\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_209_ _027_ _099_ _100_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__287__B1 _068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_190_ one_second_counter\[0\] _027_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_242_ _124_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__clkbuf_1
X_311_ _160_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__inv_2
X_173_ one_second_enable _067_ decoder.digit\[0\] VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__164__A decoder.digit\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__184__A2 _077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_225_ _095_ _110_ _111_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__and3_1
XANTENNA__249__A _095_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__235__C _114_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_208_ one_second_counter\[5\] one_second_counter\[4\] _075_ VGND VGND VPWR VPWR _100_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__167__A decoder.digit\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__220__A1 one_second_counter\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_310_ _160_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_172_ _064_ _071_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__nor2_1
X_241_ _095_ _122_ _123_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__and3_1
X_224_ one_second_counter\[10\] _109_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__nand2_1
XANTENNA__175__A one_second_counter\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_207_ one_second_counter\[4\] _075_ one_second_counter\[5\] VGND VGND VPWR VPWR _099_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__220__A2 _077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__287__A2 decoder.digit\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__286__A_N decoder.digit\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_171_ one_second_enable decoder.digit\[0\] decoder.digit\[1\] VGND VGND VPWR VPWR
+ _071_ sky130_fd_sc_hd__a21oi_1
X_240_ _121_ _119_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__or2_1
XANTENNA__196__A1 one_second_counter\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_223_ one_second_counter\[10\] _109_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__281__A _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__191__A one_second_counter\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output2_A net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_206_ _098_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__194__A _089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__279__A one_second_counter\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__196__A2 one_second_counter\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_170_ _070_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__180__C one_second_counter\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_299_ _159_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_222_ _027_ _108_ _109_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_8_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__191__B one_second_counter\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_205_ _095_ _096_ _097_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__and3_1
XANTENNA__292__A decoder.digit\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput2 net2 VGND VGND VPWR VPWR seg0 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_24_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__180__D one_second_counter\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_298_ _159_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__inv_2
XANTENNA__295__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_221_ one_second_counter\[9\] one_second_counter\[8\] _075_ _076_ VGND VGND VPWR
+ VPWR _109_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_8_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_204_ one_second_counter\[4\] _075_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__292__B decoder.digit\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__197__B _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__298__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 _069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput3 net3 VGND VGND VPWR VPWR seg1 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_24_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_297_ _159_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_220_ one_second_counter\[8\] _077_ one_second_counter\[9\] VGND VGND VPWR VPWR _108_
+ sky130_fd_sc_hd__a21oi_1
X_349_ clknet_2_2__leaf_clk _010_ _047_ VGND VGND VPWR VPWR one_second_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_203_ one_second_counter\[4\] _075_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_2 _096_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__199__A2 one_second_counter\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput4 net4 VGND VGND VPWR VPWR seg2 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_24_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_21_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_296_ _159_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_348_ clknet_2_2__leaf_clk _009_ _046_ VGND VGND VPWR VPWR one_second_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_279_ one_second_counter\[25\] _150_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_202_ _085_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__buf_2
XANTENNA__171__B1 decoder.digit\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__168__A2_N _068_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 _124_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__200__A_N _075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__199__A3 one_second_counter\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput5 net5 VGND VGND VPWR VPWR seg3 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_24_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_295_ net1 VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__buf_4
X_347_ clknet_2_3__leaf_clk _008_ _045_ VGND VGND VPWR VPWR one_second_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_278_ _027_ _149_ _150_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__nor3_1
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_201_ _094_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__buf_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__200__B _085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__171__A1 one_second_enable VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__301__A _159_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput6 net6 VGND VGND VPWR VPWR seg4 sky130_fd_sc_hd__buf_1
.ends

