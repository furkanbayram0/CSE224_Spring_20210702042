magic
tech sky130A
magscale 1 2
timestamp 1746400030
<< nwell >>
rect 1986 2159 17978 17990
<< obsli1 >>
rect 2024 2159 17940 17969
<< obsm1 >>
rect 1118 2128 17940 18000
<< metal2 >>
rect 9034 19200 9090 20000
rect 9678 19200 9734 20000
rect 10322 19200 10378 20000
rect 10966 19200 11022 20000
rect 11610 19200 11666 20000
rect 12254 19200 12310 20000
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
<< obsm2 >>
rect 1122 19144 8978 19200
rect 9146 19144 9622 19200
rect 9790 19144 10266 19200
rect 10434 19144 10910 19200
rect 11078 19144 11554 19200
rect 11722 19144 12198 19200
rect 12366 19144 17646 19200
rect 1122 856 17646 19144
rect 1122 800 7690 856
rect 7858 800 8334 856
rect 8502 800 8978 856
rect 9146 800 9622 856
rect 9790 800 10266 856
rect 10434 800 10910 856
rect 11078 800 11554 856
rect 11722 800 12198 856
rect 12366 800 17646 856
<< metal3 >>
rect 0 12248 800 12368
rect 19200 12248 20000 12368
rect 0 11568 800 11688
rect 19200 11568 20000 11688
rect 0 10888 800 11008
rect 19200 10888 20000 11008
rect 0 10208 800 10328
rect 19200 10208 20000 10328
rect 19200 9528 20000 9648
rect 0 8848 800 8968
rect 19200 8848 20000 8968
rect 19200 8168 20000 8288
rect 19200 7488 20000 7608
<< obsm3 >>
rect 800 12448 19200 17985
rect 880 12168 19120 12448
rect 800 11768 19200 12168
rect 880 11488 19120 11768
rect 800 11088 19200 11488
rect 880 10808 19120 11088
rect 800 10408 19200 10808
rect 880 10128 19120 10408
rect 800 9728 19200 10128
rect 800 9448 19120 9728
rect 800 9048 19200 9448
rect 880 8768 19120 9048
rect 800 8368 19200 8768
rect 800 8088 19120 8368
rect 800 7688 19200 8088
rect 800 7408 19120 7688
rect 800 2143 19200 7408
<< metal4 >>
rect 3853 2128 4173 18000
rect 4513 2128 4833 18000
rect 7832 2128 8152 18000
rect 8492 2128 8812 18000
rect 11811 2128 12131 18000
rect 12471 2128 12791 18000
rect 15790 2128 16110 18000
rect 16450 2128 16770 18000
<< metal5 >>
rect 1976 16480 17988 16800
rect 1976 15820 17988 16140
rect 1976 12536 17988 12856
rect 1976 11876 17988 12196
rect 1976 8592 17988 8912
rect 1976 7932 17988 8252
rect 1976 4648 17988 4968
rect 1976 3988 17988 4308
<< labels >>
rlabel metal2 s 9034 0 9090 800 6 A[0]
port 1 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 A[1]
port 2 nsew signal input
rlabel metal3 s 19200 8848 20000 8968 6 A[2]
port 3 nsew signal input
rlabel metal3 s 19200 10208 20000 10328 6 A[3]
port 4 nsew signal input
rlabel metal3 s 19200 10888 20000 11008 6 A[4]
port 5 nsew signal input
rlabel metal2 s 11610 19200 11666 20000 6 A[5]
port 6 nsew signal input
rlabel metal2 s 9678 19200 9734 20000 6 A[6]
port 7 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 A[7]
port 8 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 B[0]
port 9 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 B[1]
port 10 nsew signal input
rlabel metal3 s 19200 7488 20000 7608 6 B[2]
port 11 nsew signal input
rlabel metal3 s 19200 11568 20000 11688 6 B[3]
port 12 nsew signal input
rlabel metal3 s 19200 12248 20000 12368 6 B[4]
port 13 nsew signal input
rlabel metal2 s 10966 19200 11022 20000 6 B[5]
port 14 nsew signal input
rlabel metal2 s 9034 19200 9090 20000 6 B[6]
port 15 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 B[7]
port 16 nsew signal input
rlabel metal4 s 4513 2128 4833 18000 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 8492 2128 8812 18000 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 12471 2128 12791 18000 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 16450 2128 16770 18000 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1976 4648 17988 4968 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1976 8592 17988 8912 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1976 12536 17988 12856 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1976 16480 17988 16800 6 VGND
port 17 nsew ground bidirectional
rlabel metal4 s 3853 2128 4173 18000 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 7832 2128 8152 18000 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 11811 2128 12131 18000 6 VPWR
port 18 nsew power bidirectional
rlabel metal4 s 15790 2128 16110 18000 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1976 3988 17988 4308 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1976 7932 17988 8252 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1976 11876 17988 12196 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1976 15820 17988 16140 6 VPWR
port 18 nsew power bidirectional
rlabel metal2 s 7746 0 7802 800 6 opcode[0]
port 19 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 opcode[1]
port 20 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 opcode[2]
port 21 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 out[0]
port 22 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 out[1]
port 23 nsew signal output
rlabel metal3 s 19200 8168 20000 8288 6 out[2]
port 24 nsew signal output
rlabel metal3 s 19200 9528 20000 9648 6 out[3]
port 25 nsew signal output
rlabel metal2 s 12254 19200 12310 20000 6 out[4]
port 26 nsew signal output
rlabel metal2 s 10322 19200 10378 20000 6 out[5]
port 27 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 out[6]
port 28 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 out[7]
port 29 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 741772
string GDS_FILE /openlane/designs/project2/runs/RUN_2025.05.04_23.06.35/results/signoff/project2.magic.gds
string GDS_START 261906
<< end >>

