magic
tech sky130A
magscale 1 2
timestamp 1748901518
<< nwell >>
rect 1066 2159 58918 57681
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 1104 2128 58880 57712
<< obsm2 >>
rect 1950 2139 58586 57701
<< metal3 >>
rect 59200 55496 60000 55616
rect 59200 54680 60000 54800
rect 59200 53864 60000 53984
rect 59200 53048 60000 53168
rect 59200 52232 60000 52352
rect 59200 51416 60000 51536
rect 59200 50600 60000 50720
rect 0 49784 800 49904
rect 59200 49784 60000 49904
rect 59200 48968 60000 49088
rect 59200 48152 60000 48272
rect 59200 47336 60000 47456
rect 59200 46520 60000 46640
rect 59200 45704 60000 45824
rect 59200 44888 60000 45008
rect 59200 44072 60000 44192
rect 59200 43256 60000 43376
rect 59200 42440 60000 42560
rect 59200 41624 60000 41744
rect 59200 40808 60000 40928
rect 59200 39992 60000 40112
rect 59200 39176 60000 39296
rect 59200 38360 60000 38480
rect 59200 37544 60000 37664
rect 59200 36728 60000 36848
rect 59200 35912 60000 36032
rect 59200 35096 60000 35216
rect 59200 34280 60000 34400
rect 59200 33464 60000 33584
rect 59200 32648 60000 32768
rect 59200 31832 60000 31952
rect 59200 31016 60000 31136
rect 59200 30200 60000 30320
rect 0 29928 800 30048
rect 59200 29384 60000 29504
rect 59200 28568 60000 28688
rect 59200 27752 60000 27872
rect 59200 26936 60000 27056
rect 59200 26120 60000 26240
rect 59200 25304 60000 25424
rect 59200 24488 60000 24608
rect 59200 23672 60000 23792
rect 59200 22856 60000 22976
rect 59200 22040 60000 22160
rect 59200 21224 60000 21344
rect 59200 20408 60000 20528
rect 59200 19592 60000 19712
rect 59200 18776 60000 18896
rect 59200 17960 60000 18080
rect 59200 17144 60000 17264
rect 59200 16328 60000 16448
rect 59200 15512 60000 15632
rect 59200 14696 60000 14816
rect 59200 13880 60000 14000
rect 59200 13064 60000 13184
rect 59200 12248 60000 12368
rect 59200 11432 60000 11552
rect 59200 10616 60000 10736
rect 0 10072 800 10192
rect 59200 9800 60000 9920
rect 59200 8984 60000 9104
rect 59200 8168 60000 8288
rect 59200 7352 60000 7472
rect 59200 6536 60000 6656
rect 59200 5720 60000 5840
rect 59200 4904 60000 5024
rect 59200 4088 60000 4208
<< obsm3 >>
rect 1946 55696 59200 57697
rect 1946 55416 59120 55696
rect 1946 54880 59200 55416
rect 1946 54600 59120 54880
rect 1946 54064 59200 54600
rect 1946 53784 59120 54064
rect 1946 53248 59200 53784
rect 1946 52968 59120 53248
rect 1946 52432 59200 52968
rect 1946 52152 59120 52432
rect 1946 51616 59200 52152
rect 1946 51336 59120 51616
rect 1946 50800 59200 51336
rect 1946 50520 59120 50800
rect 1946 49984 59200 50520
rect 1946 49704 59120 49984
rect 1946 49168 59200 49704
rect 1946 48888 59120 49168
rect 1946 48352 59200 48888
rect 1946 48072 59120 48352
rect 1946 47536 59200 48072
rect 1946 47256 59120 47536
rect 1946 46720 59200 47256
rect 1946 46440 59120 46720
rect 1946 45904 59200 46440
rect 1946 45624 59120 45904
rect 1946 45088 59200 45624
rect 1946 44808 59120 45088
rect 1946 44272 59200 44808
rect 1946 43992 59120 44272
rect 1946 43456 59200 43992
rect 1946 43176 59120 43456
rect 1946 42640 59200 43176
rect 1946 42360 59120 42640
rect 1946 41824 59200 42360
rect 1946 41544 59120 41824
rect 1946 41008 59200 41544
rect 1946 40728 59120 41008
rect 1946 40192 59200 40728
rect 1946 39912 59120 40192
rect 1946 39376 59200 39912
rect 1946 39096 59120 39376
rect 1946 38560 59200 39096
rect 1946 38280 59120 38560
rect 1946 37744 59200 38280
rect 1946 37464 59120 37744
rect 1946 36928 59200 37464
rect 1946 36648 59120 36928
rect 1946 36112 59200 36648
rect 1946 35832 59120 36112
rect 1946 35296 59200 35832
rect 1946 35016 59120 35296
rect 1946 34480 59200 35016
rect 1946 34200 59120 34480
rect 1946 33664 59200 34200
rect 1946 33384 59120 33664
rect 1946 32848 59200 33384
rect 1946 32568 59120 32848
rect 1946 32032 59200 32568
rect 1946 31752 59120 32032
rect 1946 31216 59200 31752
rect 1946 30936 59120 31216
rect 1946 30400 59200 30936
rect 1946 30120 59120 30400
rect 1946 29584 59200 30120
rect 1946 29304 59120 29584
rect 1946 28768 59200 29304
rect 1946 28488 59120 28768
rect 1946 27952 59200 28488
rect 1946 27672 59120 27952
rect 1946 27136 59200 27672
rect 1946 26856 59120 27136
rect 1946 26320 59200 26856
rect 1946 26040 59120 26320
rect 1946 25504 59200 26040
rect 1946 25224 59120 25504
rect 1946 24688 59200 25224
rect 1946 24408 59120 24688
rect 1946 23872 59200 24408
rect 1946 23592 59120 23872
rect 1946 23056 59200 23592
rect 1946 22776 59120 23056
rect 1946 22240 59200 22776
rect 1946 21960 59120 22240
rect 1946 21424 59200 21960
rect 1946 21144 59120 21424
rect 1946 20608 59200 21144
rect 1946 20328 59120 20608
rect 1946 19792 59200 20328
rect 1946 19512 59120 19792
rect 1946 18976 59200 19512
rect 1946 18696 59120 18976
rect 1946 18160 59200 18696
rect 1946 17880 59120 18160
rect 1946 17344 59200 17880
rect 1946 17064 59120 17344
rect 1946 16528 59200 17064
rect 1946 16248 59120 16528
rect 1946 15712 59200 16248
rect 1946 15432 59120 15712
rect 1946 14896 59200 15432
rect 1946 14616 59120 14896
rect 1946 14080 59200 14616
rect 1946 13800 59120 14080
rect 1946 13264 59200 13800
rect 1946 12984 59120 13264
rect 1946 12448 59200 12984
rect 1946 12168 59120 12448
rect 1946 11632 59200 12168
rect 1946 11352 59120 11632
rect 1946 10816 59200 11352
rect 1946 10536 59120 10816
rect 1946 10000 59200 10536
rect 1946 9720 59120 10000
rect 1946 9184 59200 9720
rect 1946 8904 59120 9184
rect 1946 8368 59200 8904
rect 1946 8088 59120 8368
rect 1946 7552 59200 8088
rect 1946 7272 59120 7552
rect 1946 6736 59200 7272
rect 1946 6456 59120 6736
rect 1946 5920 59200 6456
rect 1946 5640 59120 5920
rect 1946 5104 59200 5640
rect 1946 4824 59120 5104
rect 1946 4288 59200 4824
rect 1946 4008 59120 4288
rect 1946 2143 59200 4008
<< metal4 >>
rect 1944 2128 2264 57712
rect 2604 2128 2924 57712
rect 6944 2128 7264 57712
rect 7604 2128 7924 57712
rect 11944 2128 12264 57712
rect 12604 2128 12924 57712
rect 16944 2128 17264 57712
rect 17604 2128 17924 57712
rect 21944 2128 22264 57712
rect 22604 2128 22924 57712
rect 26944 2128 27264 57712
rect 27604 2128 27924 57712
rect 31944 2128 32264 57712
rect 32604 2128 32924 57712
rect 36944 2128 37264 57712
rect 37604 2128 37924 57712
rect 41944 2128 42264 57712
rect 42604 2128 42924 57712
rect 46944 2128 47264 57712
rect 47604 2128 47924 57712
rect 51944 2128 52264 57712
rect 52604 2128 52924 57712
rect 56944 2128 57264 57712
rect 57604 2128 57924 57712
<< metal5 >>
rect 1056 53676 58928 53996
rect 1056 53016 58928 53336
rect 1056 48676 58928 48996
rect 1056 48016 58928 48336
rect 1056 43676 58928 43996
rect 1056 43016 58928 43336
rect 1056 38676 58928 38996
rect 1056 38016 58928 38336
rect 1056 33676 58928 33996
rect 1056 33016 58928 33336
rect 1056 28676 58928 28996
rect 1056 28016 58928 28336
rect 1056 23676 58928 23996
rect 1056 23016 58928 23336
rect 1056 18676 58928 18996
rect 1056 18016 58928 18336
rect 1056 13676 58928 13996
rect 1056 13016 58928 13336
rect 1056 8676 58928 8996
rect 1056 8016 58928 8336
rect 1056 3676 58928 3996
rect 1056 3016 58928 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 22604 2128 22924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27604 2128 27924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 32604 2128 32924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37604 2128 37924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 42604 2128 42924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47604 2128 47924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 52604 2128 52924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 57604 2128 57924 57712 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 58928 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8676 58928 8996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13676 58928 13996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18676 58928 18996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 23676 58928 23996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 28676 58928 28996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 33676 58928 33996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 38676 58928 38996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 43676 58928 43996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 48676 58928 48996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 53676 58928 53996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 21944 2128 22264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26944 2128 27264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 31944 2128 32264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 36944 2128 37264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 41944 2128 42264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46944 2128 47264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 51944 2128 52264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 56944 2128 57264 57712 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 58928 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8016 58928 8336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13016 58928 13336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 18016 58928 18336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 23016 58928 23336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 28016 58928 28336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 33016 58928 33336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 38016 58928 38336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 43016 58928 43336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 48016 58928 48336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 53016 58928 53336 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 10072 800 10192 6 clk
port 3 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 control
port 4 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 reset
port 5 nsew signal input
rlabel metal3 s 59200 29384 60000 29504 6 result1[0]
port 6 nsew signal output
rlabel metal3 s 59200 21224 60000 21344 6 result1[10]
port 7 nsew signal output
rlabel metal3 s 59200 20408 60000 20528 6 result1[11]
port 8 nsew signal output
rlabel metal3 s 59200 19592 60000 19712 6 result1[12]
port 9 nsew signal output
rlabel metal3 s 59200 18776 60000 18896 6 result1[13]
port 10 nsew signal output
rlabel metal3 s 59200 17960 60000 18080 6 result1[14]
port 11 nsew signal output
rlabel metal3 s 59200 17144 60000 17264 6 result1[15]
port 12 nsew signal output
rlabel metal3 s 59200 16328 60000 16448 6 result1[16]
port 13 nsew signal output
rlabel metal3 s 59200 15512 60000 15632 6 result1[17]
port 14 nsew signal output
rlabel metal3 s 59200 14696 60000 14816 6 result1[18]
port 15 nsew signal output
rlabel metal3 s 59200 13880 60000 14000 6 result1[19]
port 16 nsew signal output
rlabel metal3 s 59200 28568 60000 28688 6 result1[1]
port 17 nsew signal output
rlabel metal3 s 59200 13064 60000 13184 6 result1[20]
port 18 nsew signal output
rlabel metal3 s 59200 12248 60000 12368 6 result1[21]
port 19 nsew signal output
rlabel metal3 s 59200 11432 60000 11552 6 result1[22]
port 20 nsew signal output
rlabel metal3 s 59200 10616 60000 10736 6 result1[23]
port 21 nsew signal output
rlabel metal3 s 59200 9800 60000 9920 6 result1[24]
port 22 nsew signal output
rlabel metal3 s 59200 8984 60000 9104 6 result1[25]
port 23 nsew signal output
rlabel metal3 s 59200 8168 60000 8288 6 result1[26]
port 24 nsew signal output
rlabel metal3 s 59200 7352 60000 7472 6 result1[27]
port 25 nsew signal output
rlabel metal3 s 59200 6536 60000 6656 6 result1[28]
port 26 nsew signal output
rlabel metal3 s 59200 5720 60000 5840 6 result1[29]
port 27 nsew signal output
rlabel metal3 s 59200 27752 60000 27872 6 result1[2]
port 28 nsew signal output
rlabel metal3 s 59200 4904 60000 5024 6 result1[30]
port 29 nsew signal output
rlabel metal3 s 59200 4088 60000 4208 6 result1[31]
port 30 nsew signal output
rlabel metal3 s 59200 26936 60000 27056 6 result1[3]
port 31 nsew signal output
rlabel metal3 s 59200 26120 60000 26240 6 result1[4]
port 32 nsew signal output
rlabel metal3 s 59200 25304 60000 25424 6 result1[5]
port 33 nsew signal output
rlabel metal3 s 59200 24488 60000 24608 6 result1[6]
port 34 nsew signal output
rlabel metal3 s 59200 23672 60000 23792 6 result1[7]
port 35 nsew signal output
rlabel metal3 s 59200 22856 60000 22976 6 result1[8]
port 36 nsew signal output
rlabel metal3 s 59200 22040 60000 22160 6 result1[9]
port 37 nsew signal output
rlabel metal3 s 59200 55496 60000 55616 6 result2[0]
port 38 nsew signal output
rlabel metal3 s 59200 47336 60000 47456 6 result2[10]
port 39 nsew signal output
rlabel metal3 s 59200 46520 60000 46640 6 result2[11]
port 40 nsew signal output
rlabel metal3 s 59200 45704 60000 45824 6 result2[12]
port 41 nsew signal output
rlabel metal3 s 59200 44888 60000 45008 6 result2[13]
port 42 nsew signal output
rlabel metal3 s 59200 44072 60000 44192 6 result2[14]
port 43 nsew signal output
rlabel metal3 s 59200 43256 60000 43376 6 result2[15]
port 44 nsew signal output
rlabel metal3 s 59200 42440 60000 42560 6 result2[16]
port 45 nsew signal output
rlabel metal3 s 59200 41624 60000 41744 6 result2[17]
port 46 nsew signal output
rlabel metal3 s 59200 40808 60000 40928 6 result2[18]
port 47 nsew signal output
rlabel metal3 s 59200 39992 60000 40112 6 result2[19]
port 48 nsew signal output
rlabel metal3 s 59200 54680 60000 54800 6 result2[1]
port 49 nsew signal output
rlabel metal3 s 59200 39176 60000 39296 6 result2[20]
port 50 nsew signal output
rlabel metal3 s 59200 38360 60000 38480 6 result2[21]
port 51 nsew signal output
rlabel metal3 s 59200 37544 60000 37664 6 result2[22]
port 52 nsew signal output
rlabel metal3 s 59200 36728 60000 36848 6 result2[23]
port 53 nsew signal output
rlabel metal3 s 59200 35912 60000 36032 6 result2[24]
port 54 nsew signal output
rlabel metal3 s 59200 35096 60000 35216 6 result2[25]
port 55 nsew signal output
rlabel metal3 s 59200 34280 60000 34400 6 result2[26]
port 56 nsew signal output
rlabel metal3 s 59200 33464 60000 33584 6 result2[27]
port 57 nsew signal output
rlabel metal3 s 59200 32648 60000 32768 6 result2[28]
port 58 nsew signal output
rlabel metal3 s 59200 31832 60000 31952 6 result2[29]
port 59 nsew signal output
rlabel metal3 s 59200 53864 60000 53984 6 result2[2]
port 60 nsew signal output
rlabel metal3 s 59200 31016 60000 31136 6 result2[30]
port 61 nsew signal output
rlabel metal3 s 59200 30200 60000 30320 6 result2[31]
port 62 nsew signal output
rlabel metal3 s 59200 53048 60000 53168 6 result2[3]
port 63 nsew signal output
rlabel metal3 s 59200 52232 60000 52352 6 result2[4]
port 64 nsew signal output
rlabel metal3 s 59200 51416 60000 51536 6 result2[5]
port 65 nsew signal output
rlabel metal3 s 59200 50600 60000 50720 6 result2[6]
port 66 nsew signal output
rlabel metal3 s 59200 49784 60000 49904 6 result2[7]
port 67 nsew signal output
rlabel metal3 s 59200 48968 60000 49088 6 result2[8]
port 68 nsew signal output
rlabel metal3 s 59200 48152 60000 48272 6 result2[9]
port 69 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1990308
string GDS_FILE /openlane/designs/project6/runs/RUN_2025.06.02_21.58.02/results/signoff/top_module.magic.gds
string GDS_START 22340
<< end >>

