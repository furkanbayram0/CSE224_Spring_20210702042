// This is the unpowered netlist.
module top_module (clk,
    control,
    reset,
    result1,
    result2);
 input clk;
 input control;
 input reset;
 output [31:0] result1;
 output [31:0] result2;

 wire net1;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net2;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net3;
 wire net31;
 wire net32;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net33;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net34;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net35;
 wire net63;
 wire net64;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_324 ();
 sky130_fd_sc_hd__conb_1 top_module_1 (.LO(net1));
 sky130_fd_sc_hd__conb_1 top_module_10 (.LO(net10));
 sky130_fd_sc_hd__conb_1 top_module_11 (.LO(net11));
 sky130_fd_sc_hd__conb_1 top_module_12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 top_module_13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 top_module_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 top_module_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 top_module_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 top_module_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 top_module_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 top_module_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 top_module_2 (.LO(net2));
 sky130_fd_sc_hd__conb_1 top_module_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 top_module_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 top_module_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 top_module_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 top_module_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 top_module_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 top_module_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 top_module_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 top_module_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 top_module_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 top_module_3 (.LO(net3));
 sky130_fd_sc_hd__conb_1 top_module_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 top_module_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 top_module_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 top_module_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 top_module_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 top_module_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 top_module_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 top_module_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 top_module_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 top_module_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 top_module_4 (.LO(net4));
 sky130_fd_sc_hd__conb_1 top_module_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 top_module_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 top_module_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 top_module_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 top_module_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 top_module_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 top_module_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 top_module_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 top_module_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 top_module_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 top_module_5 (.LO(net5));
 sky130_fd_sc_hd__conb_1 top_module_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 top_module_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 top_module_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 top_module_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 top_module_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 top_module_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 top_module_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 top_module_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 top_module_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 top_module_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 top_module_6 (.LO(net6));
 sky130_fd_sc_hd__conb_1 top_module_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 top_module_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 top_module_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 top_module_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 top_module_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 top_module_7 (.LO(net7));
 sky130_fd_sc_hd__conb_1 top_module_8 (.LO(net8));
 sky130_fd_sc_hd__conb_1 top_module_9 (.LO(net9));
 assign result1[0] = net1;
 assign result1[10] = net11;
 assign result1[11] = net12;
 assign result1[12] = net13;
 assign result1[13] = net14;
 assign result1[14] = net15;
 assign result1[15] = net16;
 assign result1[16] = net17;
 assign result1[17] = net18;
 assign result1[18] = net19;
 assign result1[19] = net20;
 assign result1[1] = net2;
 assign result1[20] = net21;
 assign result1[21] = net22;
 assign result1[22] = net23;
 assign result1[23] = net24;
 assign result1[24] = net25;
 assign result1[25] = net26;
 assign result1[26] = net27;
 assign result1[27] = net28;
 assign result1[28] = net29;
 assign result1[29] = net30;
 assign result1[2] = net3;
 assign result1[30] = net31;
 assign result1[31] = net32;
 assign result1[3] = net4;
 assign result1[4] = net5;
 assign result1[5] = net6;
 assign result1[6] = net7;
 assign result1[7] = net8;
 assign result1[8] = net9;
 assign result1[9] = net10;
 assign result2[0] = net33;
 assign result2[10] = net43;
 assign result2[11] = net44;
 assign result2[12] = net45;
 assign result2[13] = net46;
 assign result2[14] = net47;
 assign result2[15] = net48;
 assign result2[16] = net49;
 assign result2[17] = net50;
 assign result2[18] = net51;
 assign result2[19] = net52;
 assign result2[1] = net34;
 assign result2[20] = net53;
 assign result2[21] = net54;
 assign result2[22] = net55;
 assign result2[23] = net56;
 assign result2[24] = net57;
 assign result2[25] = net58;
 assign result2[26] = net59;
 assign result2[27] = net60;
 assign result2[28] = net61;
 assign result2[29] = net62;
 assign result2[2] = net35;
 assign result2[30] = net63;
 assign result2[31] = net64;
 assign result2[3] = net36;
 assign result2[4] = net37;
 assign result2[5] = net38;
 assign result2[6] = net39;
 assign result2[7] = net40;
 assign result2[8] = net41;
 assign result2[9] = net42;
endmodule

