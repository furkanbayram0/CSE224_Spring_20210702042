magic
tech sky130A
magscale 1 2
timestamp 1747871249
<< nwell >>
rect 1066 2159 14850 15814
<< obsli1 >>
rect 1104 2159 14812 15793
<< obsm1 >>
rect 658 1640 15718 15972
<< obsm2 >>
rect 664 1119 15712 16425
<< metal3 >>
rect 15200 16328 16000 16448
rect 15200 15240 16000 15360
rect 15200 14152 16000 14272
rect 0 13336 800 13456
rect 15200 13064 16000 13184
rect 15200 11976 16000 12096
rect 15200 10888 16000 11008
rect 15200 9800 16000 9920
rect 15200 8712 16000 8832
rect 15200 7624 16000 7744
rect 15200 6536 16000 6656
rect 15200 5448 16000 5568
rect 0 4360 800 4480
rect 15200 4360 16000 4480
rect 15200 3272 16000 3392
rect 15200 2184 16000 2304
rect 15200 1096 16000 1216
<< obsm3 >>
rect 606 16248 15120 16421
rect 606 15440 15200 16248
rect 606 15160 15120 15440
rect 606 14352 15200 15160
rect 606 14072 15120 14352
rect 606 13536 15200 14072
rect 880 13264 15200 13536
rect 880 13256 15120 13264
rect 606 12984 15120 13256
rect 606 12176 15200 12984
rect 606 11896 15120 12176
rect 606 11088 15200 11896
rect 606 10808 15120 11088
rect 606 10000 15200 10808
rect 606 9720 15120 10000
rect 606 8912 15200 9720
rect 606 8632 15120 8912
rect 606 7824 15200 8632
rect 606 7544 15120 7824
rect 606 6736 15200 7544
rect 606 6456 15120 6736
rect 606 5648 15200 6456
rect 606 5368 15120 5648
rect 606 4560 15200 5368
rect 880 4280 15120 4560
rect 606 3472 15200 4280
rect 606 3192 15120 3472
rect 606 2384 15200 3192
rect 606 2104 15120 2384
rect 606 1296 15200 2104
rect 606 1123 15120 1296
<< metal4 >>
rect 1944 2128 2264 15824
rect 2604 2128 2924 15824
rect 6944 2128 7264 15824
rect 7604 2128 7924 15824
rect 11944 2128 12264 15824
rect 12604 2128 12924 15824
<< obsm4 >>
rect 611 2048 1864 15469
rect 2344 2048 2524 15469
rect 3004 2048 6864 15469
rect 7344 2048 7524 15469
rect 8004 2048 11864 15469
rect 12344 2048 12524 15469
rect 13004 2048 14109 15469
rect 611 1531 14109 2048
<< metal5 >>
rect 1056 13676 14860 13996
rect 1056 13016 14860 13336
rect 1056 8676 14860 8996
rect 1056 8016 14860 8336
rect 1056 3676 14860 3996
rect 1056 3016 14860 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 15824 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 15824 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 15824 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 14860 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8676 14860 8996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13676 14860 13996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 15824 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 15824 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 15824 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 14860 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8016 14860 8336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13016 14860 13336 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 15200 8712 16000 8832 6 an0
port 3 nsew signal output
rlabel metal3 s 15200 9800 16000 9920 6 an1
port 4 nsew signal output
rlabel metal3 s 15200 10888 16000 11008 6 an2
port 5 nsew signal output
rlabel metal3 s 15200 11976 16000 12096 6 an3
port 6 nsew signal output
rlabel metal3 s 15200 13064 16000 13184 6 an4
port 7 nsew signal output
rlabel metal3 s 15200 14152 16000 14272 6 an5
port 8 nsew signal output
rlabel metal3 s 15200 15240 16000 15360 6 an6
port 9 nsew signal output
rlabel metal3 s 15200 16328 16000 16448 6 an7
port 10 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 clk
port 11 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 rst
port 12 nsew signal input
rlabel metal3 s 15200 1096 16000 1216 6 seg0
port 13 nsew signal output
rlabel metal3 s 15200 2184 16000 2304 6 seg1
port 14 nsew signal output
rlabel metal3 s 15200 3272 16000 3392 6 seg2
port 15 nsew signal output
rlabel metal3 s 15200 4360 16000 4480 6 seg3
port 16 nsew signal output
rlabel metal3 s 15200 5448 16000 5568 6 seg4
port 17 nsew signal output
rlabel metal3 s 15200 6536 16000 6656 6 seg5
port 18 nsew signal output
rlabel metal3 s 15200 7624 16000 7744 6 seg6
port 19 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 16000 18000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1230036
string GDS_FILE /openlane/designs/project3/runs/RUN_2025.05.21_23.45.57/results/signoff/project3.magic.gds
string GDS_START 315288
<< end >>

