magic
tech sky130A
magscale 1 2
timestamp 1748901528
<< checkpaint >>
rect -3932 -1804 63932 61644
<< viali >>
rect 58541 55709 58575 55743
rect 58541 55029 58575 55063
rect 58541 53941 58575 53975
rect 58541 53533 58575 53567
rect 58541 52445 58575 52479
rect 58541 51765 58575 51799
rect 58541 50677 58575 50711
rect 58541 50269 58575 50303
rect 58541 49181 58575 49215
rect 58541 48501 58575 48535
rect 58541 47413 58575 47447
rect 58541 47005 58575 47039
rect 58541 45917 58575 45951
rect 58541 45237 58575 45271
rect 58541 44149 58575 44183
rect 58541 43741 58575 43775
rect 58541 42653 58575 42687
rect 58541 41973 58575 42007
rect 58541 40885 58575 40919
rect 58541 40477 58575 40511
rect 58541 39389 58575 39423
rect 58541 38709 58575 38743
rect 58541 37621 58575 37655
rect 58541 37281 58575 37315
rect 58541 36125 58575 36159
rect 58541 35445 58575 35479
rect 58541 34357 58575 34391
rect 58541 33949 58575 33983
rect 58541 32861 58575 32895
rect 58541 32181 58575 32215
rect 58541 31093 58575 31127
rect 58541 30685 58575 30719
rect 58541 29597 58575 29631
rect 58541 28985 58575 29019
rect 58541 27829 58575 27863
rect 58541 27421 58575 27455
rect 58541 26333 58575 26367
rect 58541 25653 58575 25687
rect 58541 24565 58575 24599
rect 58541 24157 58575 24191
rect 58541 23069 58575 23103
rect 58541 22389 58575 22423
rect 58541 21301 58575 21335
rect 58541 20893 58575 20927
rect 58541 19805 58575 19839
rect 58541 19125 58575 19159
rect 58541 18037 58575 18071
rect 58541 17629 58575 17663
rect 58541 16609 58575 16643
rect 58541 15861 58575 15895
rect 58541 14773 58575 14807
rect 58541 14365 58575 14399
rect 58541 13277 58575 13311
rect 58541 12597 58575 12631
rect 58541 11509 58575 11543
rect 58541 11101 58575 11135
rect 58541 10013 58575 10047
rect 58541 9333 58575 9367
rect 58541 8313 58575 8347
rect 58541 7837 58575 7871
rect 58541 6749 58575 6783
rect 58541 6069 58575 6103
rect 58541 4981 58575 5015
rect 58541 4573 58575 4607
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 2610 57690
rect 2662 57638 2674 57690
rect 2726 57638 2738 57690
rect 2790 57638 2802 57690
rect 2854 57638 2866 57690
rect 2918 57638 7610 57690
rect 7662 57638 7674 57690
rect 7726 57638 7738 57690
rect 7790 57638 7802 57690
rect 7854 57638 7866 57690
rect 7918 57638 12610 57690
rect 12662 57638 12674 57690
rect 12726 57638 12738 57690
rect 12790 57638 12802 57690
rect 12854 57638 12866 57690
rect 12918 57638 17610 57690
rect 17662 57638 17674 57690
rect 17726 57638 17738 57690
rect 17790 57638 17802 57690
rect 17854 57638 17866 57690
rect 17918 57638 22610 57690
rect 22662 57638 22674 57690
rect 22726 57638 22738 57690
rect 22790 57638 22802 57690
rect 22854 57638 22866 57690
rect 22918 57638 27610 57690
rect 27662 57638 27674 57690
rect 27726 57638 27738 57690
rect 27790 57638 27802 57690
rect 27854 57638 27866 57690
rect 27918 57638 32610 57690
rect 32662 57638 32674 57690
rect 32726 57638 32738 57690
rect 32790 57638 32802 57690
rect 32854 57638 32866 57690
rect 32918 57638 37610 57690
rect 37662 57638 37674 57690
rect 37726 57638 37738 57690
rect 37790 57638 37802 57690
rect 37854 57638 37866 57690
rect 37918 57638 42610 57690
rect 42662 57638 42674 57690
rect 42726 57638 42738 57690
rect 42790 57638 42802 57690
rect 42854 57638 42866 57690
rect 42918 57638 47610 57690
rect 47662 57638 47674 57690
rect 47726 57638 47738 57690
rect 47790 57638 47802 57690
rect 47854 57638 47866 57690
rect 47918 57638 52610 57690
rect 52662 57638 52674 57690
rect 52726 57638 52738 57690
rect 52790 57638 52802 57690
rect 52854 57638 52866 57690
rect 52918 57638 57610 57690
rect 57662 57638 57674 57690
rect 57726 57638 57738 57690
rect 57790 57638 57802 57690
rect 57854 57638 57866 57690
rect 57918 57638 58880 57690
rect 1104 57616 58880 57638
rect 1104 57146 58880 57168
rect 1104 57094 1950 57146
rect 2002 57094 2014 57146
rect 2066 57094 2078 57146
rect 2130 57094 2142 57146
rect 2194 57094 2206 57146
rect 2258 57094 6950 57146
rect 7002 57094 7014 57146
rect 7066 57094 7078 57146
rect 7130 57094 7142 57146
rect 7194 57094 7206 57146
rect 7258 57094 11950 57146
rect 12002 57094 12014 57146
rect 12066 57094 12078 57146
rect 12130 57094 12142 57146
rect 12194 57094 12206 57146
rect 12258 57094 16950 57146
rect 17002 57094 17014 57146
rect 17066 57094 17078 57146
rect 17130 57094 17142 57146
rect 17194 57094 17206 57146
rect 17258 57094 21950 57146
rect 22002 57094 22014 57146
rect 22066 57094 22078 57146
rect 22130 57094 22142 57146
rect 22194 57094 22206 57146
rect 22258 57094 26950 57146
rect 27002 57094 27014 57146
rect 27066 57094 27078 57146
rect 27130 57094 27142 57146
rect 27194 57094 27206 57146
rect 27258 57094 31950 57146
rect 32002 57094 32014 57146
rect 32066 57094 32078 57146
rect 32130 57094 32142 57146
rect 32194 57094 32206 57146
rect 32258 57094 36950 57146
rect 37002 57094 37014 57146
rect 37066 57094 37078 57146
rect 37130 57094 37142 57146
rect 37194 57094 37206 57146
rect 37258 57094 41950 57146
rect 42002 57094 42014 57146
rect 42066 57094 42078 57146
rect 42130 57094 42142 57146
rect 42194 57094 42206 57146
rect 42258 57094 46950 57146
rect 47002 57094 47014 57146
rect 47066 57094 47078 57146
rect 47130 57094 47142 57146
rect 47194 57094 47206 57146
rect 47258 57094 51950 57146
rect 52002 57094 52014 57146
rect 52066 57094 52078 57146
rect 52130 57094 52142 57146
rect 52194 57094 52206 57146
rect 52258 57094 56950 57146
rect 57002 57094 57014 57146
rect 57066 57094 57078 57146
rect 57130 57094 57142 57146
rect 57194 57094 57206 57146
rect 57258 57094 58880 57146
rect 1104 57072 58880 57094
rect 1104 56602 58880 56624
rect 1104 56550 2610 56602
rect 2662 56550 2674 56602
rect 2726 56550 2738 56602
rect 2790 56550 2802 56602
rect 2854 56550 2866 56602
rect 2918 56550 7610 56602
rect 7662 56550 7674 56602
rect 7726 56550 7738 56602
rect 7790 56550 7802 56602
rect 7854 56550 7866 56602
rect 7918 56550 12610 56602
rect 12662 56550 12674 56602
rect 12726 56550 12738 56602
rect 12790 56550 12802 56602
rect 12854 56550 12866 56602
rect 12918 56550 17610 56602
rect 17662 56550 17674 56602
rect 17726 56550 17738 56602
rect 17790 56550 17802 56602
rect 17854 56550 17866 56602
rect 17918 56550 22610 56602
rect 22662 56550 22674 56602
rect 22726 56550 22738 56602
rect 22790 56550 22802 56602
rect 22854 56550 22866 56602
rect 22918 56550 27610 56602
rect 27662 56550 27674 56602
rect 27726 56550 27738 56602
rect 27790 56550 27802 56602
rect 27854 56550 27866 56602
rect 27918 56550 32610 56602
rect 32662 56550 32674 56602
rect 32726 56550 32738 56602
rect 32790 56550 32802 56602
rect 32854 56550 32866 56602
rect 32918 56550 37610 56602
rect 37662 56550 37674 56602
rect 37726 56550 37738 56602
rect 37790 56550 37802 56602
rect 37854 56550 37866 56602
rect 37918 56550 42610 56602
rect 42662 56550 42674 56602
rect 42726 56550 42738 56602
rect 42790 56550 42802 56602
rect 42854 56550 42866 56602
rect 42918 56550 47610 56602
rect 47662 56550 47674 56602
rect 47726 56550 47738 56602
rect 47790 56550 47802 56602
rect 47854 56550 47866 56602
rect 47918 56550 52610 56602
rect 52662 56550 52674 56602
rect 52726 56550 52738 56602
rect 52790 56550 52802 56602
rect 52854 56550 52866 56602
rect 52918 56550 57610 56602
rect 57662 56550 57674 56602
rect 57726 56550 57738 56602
rect 57790 56550 57802 56602
rect 57854 56550 57866 56602
rect 57918 56550 58880 56602
rect 1104 56528 58880 56550
rect 1104 56058 58880 56080
rect 1104 56006 1950 56058
rect 2002 56006 2014 56058
rect 2066 56006 2078 56058
rect 2130 56006 2142 56058
rect 2194 56006 2206 56058
rect 2258 56006 6950 56058
rect 7002 56006 7014 56058
rect 7066 56006 7078 56058
rect 7130 56006 7142 56058
rect 7194 56006 7206 56058
rect 7258 56006 11950 56058
rect 12002 56006 12014 56058
rect 12066 56006 12078 56058
rect 12130 56006 12142 56058
rect 12194 56006 12206 56058
rect 12258 56006 16950 56058
rect 17002 56006 17014 56058
rect 17066 56006 17078 56058
rect 17130 56006 17142 56058
rect 17194 56006 17206 56058
rect 17258 56006 21950 56058
rect 22002 56006 22014 56058
rect 22066 56006 22078 56058
rect 22130 56006 22142 56058
rect 22194 56006 22206 56058
rect 22258 56006 26950 56058
rect 27002 56006 27014 56058
rect 27066 56006 27078 56058
rect 27130 56006 27142 56058
rect 27194 56006 27206 56058
rect 27258 56006 31950 56058
rect 32002 56006 32014 56058
rect 32066 56006 32078 56058
rect 32130 56006 32142 56058
rect 32194 56006 32206 56058
rect 32258 56006 36950 56058
rect 37002 56006 37014 56058
rect 37066 56006 37078 56058
rect 37130 56006 37142 56058
rect 37194 56006 37206 56058
rect 37258 56006 41950 56058
rect 42002 56006 42014 56058
rect 42066 56006 42078 56058
rect 42130 56006 42142 56058
rect 42194 56006 42206 56058
rect 42258 56006 46950 56058
rect 47002 56006 47014 56058
rect 47066 56006 47078 56058
rect 47130 56006 47142 56058
rect 47194 56006 47206 56058
rect 47258 56006 51950 56058
rect 52002 56006 52014 56058
rect 52066 56006 52078 56058
rect 52130 56006 52142 56058
rect 52194 56006 52206 56058
rect 52258 56006 56950 56058
rect 57002 56006 57014 56058
rect 57066 56006 57078 56058
rect 57130 56006 57142 56058
rect 57194 56006 57206 56058
rect 57258 56006 58880 56058
rect 1104 55984 58880 56006
rect 58526 55700 58532 55752
rect 58584 55700 58590 55752
rect 1104 55514 58880 55536
rect 1104 55462 2610 55514
rect 2662 55462 2674 55514
rect 2726 55462 2738 55514
rect 2790 55462 2802 55514
rect 2854 55462 2866 55514
rect 2918 55462 7610 55514
rect 7662 55462 7674 55514
rect 7726 55462 7738 55514
rect 7790 55462 7802 55514
rect 7854 55462 7866 55514
rect 7918 55462 12610 55514
rect 12662 55462 12674 55514
rect 12726 55462 12738 55514
rect 12790 55462 12802 55514
rect 12854 55462 12866 55514
rect 12918 55462 17610 55514
rect 17662 55462 17674 55514
rect 17726 55462 17738 55514
rect 17790 55462 17802 55514
rect 17854 55462 17866 55514
rect 17918 55462 22610 55514
rect 22662 55462 22674 55514
rect 22726 55462 22738 55514
rect 22790 55462 22802 55514
rect 22854 55462 22866 55514
rect 22918 55462 27610 55514
rect 27662 55462 27674 55514
rect 27726 55462 27738 55514
rect 27790 55462 27802 55514
rect 27854 55462 27866 55514
rect 27918 55462 32610 55514
rect 32662 55462 32674 55514
rect 32726 55462 32738 55514
rect 32790 55462 32802 55514
rect 32854 55462 32866 55514
rect 32918 55462 37610 55514
rect 37662 55462 37674 55514
rect 37726 55462 37738 55514
rect 37790 55462 37802 55514
rect 37854 55462 37866 55514
rect 37918 55462 42610 55514
rect 42662 55462 42674 55514
rect 42726 55462 42738 55514
rect 42790 55462 42802 55514
rect 42854 55462 42866 55514
rect 42918 55462 47610 55514
rect 47662 55462 47674 55514
rect 47726 55462 47738 55514
rect 47790 55462 47802 55514
rect 47854 55462 47866 55514
rect 47918 55462 52610 55514
rect 52662 55462 52674 55514
rect 52726 55462 52738 55514
rect 52790 55462 52802 55514
rect 52854 55462 52866 55514
rect 52918 55462 57610 55514
rect 57662 55462 57674 55514
rect 57726 55462 57738 55514
rect 57790 55462 57802 55514
rect 57854 55462 57866 55514
rect 57918 55462 58880 55514
rect 1104 55440 58880 55462
rect 58526 55020 58532 55072
rect 58584 55020 58590 55072
rect 1104 54970 58880 54992
rect 1104 54918 1950 54970
rect 2002 54918 2014 54970
rect 2066 54918 2078 54970
rect 2130 54918 2142 54970
rect 2194 54918 2206 54970
rect 2258 54918 6950 54970
rect 7002 54918 7014 54970
rect 7066 54918 7078 54970
rect 7130 54918 7142 54970
rect 7194 54918 7206 54970
rect 7258 54918 11950 54970
rect 12002 54918 12014 54970
rect 12066 54918 12078 54970
rect 12130 54918 12142 54970
rect 12194 54918 12206 54970
rect 12258 54918 16950 54970
rect 17002 54918 17014 54970
rect 17066 54918 17078 54970
rect 17130 54918 17142 54970
rect 17194 54918 17206 54970
rect 17258 54918 21950 54970
rect 22002 54918 22014 54970
rect 22066 54918 22078 54970
rect 22130 54918 22142 54970
rect 22194 54918 22206 54970
rect 22258 54918 26950 54970
rect 27002 54918 27014 54970
rect 27066 54918 27078 54970
rect 27130 54918 27142 54970
rect 27194 54918 27206 54970
rect 27258 54918 31950 54970
rect 32002 54918 32014 54970
rect 32066 54918 32078 54970
rect 32130 54918 32142 54970
rect 32194 54918 32206 54970
rect 32258 54918 36950 54970
rect 37002 54918 37014 54970
rect 37066 54918 37078 54970
rect 37130 54918 37142 54970
rect 37194 54918 37206 54970
rect 37258 54918 41950 54970
rect 42002 54918 42014 54970
rect 42066 54918 42078 54970
rect 42130 54918 42142 54970
rect 42194 54918 42206 54970
rect 42258 54918 46950 54970
rect 47002 54918 47014 54970
rect 47066 54918 47078 54970
rect 47130 54918 47142 54970
rect 47194 54918 47206 54970
rect 47258 54918 51950 54970
rect 52002 54918 52014 54970
rect 52066 54918 52078 54970
rect 52130 54918 52142 54970
rect 52194 54918 52206 54970
rect 52258 54918 56950 54970
rect 57002 54918 57014 54970
rect 57066 54918 57078 54970
rect 57130 54918 57142 54970
rect 57194 54918 57206 54970
rect 57258 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 2610 54426
rect 2662 54374 2674 54426
rect 2726 54374 2738 54426
rect 2790 54374 2802 54426
rect 2854 54374 2866 54426
rect 2918 54374 7610 54426
rect 7662 54374 7674 54426
rect 7726 54374 7738 54426
rect 7790 54374 7802 54426
rect 7854 54374 7866 54426
rect 7918 54374 12610 54426
rect 12662 54374 12674 54426
rect 12726 54374 12738 54426
rect 12790 54374 12802 54426
rect 12854 54374 12866 54426
rect 12918 54374 17610 54426
rect 17662 54374 17674 54426
rect 17726 54374 17738 54426
rect 17790 54374 17802 54426
rect 17854 54374 17866 54426
rect 17918 54374 22610 54426
rect 22662 54374 22674 54426
rect 22726 54374 22738 54426
rect 22790 54374 22802 54426
rect 22854 54374 22866 54426
rect 22918 54374 27610 54426
rect 27662 54374 27674 54426
rect 27726 54374 27738 54426
rect 27790 54374 27802 54426
rect 27854 54374 27866 54426
rect 27918 54374 32610 54426
rect 32662 54374 32674 54426
rect 32726 54374 32738 54426
rect 32790 54374 32802 54426
rect 32854 54374 32866 54426
rect 32918 54374 37610 54426
rect 37662 54374 37674 54426
rect 37726 54374 37738 54426
rect 37790 54374 37802 54426
rect 37854 54374 37866 54426
rect 37918 54374 42610 54426
rect 42662 54374 42674 54426
rect 42726 54374 42738 54426
rect 42790 54374 42802 54426
rect 42854 54374 42866 54426
rect 42918 54374 47610 54426
rect 47662 54374 47674 54426
rect 47726 54374 47738 54426
rect 47790 54374 47802 54426
rect 47854 54374 47866 54426
rect 47918 54374 52610 54426
rect 52662 54374 52674 54426
rect 52726 54374 52738 54426
rect 52790 54374 52802 54426
rect 52854 54374 52866 54426
rect 52918 54374 57610 54426
rect 57662 54374 57674 54426
rect 57726 54374 57738 54426
rect 57790 54374 57802 54426
rect 57854 54374 57866 54426
rect 57918 54374 58880 54426
rect 1104 54352 58880 54374
rect 58526 53932 58532 53984
rect 58584 53932 58590 53984
rect 1104 53882 58880 53904
rect 1104 53830 1950 53882
rect 2002 53830 2014 53882
rect 2066 53830 2078 53882
rect 2130 53830 2142 53882
rect 2194 53830 2206 53882
rect 2258 53830 6950 53882
rect 7002 53830 7014 53882
rect 7066 53830 7078 53882
rect 7130 53830 7142 53882
rect 7194 53830 7206 53882
rect 7258 53830 11950 53882
rect 12002 53830 12014 53882
rect 12066 53830 12078 53882
rect 12130 53830 12142 53882
rect 12194 53830 12206 53882
rect 12258 53830 16950 53882
rect 17002 53830 17014 53882
rect 17066 53830 17078 53882
rect 17130 53830 17142 53882
rect 17194 53830 17206 53882
rect 17258 53830 21950 53882
rect 22002 53830 22014 53882
rect 22066 53830 22078 53882
rect 22130 53830 22142 53882
rect 22194 53830 22206 53882
rect 22258 53830 26950 53882
rect 27002 53830 27014 53882
rect 27066 53830 27078 53882
rect 27130 53830 27142 53882
rect 27194 53830 27206 53882
rect 27258 53830 31950 53882
rect 32002 53830 32014 53882
rect 32066 53830 32078 53882
rect 32130 53830 32142 53882
rect 32194 53830 32206 53882
rect 32258 53830 36950 53882
rect 37002 53830 37014 53882
rect 37066 53830 37078 53882
rect 37130 53830 37142 53882
rect 37194 53830 37206 53882
rect 37258 53830 41950 53882
rect 42002 53830 42014 53882
rect 42066 53830 42078 53882
rect 42130 53830 42142 53882
rect 42194 53830 42206 53882
rect 42258 53830 46950 53882
rect 47002 53830 47014 53882
rect 47066 53830 47078 53882
rect 47130 53830 47142 53882
rect 47194 53830 47206 53882
rect 47258 53830 51950 53882
rect 52002 53830 52014 53882
rect 52066 53830 52078 53882
rect 52130 53830 52142 53882
rect 52194 53830 52206 53882
rect 52258 53830 56950 53882
rect 57002 53830 57014 53882
rect 57066 53830 57078 53882
rect 57130 53830 57142 53882
rect 57194 53830 57206 53882
rect 57258 53830 58880 53882
rect 1104 53808 58880 53830
rect 58526 53524 58532 53576
rect 58584 53524 58590 53576
rect 1104 53338 58880 53360
rect 1104 53286 2610 53338
rect 2662 53286 2674 53338
rect 2726 53286 2738 53338
rect 2790 53286 2802 53338
rect 2854 53286 2866 53338
rect 2918 53286 7610 53338
rect 7662 53286 7674 53338
rect 7726 53286 7738 53338
rect 7790 53286 7802 53338
rect 7854 53286 7866 53338
rect 7918 53286 12610 53338
rect 12662 53286 12674 53338
rect 12726 53286 12738 53338
rect 12790 53286 12802 53338
rect 12854 53286 12866 53338
rect 12918 53286 17610 53338
rect 17662 53286 17674 53338
rect 17726 53286 17738 53338
rect 17790 53286 17802 53338
rect 17854 53286 17866 53338
rect 17918 53286 22610 53338
rect 22662 53286 22674 53338
rect 22726 53286 22738 53338
rect 22790 53286 22802 53338
rect 22854 53286 22866 53338
rect 22918 53286 27610 53338
rect 27662 53286 27674 53338
rect 27726 53286 27738 53338
rect 27790 53286 27802 53338
rect 27854 53286 27866 53338
rect 27918 53286 32610 53338
rect 32662 53286 32674 53338
rect 32726 53286 32738 53338
rect 32790 53286 32802 53338
rect 32854 53286 32866 53338
rect 32918 53286 37610 53338
rect 37662 53286 37674 53338
rect 37726 53286 37738 53338
rect 37790 53286 37802 53338
rect 37854 53286 37866 53338
rect 37918 53286 42610 53338
rect 42662 53286 42674 53338
rect 42726 53286 42738 53338
rect 42790 53286 42802 53338
rect 42854 53286 42866 53338
rect 42918 53286 47610 53338
rect 47662 53286 47674 53338
rect 47726 53286 47738 53338
rect 47790 53286 47802 53338
rect 47854 53286 47866 53338
rect 47918 53286 52610 53338
rect 52662 53286 52674 53338
rect 52726 53286 52738 53338
rect 52790 53286 52802 53338
rect 52854 53286 52866 53338
rect 52918 53286 57610 53338
rect 57662 53286 57674 53338
rect 57726 53286 57738 53338
rect 57790 53286 57802 53338
rect 57854 53286 57866 53338
rect 57918 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 1950 52794
rect 2002 52742 2014 52794
rect 2066 52742 2078 52794
rect 2130 52742 2142 52794
rect 2194 52742 2206 52794
rect 2258 52742 6950 52794
rect 7002 52742 7014 52794
rect 7066 52742 7078 52794
rect 7130 52742 7142 52794
rect 7194 52742 7206 52794
rect 7258 52742 11950 52794
rect 12002 52742 12014 52794
rect 12066 52742 12078 52794
rect 12130 52742 12142 52794
rect 12194 52742 12206 52794
rect 12258 52742 16950 52794
rect 17002 52742 17014 52794
rect 17066 52742 17078 52794
rect 17130 52742 17142 52794
rect 17194 52742 17206 52794
rect 17258 52742 21950 52794
rect 22002 52742 22014 52794
rect 22066 52742 22078 52794
rect 22130 52742 22142 52794
rect 22194 52742 22206 52794
rect 22258 52742 26950 52794
rect 27002 52742 27014 52794
rect 27066 52742 27078 52794
rect 27130 52742 27142 52794
rect 27194 52742 27206 52794
rect 27258 52742 31950 52794
rect 32002 52742 32014 52794
rect 32066 52742 32078 52794
rect 32130 52742 32142 52794
rect 32194 52742 32206 52794
rect 32258 52742 36950 52794
rect 37002 52742 37014 52794
rect 37066 52742 37078 52794
rect 37130 52742 37142 52794
rect 37194 52742 37206 52794
rect 37258 52742 41950 52794
rect 42002 52742 42014 52794
rect 42066 52742 42078 52794
rect 42130 52742 42142 52794
rect 42194 52742 42206 52794
rect 42258 52742 46950 52794
rect 47002 52742 47014 52794
rect 47066 52742 47078 52794
rect 47130 52742 47142 52794
rect 47194 52742 47206 52794
rect 47258 52742 51950 52794
rect 52002 52742 52014 52794
rect 52066 52742 52078 52794
rect 52130 52742 52142 52794
rect 52194 52742 52206 52794
rect 52258 52742 56950 52794
rect 57002 52742 57014 52794
rect 57066 52742 57078 52794
rect 57130 52742 57142 52794
rect 57194 52742 57206 52794
rect 57258 52742 58880 52794
rect 1104 52720 58880 52742
rect 58526 52436 58532 52488
rect 58584 52436 58590 52488
rect 1104 52250 58880 52272
rect 1104 52198 2610 52250
rect 2662 52198 2674 52250
rect 2726 52198 2738 52250
rect 2790 52198 2802 52250
rect 2854 52198 2866 52250
rect 2918 52198 7610 52250
rect 7662 52198 7674 52250
rect 7726 52198 7738 52250
rect 7790 52198 7802 52250
rect 7854 52198 7866 52250
rect 7918 52198 12610 52250
rect 12662 52198 12674 52250
rect 12726 52198 12738 52250
rect 12790 52198 12802 52250
rect 12854 52198 12866 52250
rect 12918 52198 17610 52250
rect 17662 52198 17674 52250
rect 17726 52198 17738 52250
rect 17790 52198 17802 52250
rect 17854 52198 17866 52250
rect 17918 52198 22610 52250
rect 22662 52198 22674 52250
rect 22726 52198 22738 52250
rect 22790 52198 22802 52250
rect 22854 52198 22866 52250
rect 22918 52198 27610 52250
rect 27662 52198 27674 52250
rect 27726 52198 27738 52250
rect 27790 52198 27802 52250
rect 27854 52198 27866 52250
rect 27918 52198 32610 52250
rect 32662 52198 32674 52250
rect 32726 52198 32738 52250
rect 32790 52198 32802 52250
rect 32854 52198 32866 52250
rect 32918 52198 37610 52250
rect 37662 52198 37674 52250
rect 37726 52198 37738 52250
rect 37790 52198 37802 52250
rect 37854 52198 37866 52250
rect 37918 52198 42610 52250
rect 42662 52198 42674 52250
rect 42726 52198 42738 52250
rect 42790 52198 42802 52250
rect 42854 52198 42866 52250
rect 42918 52198 47610 52250
rect 47662 52198 47674 52250
rect 47726 52198 47738 52250
rect 47790 52198 47802 52250
rect 47854 52198 47866 52250
rect 47918 52198 52610 52250
rect 52662 52198 52674 52250
rect 52726 52198 52738 52250
rect 52790 52198 52802 52250
rect 52854 52198 52866 52250
rect 52918 52198 57610 52250
rect 57662 52198 57674 52250
rect 57726 52198 57738 52250
rect 57790 52198 57802 52250
rect 57854 52198 57866 52250
rect 57918 52198 58880 52250
rect 1104 52176 58880 52198
rect 58526 51756 58532 51808
rect 58584 51756 58590 51808
rect 1104 51706 58880 51728
rect 1104 51654 1950 51706
rect 2002 51654 2014 51706
rect 2066 51654 2078 51706
rect 2130 51654 2142 51706
rect 2194 51654 2206 51706
rect 2258 51654 6950 51706
rect 7002 51654 7014 51706
rect 7066 51654 7078 51706
rect 7130 51654 7142 51706
rect 7194 51654 7206 51706
rect 7258 51654 11950 51706
rect 12002 51654 12014 51706
rect 12066 51654 12078 51706
rect 12130 51654 12142 51706
rect 12194 51654 12206 51706
rect 12258 51654 16950 51706
rect 17002 51654 17014 51706
rect 17066 51654 17078 51706
rect 17130 51654 17142 51706
rect 17194 51654 17206 51706
rect 17258 51654 21950 51706
rect 22002 51654 22014 51706
rect 22066 51654 22078 51706
rect 22130 51654 22142 51706
rect 22194 51654 22206 51706
rect 22258 51654 26950 51706
rect 27002 51654 27014 51706
rect 27066 51654 27078 51706
rect 27130 51654 27142 51706
rect 27194 51654 27206 51706
rect 27258 51654 31950 51706
rect 32002 51654 32014 51706
rect 32066 51654 32078 51706
rect 32130 51654 32142 51706
rect 32194 51654 32206 51706
rect 32258 51654 36950 51706
rect 37002 51654 37014 51706
rect 37066 51654 37078 51706
rect 37130 51654 37142 51706
rect 37194 51654 37206 51706
rect 37258 51654 41950 51706
rect 42002 51654 42014 51706
rect 42066 51654 42078 51706
rect 42130 51654 42142 51706
rect 42194 51654 42206 51706
rect 42258 51654 46950 51706
rect 47002 51654 47014 51706
rect 47066 51654 47078 51706
rect 47130 51654 47142 51706
rect 47194 51654 47206 51706
rect 47258 51654 51950 51706
rect 52002 51654 52014 51706
rect 52066 51654 52078 51706
rect 52130 51654 52142 51706
rect 52194 51654 52206 51706
rect 52258 51654 56950 51706
rect 57002 51654 57014 51706
rect 57066 51654 57078 51706
rect 57130 51654 57142 51706
rect 57194 51654 57206 51706
rect 57258 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 2610 51162
rect 2662 51110 2674 51162
rect 2726 51110 2738 51162
rect 2790 51110 2802 51162
rect 2854 51110 2866 51162
rect 2918 51110 7610 51162
rect 7662 51110 7674 51162
rect 7726 51110 7738 51162
rect 7790 51110 7802 51162
rect 7854 51110 7866 51162
rect 7918 51110 12610 51162
rect 12662 51110 12674 51162
rect 12726 51110 12738 51162
rect 12790 51110 12802 51162
rect 12854 51110 12866 51162
rect 12918 51110 17610 51162
rect 17662 51110 17674 51162
rect 17726 51110 17738 51162
rect 17790 51110 17802 51162
rect 17854 51110 17866 51162
rect 17918 51110 22610 51162
rect 22662 51110 22674 51162
rect 22726 51110 22738 51162
rect 22790 51110 22802 51162
rect 22854 51110 22866 51162
rect 22918 51110 27610 51162
rect 27662 51110 27674 51162
rect 27726 51110 27738 51162
rect 27790 51110 27802 51162
rect 27854 51110 27866 51162
rect 27918 51110 32610 51162
rect 32662 51110 32674 51162
rect 32726 51110 32738 51162
rect 32790 51110 32802 51162
rect 32854 51110 32866 51162
rect 32918 51110 37610 51162
rect 37662 51110 37674 51162
rect 37726 51110 37738 51162
rect 37790 51110 37802 51162
rect 37854 51110 37866 51162
rect 37918 51110 42610 51162
rect 42662 51110 42674 51162
rect 42726 51110 42738 51162
rect 42790 51110 42802 51162
rect 42854 51110 42866 51162
rect 42918 51110 47610 51162
rect 47662 51110 47674 51162
rect 47726 51110 47738 51162
rect 47790 51110 47802 51162
rect 47854 51110 47866 51162
rect 47918 51110 52610 51162
rect 52662 51110 52674 51162
rect 52726 51110 52738 51162
rect 52790 51110 52802 51162
rect 52854 51110 52866 51162
rect 52918 51110 57610 51162
rect 57662 51110 57674 51162
rect 57726 51110 57738 51162
rect 57790 51110 57802 51162
rect 57854 51110 57866 51162
rect 57918 51110 58880 51162
rect 1104 51088 58880 51110
rect 58526 50668 58532 50720
rect 58584 50668 58590 50720
rect 1104 50618 58880 50640
rect 1104 50566 1950 50618
rect 2002 50566 2014 50618
rect 2066 50566 2078 50618
rect 2130 50566 2142 50618
rect 2194 50566 2206 50618
rect 2258 50566 6950 50618
rect 7002 50566 7014 50618
rect 7066 50566 7078 50618
rect 7130 50566 7142 50618
rect 7194 50566 7206 50618
rect 7258 50566 11950 50618
rect 12002 50566 12014 50618
rect 12066 50566 12078 50618
rect 12130 50566 12142 50618
rect 12194 50566 12206 50618
rect 12258 50566 16950 50618
rect 17002 50566 17014 50618
rect 17066 50566 17078 50618
rect 17130 50566 17142 50618
rect 17194 50566 17206 50618
rect 17258 50566 21950 50618
rect 22002 50566 22014 50618
rect 22066 50566 22078 50618
rect 22130 50566 22142 50618
rect 22194 50566 22206 50618
rect 22258 50566 26950 50618
rect 27002 50566 27014 50618
rect 27066 50566 27078 50618
rect 27130 50566 27142 50618
rect 27194 50566 27206 50618
rect 27258 50566 31950 50618
rect 32002 50566 32014 50618
rect 32066 50566 32078 50618
rect 32130 50566 32142 50618
rect 32194 50566 32206 50618
rect 32258 50566 36950 50618
rect 37002 50566 37014 50618
rect 37066 50566 37078 50618
rect 37130 50566 37142 50618
rect 37194 50566 37206 50618
rect 37258 50566 41950 50618
rect 42002 50566 42014 50618
rect 42066 50566 42078 50618
rect 42130 50566 42142 50618
rect 42194 50566 42206 50618
rect 42258 50566 46950 50618
rect 47002 50566 47014 50618
rect 47066 50566 47078 50618
rect 47130 50566 47142 50618
rect 47194 50566 47206 50618
rect 47258 50566 51950 50618
rect 52002 50566 52014 50618
rect 52066 50566 52078 50618
rect 52130 50566 52142 50618
rect 52194 50566 52206 50618
rect 52258 50566 56950 50618
rect 57002 50566 57014 50618
rect 57066 50566 57078 50618
rect 57130 50566 57142 50618
rect 57194 50566 57206 50618
rect 57258 50566 58880 50618
rect 1104 50544 58880 50566
rect 58526 50260 58532 50312
rect 58584 50260 58590 50312
rect 1104 50074 58880 50096
rect 1104 50022 2610 50074
rect 2662 50022 2674 50074
rect 2726 50022 2738 50074
rect 2790 50022 2802 50074
rect 2854 50022 2866 50074
rect 2918 50022 7610 50074
rect 7662 50022 7674 50074
rect 7726 50022 7738 50074
rect 7790 50022 7802 50074
rect 7854 50022 7866 50074
rect 7918 50022 12610 50074
rect 12662 50022 12674 50074
rect 12726 50022 12738 50074
rect 12790 50022 12802 50074
rect 12854 50022 12866 50074
rect 12918 50022 17610 50074
rect 17662 50022 17674 50074
rect 17726 50022 17738 50074
rect 17790 50022 17802 50074
rect 17854 50022 17866 50074
rect 17918 50022 22610 50074
rect 22662 50022 22674 50074
rect 22726 50022 22738 50074
rect 22790 50022 22802 50074
rect 22854 50022 22866 50074
rect 22918 50022 27610 50074
rect 27662 50022 27674 50074
rect 27726 50022 27738 50074
rect 27790 50022 27802 50074
rect 27854 50022 27866 50074
rect 27918 50022 32610 50074
rect 32662 50022 32674 50074
rect 32726 50022 32738 50074
rect 32790 50022 32802 50074
rect 32854 50022 32866 50074
rect 32918 50022 37610 50074
rect 37662 50022 37674 50074
rect 37726 50022 37738 50074
rect 37790 50022 37802 50074
rect 37854 50022 37866 50074
rect 37918 50022 42610 50074
rect 42662 50022 42674 50074
rect 42726 50022 42738 50074
rect 42790 50022 42802 50074
rect 42854 50022 42866 50074
rect 42918 50022 47610 50074
rect 47662 50022 47674 50074
rect 47726 50022 47738 50074
rect 47790 50022 47802 50074
rect 47854 50022 47866 50074
rect 47918 50022 52610 50074
rect 52662 50022 52674 50074
rect 52726 50022 52738 50074
rect 52790 50022 52802 50074
rect 52854 50022 52866 50074
rect 52918 50022 57610 50074
rect 57662 50022 57674 50074
rect 57726 50022 57738 50074
rect 57790 50022 57802 50074
rect 57854 50022 57866 50074
rect 57918 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 1950 49530
rect 2002 49478 2014 49530
rect 2066 49478 2078 49530
rect 2130 49478 2142 49530
rect 2194 49478 2206 49530
rect 2258 49478 6950 49530
rect 7002 49478 7014 49530
rect 7066 49478 7078 49530
rect 7130 49478 7142 49530
rect 7194 49478 7206 49530
rect 7258 49478 11950 49530
rect 12002 49478 12014 49530
rect 12066 49478 12078 49530
rect 12130 49478 12142 49530
rect 12194 49478 12206 49530
rect 12258 49478 16950 49530
rect 17002 49478 17014 49530
rect 17066 49478 17078 49530
rect 17130 49478 17142 49530
rect 17194 49478 17206 49530
rect 17258 49478 21950 49530
rect 22002 49478 22014 49530
rect 22066 49478 22078 49530
rect 22130 49478 22142 49530
rect 22194 49478 22206 49530
rect 22258 49478 26950 49530
rect 27002 49478 27014 49530
rect 27066 49478 27078 49530
rect 27130 49478 27142 49530
rect 27194 49478 27206 49530
rect 27258 49478 31950 49530
rect 32002 49478 32014 49530
rect 32066 49478 32078 49530
rect 32130 49478 32142 49530
rect 32194 49478 32206 49530
rect 32258 49478 36950 49530
rect 37002 49478 37014 49530
rect 37066 49478 37078 49530
rect 37130 49478 37142 49530
rect 37194 49478 37206 49530
rect 37258 49478 41950 49530
rect 42002 49478 42014 49530
rect 42066 49478 42078 49530
rect 42130 49478 42142 49530
rect 42194 49478 42206 49530
rect 42258 49478 46950 49530
rect 47002 49478 47014 49530
rect 47066 49478 47078 49530
rect 47130 49478 47142 49530
rect 47194 49478 47206 49530
rect 47258 49478 51950 49530
rect 52002 49478 52014 49530
rect 52066 49478 52078 49530
rect 52130 49478 52142 49530
rect 52194 49478 52206 49530
rect 52258 49478 56950 49530
rect 57002 49478 57014 49530
rect 57066 49478 57078 49530
rect 57130 49478 57142 49530
rect 57194 49478 57206 49530
rect 57258 49478 58880 49530
rect 1104 49456 58880 49478
rect 58526 49172 58532 49224
rect 58584 49172 58590 49224
rect 1104 48986 58880 49008
rect 1104 48934 2610 48986
rect 2662 48934 2674 48986
rect 2726 48934 2738 48986
rect 2790 48934 2802 48986
rect 2854 48934 2866 48986
rect 2918 48934 7610 48986
rect 7662 48934 7674 48986
rect 7726 48934 7738 48986
rect 7790 48934 7802 48986
rect 7854 48934 7866 48986
rect 7918 48934 12610 48986
rect 12662 48934 12674 48986
rect 12726 48934 12738 48986
rect 12790 48934 12802 48986
rect 12854 48934 12866 48986
rect 12918 48934 17610 48986
rect 17662 48934 17674 48986
rect 17726 48934 17738 48986
rect 17790 48934 17802 48986
rect 17854 48934 17866 48986
rect 17918 48934 22610 48986
rect 22662 48934 22674 48986
rect 22726 48934 22738 48986
rect 22790 48934 22802 48986
rect 22854 48934 22866 48986
rect 22918 48934 27610 48986
rect 27662 48934 27674 48986
rect 27726 48934 27738 48986
rect 27790 48934 27802 48986
rect 27854 48934 27866 48986
rect 27918 48934 32610 48986
rect 32662 48934 32674 48986
rect 32726 48934 32738 48986
rect 32790 48934 32802 48986
rect 32854 48934 32866 48986
rect 32918 48934 37610 48986
rect 37662 48934 37674 48986
rect 37726 48934 37738 48986
rect 37790 48934 37802 48986
rect 37854 48934 37866 48986
rect 37918 48934 42610 48986
rect 42662 48934 42674 48986
rect 42726 48934 42738 48986
rect 42790 48934 42802 48986
rect 42854 48934 42866 48986
rect 42918 48934 47610 48986
rect 47662 48934 47674 48986
rect 47726 48934 47738 48986
rect 47790 48934 47802 48986
rect 47854 48934 47866 48986
rect 47918 48934 52610 48986
rect 52662 48934 52674 48986
rect 52726 48934 52738 48986
rect 52790 48934 52802 48986
rect 52854 48934 52866 48986
rect 52918 48934 57610 48986
rect 57662 48934 57674 48986
rect 57726 48934 57738 48986
rect 57790 48934 57802 48986
rect 57854 48934 57866 48986
rect 57918 48934 58880 48986
rect 1104 48912 58880 48934
rect 58526 48492 58532 48544
rect 58584 48492 58590 48544
rect 1104 48442 58880 48464
rect 1104 48390 1950 48442
rect 2002 48390 2014 48442
rect 2066 48390 2078 48442
rect 2130 48390 2142 48442
rect 2194 48390 2206 48442
rect 2258 48390 6950 48442
rect 7002 48390 7014 48442
rect 7066 48390 7078 48442
rect 7130 48390 7142 48442
rect 7194 48390 7206 48442
rect 7258 48390 11950 48442
rect 12002 48390 12014 48442
rect 12066 48390 12078 48442
rect 12130 48390 12142 48442
rect 12194 48390 12206 48442
rect 12258 48390 16950 48442
rect 17002 48390 17014 48442
rect 17066 48390 17078 48442
rect 17130 48390 17142 48442
rect 17194 48390 17206 48442
rect 17258 48390 21950 48442
rect 22002 48390 22014 48442
rect 22066 48390 22078 48442
rect 22130 48390 22142 48442
rect 22194 48390 22206 48442
rect 22258 48390 26950 48442
rect 27002 48390 27014 48442
rect 27066 48390 27078 48442
rect 27130 48390 27142 48442
rect 27194 48390 27206 48442
rect 27258 48390 31950 48442
rect 32002 48390 32014 48442
rect 32066 48390 32078 48442
rect 32130 48390 32142 48442
rect 32194 48390 32206 48442
rect 32258 48390 36950 48442
rect 37002 48390 37014 48442
rect 37066 48390 37078 48442
rect 37130 48390 37142 48442
rect 37194 48390 37206 48442
rect 37258 48390 41950 48442
rect 42002 48390 42014 48442
rect 42066 48390 42078 48442
rect 42130 48390 42142 48442
rect 42194 48390 42206 48442
rect 42258 48390 46950 48442
rect 47002 48390 47014 48442
rect 47066 48390 47078 48442
rect 47130 48390 47142 48442
rect 47194 48390 47206 48442
rect 47258 48390 51950 48442
rect 52002 48390 52014 48442
rect 52066 48390 52078 48442
rect 52130 48390 52142 48442
rect 52194 48390 52206 48442
rect 52258 48390 56950 48442
rect 57002 48390 57014 48442
rect 57066 48390 57078 48442
rect 57130 48390 57142 48442
rect 57194 48390 57206 48442
rect 57258 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 2610 47898
rect 2662 47846 2674 47898
rect 2726 47846 2738 47898
rect 2790 47846 2802 47898
rect 2854 47846 2866 47898
rect 2918 47846 7610 47898
rect 7662 47846 7674 47898
rect 7726 47846 7738 47898
rect 7790 47846 7802 47898
rect 7854 47846 7866 47898
rect 7918 47846 12610 47898
rect 12662 47846 12674 47898
rect 12726 47846 12738 47898
rect 12790 47846 12802 47898
rect 12854 47846 12866 47898
rect 12918 47846 17610 47898
rect 17662 47846 17674 47898
rect 17726 47846 17738 47898
rect 17790 47846 17802 47898
rect 17854 47846 17866 47898
rect 17918 47846 22610 47898
rect 22662 47846 22674 47898
rect 22726 47846 22738 47898
rect 22790 47846 22802 47898
rect 22854 47846 22866 47898
rect 22918 47846 27610 47898
rect 27662 47846 27674 47898
rect 27726 47846 27738 47898
rect 27790 47846 27802 47898
rect 27854 47846 27866 47898
rect 27918 47846 32610 47898
rect 32662 47846 32674 47898
rect 32726 47846 32738 47898
rect 32790 47846 32802 47898
rect 32854 47846 32866 47898
rect 32918 47846 37610 47898
rect 37662 47846 37674 47898
rect 37726 47846 37738 47898
rect 37790 47846 37802 47898
rect 37854 47846 37866 47898
rect 37918 47846 42610 47898
rect 42662 47846 42674 47898
rect 42726 47846 42738 47898
rect 42790 47846 42802 47898
rect 42854 47846 42866 47898
rect 42918 47846 47610 47898
rect 47662 47846 47674 47898
rect 47726 47846 47738 47898
rect 47790 47846 47802 47898
rect 47854 47846 47866 47898
rect 47918 47846 52610 47898
rect 52662 47846 52674 47898
rect 52726 47846 52738 47898
rect 52790 47846 52802 47898
rect 52854 47846 52866 47898
rect 52918 47846 57610 47898
rect 57662 47846 57674 47898
rect 57726 47846 57738 47898
rect 57790 47846 57802 47898
rect 57854 47846 57866 47898
rect 57918 47846 58880 47898
rect 1104 47824 58880 47846
rect 58526 47404 58532 47456
rect 58584 47404 58590 47456
rect 1104 47354 58880 47376
rect 1104 47302 1950 47354
rect 2002 47302 2014 47354
rect 2066 47302 2078 47354
rect 2130 47302 2142 47354
rect 2194 47302 2206 47354
rect 2258 47302 6950 47354
rect 7002 47302 7014 47354
rect 7066 47302 7078 47354
rect 7130 47302 7142 47354
rect 7194 47302 7206 47354
rect 7258 47302 11950 47354
rect 12002 47302 12014 47354
rect 12066 47302 12078 47354
rect 12130 47302 12142 47354
rect 12194 47302 12206 47354
rect 12258 47302 16950 47354
rect 17002 47302 17014 47354
rect 17066 47302 17078 47354
rect 17130 47302 17142 47354
rect 17194 47302 17206 47354
rect 17258 47302 21950 47354
rect 22002 47302 22014 47354
rect 22066 47302 22078 47354
rect 22130 47302 22142 47354
rect 22194 47302 22206 47354
rect 22258 47302 26950 47354
rect 27002 47302 27014 47354
rect 27066 47302 27078 47354
rect 27130 47302 27142 47354
rect 27194 47302 27206 47354
rect 27258 47302 31950 47354
rect 32002 47302 32014 47354
rect 32066 47302 32078 47354
rect 32130 47302 32142 47354
rect 32194 47302 32206 47354
rect 32258 47302 36950 47354
rect 37002 47302 37014 47354
rect 37066 47302 37078 47354
rect 37130 47302 37142 47354
rect 37194 47302 37206 47354
rect 37258 47302 41950 47354
rect 42002 47302 42014 47354
rect 42066 47302 42078 47354
rect 42130 47302 42142 47354
rect 42194 47302 42206 47354
rect 42258 47302 46950 47354
rect 47002 47302 47014 47354
rect 47066 47302 47078 47354
rect 47130 47302 47142 47354
rect 47194 47302 47206 47354
rect 47258 47302 51950 47354
rect 52002 47302 52014 47354
rect 52066 47302 52078 47354
rect 52130 47302 52142 47354
rect 52194 47302 52206 47354
rect 52258 47302 56950 47354
rect 57002 47302 57014 47354
rect 57066 47302 57078 47354
rect 57130 47302 57142 47354
rect 57194 47302 57206 47354
rect 57258 47302 58880 47354
rect 1104 47280 58880 47302
rect 58526 46996 58532 47048
rect 58584 46996 58590 47048
rect 1104 46810 58880 46832
rect 1104 46758 2610 46810
rect 2662 46758 2674 46810
rect 2726 46758 2738 46810
rect 2790 46758 2802 46810
rect 2854 46758 2866 46810
rect 2918 46758 7610 46810
rect 7662 46758 7674 46810
rect 7726 46758 7738 46810
rect 7790 46758 7802 46810
rect 7854 46758 7866 46810
rect 7918 46758 12610 46810
rect 12662 46758 12674 46810
rect 12726 46758 12738 46810
rect 12790 46758 12802 46810
rect 12854 46758 12866 46810
rect 12918 46758 17610 46810
rect 17662 46758 17674 46810
rect 17726 46758 17738 46810
rect 17790 46758 17802 46810
rect 17854 46758 17866 46810
rect 17918 46758 22610 46810
rect 22662 46758 22674 46810
rect 22726 46758 22738 46810
rect 22790 46758 22802 46810
rect 22854 46758 22866 46810
rect 22918 46758 27610 46810
rect 27662 46758 27674 46810
rect 27726 46758 27738 46810
rect 27790 46758 27802 46810
rect 27854 46758 27866 46810
rect 27918 46758 32610 46810
rect 32662 46758 32674 46810
rect 32726 46758 32738 46810
rect 32790 46758 32802 46810
rect 32854 46758 32866 46810
rect 32918 46758 37610 46810
rect 37662 46758 37674 46810
rect 37726 46758 37738 46810
rect 37790 46758 37802 46810
rect 37854 46758 37866 46810
rect 37918 46758 42610 46810
rect 42662 46758 42674 46810
rect 42726 46758 42738 46810
rect 42790 46758 42802 46810
rect 42854 46758 42866 46810
rect 42918 46758 47610 46810
rect 47662 46758 47674 46810
rect 47726 46758 47738 46810
rect 47790 46758 47802 46810
rect 47854 46758 47866 46810
rect 47918 46758 52610 46810
rect 52662 46758 52674 46810
rect 52726 46758 52738 46810
rect 52790 46758 52802 46810
rect 52854 46758 52866 46810
rect 52918 46758 57610 46810
rect 57662 46758 57674 46810
rect 57726 46758 57738 46810
rect 57790 46758 57802 46810
rect 57854 46758 57866 46810
rect 57918 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 1950 46266
rect 2002 46214 2014 46266
rect 2066 46214 2078 46266
rect 2130 46214 2142 46266
rect 2194 46214 2206 46266
rect 2258 46214 6950 46266
rect 7002 46214 7014 46266
rect 7066 46214 7078 46266
rect 7130 46214 7142 46266
rect 7194 46214 7206 46266
rect 7258 46214 11950 46266
rect 12002 46214 12014 46266
rect 12066 46214 12078 46266
rect 12130 46214 12142 46266
rect 12194 46214 12206 46266
rect 12258 46214 16950 46266
rect 17002 46214 17014 46266
rect 17066 46214 17078 46266
rect 17130 46214 17142 46266
rect 17194 46214 17206 46266
rect 17258 46214 21950 46266
rect 22002 46214 22014 46266
rect 22066 46214 22078 46266
rect 22130 46214 22142 46266
rect 22194 46214 22206 46266
rect 22258 46214 26950 46266
rect 27002 46214 27014 46266
rect 27066 46214 27078 46266
rect 27130 46214 27142 46266
rect 27194 46214 27206 46266
rect 27258 46214 31950 46266
rect 32002 46214 32014 46266
rect 32066 46214 32078 46266
rect 32130 46214 32142 46266
rect 32194 46214 32206 46266
rect 32258 46214 36950 46266
rect 37002 46214 37014 46266
rect 37066 46214 37078 46266
rect 37130 46214 37142 46266
rect 37194 46214 37206 46266
rect 37258 46214 41950 46266
rect 42002 46214 42014 46266
rect 42066 46214 42078 46266
rect 42130 46214 42142 46266
rect 42194 46214 42206 46266
rect 42258 46214 46950 46266
rect 47002 46214 47014 46266
rect 47066 46214 47078 46266
rect 47130 46214 47142 46266
rect 47194 46214 47206 46266
rect 47258 46214 51950 46266
rect 52002 46214 52014 46266
rect 52066 46214 52078 46266
rect 52130 46214 52142 46266
rect 52194 46214 52206 46266
rect 52258 46214 56950 46266
rect 57002 46214 57014 46266
rect 57066 46214 57078 46266
rect 57130 46214 57142 46266
rect 57194 46214 57206 46266
rect 57258 46214 58880 46266
rect 1104 46192 58880 46214
rect 58526 45908 58532 45960
rect 58584 45908 58590 45960
rect 1104 45722 58880 45744
rect 1104 45670 2610 45722
rect 2662 45670 2674 45722
rect 2726 45670 2738 45722
rect 2790 45670 2802 45722
rect 2854 45670 2866 45722
rect 2918 45670 7610 45722
rect 7662 45670 7674 45722
rect 7726 45670 7738 45722
rect 7790 45670 7802 45722
rect 7854 45670 7866 45722
rect 7918 45670 12610 45722
rect 12662 45670 12674 45722
rect 12726 45670 12738 45722
rect 12790 45670 12802 45722
rect 12854 45670 12866 45722
rect 12918 45670 17610 45722
rect 17662 45670 17674 45722
rect 17726 45670 17738 45722
rect 17790 45670 17802 45722
rect 17854 45670 17866 45722
rect 17918 45670 22610 45722
rect 22662 45670 22674 45722
rect 22726 45670 22738 45722
rect 22790 45670 22802 45722
rect 22854 45670 22866 45722
rect 22918 45670 27610 45722
rect 27662 45670 27674 45722
rect 27726 45670 27738 45722
rect 27790 45670 27802 45722
rect 27854 45670 27866 45722
rect 27918 45670 32610 45722
rect 32662 45670 32674 45722
rect 32726 45670 32738 45722
rect 32790 45670 32802 45722
rect 32854 45670 32866 45722
rect 32918 45670 37610 45722
rect 37662 45670 37674 45722
rect 37726 45670 37738 45722
rect 37790 45670 37802 45722
rect 37854 45670 37866 45722
rect 37918 45670 42610 45722
rect 42662 45670 42674 45722
rect 42726 45670 42738 45722
rect 42790 45670 42802 45722
rect 42854 45670 42866 45722
rect 42918 45670 47610 45722
rect 47662 45670 47674 45722
rect 47726 45670 47738 45722
rect 47790 45670 47802 45722
rect 47854 45670 47866 45722
rect 47918 45670 52610 45722
rect 52662 45670 52674 45722
rect 52726 45670 52738 45722
rect 52790 45670 52802 45722
rect 52854 45670 52866 45722
rect 52918 45670 57610 45722
rect 57662 45670 57674 45722
rect 57726 45670 57738 45722
rect 57790 45670 57802 45722
rect 57854 45670 57866 45722
rect 57918 45670 58880 45722
rect 1104 45648 58880 45670
rect 58526 45228 58532 45280
rect 58584 45228 58590 45280
rect 1104 45178 58880 45200
rect 1104 45126 1950 45178
rect 2002 45126 2014 45178
rect 2066 45126 2078 45178
rect 2130 45126 2142 45178
rect 2194 45126 2206 45178
rect 2258 45126 6950 45178
rect 7002 45126 7014 45178
rect 7066 45126 7078 45178
rect 7130 45126 7142 45178
rect 7194 45126 7206 45178
rect 7258 45126 11950 45178
rect 12002 45126 12014 45178
rect 12066 45126 12078 45178
rect 12130 45126 12142 45178
rect 12194 45126 12206 45178
rect 12258 45126 16950 45178
rect 17002 45126 17014 45178
rect 17066 45126 17078 45178
rect 17130 45126 17142 45178
rect 17194 45126 17206 45178
rect 17258 45126 21950 45178
rect 22002 45126 22014 45178
rect 22066 45126 22078 45178
rect 22130 45126 22142 45178
rect 22194 45126 22206 45178
rect 22258 45126 26950 45178
rect 27002 45126 27014 45178
rect 27066 45126 27078 45178
rect 27130 45126 27142 45178
rect 27194 45126 27206 45178
rect 27258 45126 31950 45178
rect 32002 45126 32014 45178
rect 32066 45126 32078 45178
rect 32130 45126 32142 45178
rect 32194 45126 32206 45178
rect 32258 45126 36950 45178
rect 37002 45126 37014 45178
rect 37066 45126 37078 45178
rect 37130 45126 37142 45178
rect 37194 45126 37206 45178
rect 37258 45126 41950 45178
rect 42002 45126 42014 45178
rect 42066 45126 42078 45178
rect 42130 45126 42142 45178
rect 42194 45126 42206 45178
rect 42258 45126 46950 45178
rect 47002 45126 47014 45178
rect 47066 45126 47078 45178
rect 47130 45126 47142 45178
rect 47194 45126 47206 45178
rect 47258 45126 51950 45178
rect 52002 45126 52014 45178
rect 52066 45126 52078 45178
rect 52130 45126 52142 45178
rect 52194 45126 52206 45178
rect 52258 45126 56950 45178
rect 57002 45126 57014 45178
rect 57066 45126 57078 45178
rect 57130 45126 57142 45178
rect 57194 45126 57206 45178
rect 57258 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 2610 44634
rect 2662 44582 2674 44634
rect 2726 44582 2738 44634
rect 2790 44582 2802 44634
rect 2854 44582 2866 44634
rect 2918 44582 7610 44634
rect 7662 44582 7674 44634
rect 7726 44582 7738 44634
rect 7790 44582 7802 44634
rect 7854 44582 7866 44634
rect 7918 44582 12610 44634
rect 12662 44582 12674 44634
rect 12726 44582 12738 44634
rect 12790 44582 12802 44634
rect 12854 44582 12866 44634
rect 12918 44582 17610 44634
rect 17662 44582 17674 44634
rect 17726 44582 17738 44634
rect 17790 44582 17802 44634
rect 17854 44582 17866 44634
rect 17918 44582 22610 44634
rect 22662 44582 22674 44634
rect 22726 44582 22738 44634
rect 22790 44582 22802 44634
rect 22854 44582 22866 44634
rect 22918 44582 27610 44634
rect 27662 44582 27674 44634
rect 27726 44582 27738 44634
rect 27790 44582 27802 44634
rect 27854 44582 27866 44634
rect 27918 44582 32610 44634
rect 32662 44582 32674 44634
rect 32726 44582 32738 44634
rect 32790 44582 32802 44634
rect 32854 44582 32866 44634
rect 32918 44582 37610 44634
rect 37662 44582 37674 44634
rect 37726 44582 37738 44634
rect 37790 44582 37802 44634
rect 37854 44582 37866 44634
rect 37918 44582 42610 44634
rect 42662 44582 42674 44634
rect 42726 44582 42738 44634
rect 42790 44582 42802 44634
rect 42854 44582 42866 44634
rect 42918 44582 47610 44634
rect 47662 44582 47674 44634
rect 47726 44582 47738 44634
rect 47790 44582 47802 44634
rect 47854 44582 47866 44634
rect 47918 44582 52610 44634
rect 52662 44582 52674 44634
rect 52726 44582 52738 44634
rect 52790 44582 52802 44634
rect 52854 44582 52866 44634
rect 52918 44582 57610 44634
rect 57662 44582 57674 44634
rect 57726 44582 57738 44634
rect 57790 44582 57802 44634
rect 57854 44582 57866 44634
rect 57918 44582 58880 44634
rect 1104 44560 58880 44582
rect 58526 44140 58532 44192
rect 58584 44140 58590 44192
rect 1104 44090 58880 44112
rect 1104 44038 1950 44090
rect 2002 44038 2014 44090
rect 2066 44038 2078 44090
rect 2130 44038 2142 44090
rect 2194 44038 2206 44090
rect 2258 44038 6950 44090
rect 7002 44038 7014 44090
rect 7066 44038 7078 44090
rect 7130 44038 7142 44090
rect 7194 44038 7206 44090
rect 7258 44038 11950 44090
rect 12002 44038 12014 44090
rect 12066 44038 12078 44090
rect 12130 44038 12142 44090
rect 12194 44038 12206 44090
rect 12258 44038 16950 44090
rect 17002 44038 17014 44090
rect 17066 44038 17078 44090
rect 17130 44038 17142 44090
rect 17194 44038 17206 44090
rect 17258 44038 21950 44090
rect 22002 44038 22014 44090
rect 22066 44038 22078 44090
rect 22130 44038 22142 44090
rect 22194 44038 22206 44090
rect 22258 44038 26950 44090
rect 27002 44038 27014 44090
rect 27066 44038 27078 44090
rect 27130 44038 27142 44090
rect 27194 44038 27206 44090
rect 27258 44038 31950 44090
rect 32002 44038 32014 44090
rect 32066 44038 32078 44090
rect 32130 44038 32142 44090
rect 32194 44038 32206 44090
rect 32258 44038 36950 44090
rect 37002 44038 37014 44090
rect 37066 44038 37078 44090
rect 37130 44038 37142 44090
rect 37194 44038 37206 44090
rect 37258 44038 41950 44090
rect 42002 44038 42014 44090
rect 42066 44038 42078 44090
rect 42130 44038 42142 44090
rect 42194 44038 42206 44090
rect 42258 44038 46950 44090
rect 47002 44038 47014 44090
rect 47066 44038 47078 44090
rect 47130 44038 47142 44090
rect 47194 44038 47206 44090
rect 47258 44038 51950 44090
rect 52002 44038 52014 44090
rect 52066 44038 52078 44090
rect 52130 44038 52142 44090
rect 52194 44038 52206 44090
rect 52258 44038 56950 44090
rect 57002 44038 57014 44090
rect 57066 44038 57078 44090
rect 57130 44038 57142 44090
rect 57194 44038 57206 44090
rect 57258 44038 58880 44090
rect 1104 44016 58880 44038
rect 58526 43732 58532 43784
rect 58584 43732 58590 43784
rect 1104 43546 58880 43568
rect 1104 43494 2610 43546
rect 2662 43494 2674 43546
rect 2726 43494 2738 43546
rect 2790 43494 2802 43546
rect 2854 43494 2866 43546
rect 2918 43494 7610 43546
rect 7662 43494 7674 43546
rect 7726 43494 7738 43546
rect 7790 43494 7802 43546
rect 7854 43494 7866 43546
rect 7918 43494 12610 43546
rect 12662 43494 12674 43546
rect 12726 43494 12738 43546
rect 12790 43494 12802 43546
rect 12854 43494 12866 43546
rect 12918 43494 17610 43546
rect 17662 43494 17674 43546
rect 17726 43494 17738 43546
rect 17790 43494 17802 43546
rect 17854 43494 17866 43546
rect 17918 43494 22610 43546
rect 22662 43494 22674 43546
rect 22726 43494 22738 43546
rect 22790 43494 22802 43546
rect 22854 43494 22866 43546
rect 22918 43494 27610 43546
rect 27662 43494 27674 43546
rect 27726 43494 27738 43546
rect 27790 43494 27802 43546
rect 27854 43494 27866 43546
rect 27918 43494 32610 43546
rect 32662 43494 32674 43546
rect 32726 43494 32738 43546
rect 32790 43494 32802 43546
rect 32854 43494 32866 43546
rect 32918 43494 37610 43546
rect 37662 43494 37674 43546
rect 37726 43494 37738 43546
rect 37790 43494 37802 43546
rect 37854 43494 37866 43546
rect 37918 43494 42610 43546
rect 42662 43494 42674 43546
rect 42726 43494 42738 43546
rect 42790 43494 42802 43546
rect 42854 43494 42866 43546
rect 42918 43494 47610 43546
rect 47662 43494 47674 43546
rect 47726 43494 47738 43546
rect 47790 43494 47802 43546
rect 47854 43494 47866 43546
rect 47918 43494 52610 43546
rect 52662 43494 52674 43546
rect 52726 43494 52738 43546
rect 52790 43494 52802 43546
rect 52854 43494 52866 43546
rect 52918 43494 57610 43546
rect 57662 43494 57674 43546
rect 57726 43494 57738 43546
rect 57790 43494 57802 43546
rect 57854 43494 57866 43546
rect 57918 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 1950 43002
rect 2002 42950 2014 43002
rect 2066 42950 2078 43002
rect 2130 42950 2142 43002
rect 2194 42950 2206 43002
rect 2258 42950 6950 43002
rect 7002 42950 7014 43002
rect 7066 42950 7078 43002
rect 7130 42950 7142 43002
rect 7194 42950 7206 43002
rect 7258 42950 11950 43002
rect 12002 42950 12014 43002
rect 12066 42950 12078 43002
rect 12130 42950 12142 43002
rect 12194 42950 12206 43002
rect 12258 42950 16950 43002
rect 17002 42950 17014 43002
rect 17066 42950 17078 43002
rect 17130 42950 17142 43002
rect 17194 42950 17206 43002
rect 17258 42950 21950 43002
rect 22002 42950 22014 43002
rect 22066 42950 22078 43002
rect 22130 42950 22142 43002
rect 22194 42950 22206 43002
rect 22258 42950 26950 43002
rect 27002 42950 27014 43002
rect 27066 42950 27078 43002
rect 27130 42950 27142 43002
rect 27194 42950 27206 43002
rect 27258 42950 31950 43002
rect 32002 42950 32014 43002
rect 32066 42950 32078 43002
rect 32130 42950 32142 43002
rect 32194 42950 32206 43002
rect 32258 42950 36950 43002
rect 37002 42950 37014 43002
rect 37066 42950 37078 43002
rect 37130 42950 37142 43002
rect 37194 42950 37206 43002
rect 37258 42950 41950 43002
rect 42002 42950 42014 43002
rect 42066 42950 42078 43002
rect 42130 42950 42142 43002
rect 42194 42950 42206 43002
rect 42258 42950 46950 43002
rect 47002 42950 47014 43002
rect 47066 42950 47078 43002
rect 47130 42950 47142 43002
rect 47194 42950 47206 43002
rect 47258 42950 51950 43002
rect 52002 42950 52014 43002
rect 52066 42950 52078 43002
rect 52130 42950 52142 43002
rect 52194 42950 52206 43002
rect 52258 42950 56950 43002
rect 57002 42950 57014 43002
rect 57066 42950 57078 43002
rect 57130 42950 57142 43002
rect 57194 42950 57206 43002
rect 57258 42950 58880 43002
rect 1104 42928 58880 42950
rect 58526 42644 58532 42696
rect 58584 42644 58590 42696
rect 1104 42458 58880 42480
rect 1104 42406 2610 42458
rect 2662 42406 2674 42458
rect 2726 42406 2738 42458
rect 2790 42406 2802 42458
rect 2854 42406 2866 42458
rect 2918 42406 7610 42458
rect 7662 42406 7674 42458
rect 7726 42406 7738 42458
rect 7790 42406 7802 42458
rect 7854 42406 7866 42458
rect 7918 42406 12610 42458
rect 12662 42406 12674 42458
rect 12726 42406 12738 42458
rect 12790 42406 12802 42458
rect 12854 42406 12866 42458
rect 12918 42406 17610 42458
rect 17662 42406 17674 42458
rect 17726 42406 17738 42458
rect 17790 42406 17802 42458
rect 17854 42406 17866 42458
rect 17918 42406 22610 42458
rect 22662 42406 22674 42458
rect 22726 42406 22738 42458
rect 22790 42406 22802 42458
rect 22854 42406 22866 42458
rect 22918 42406 27610 42458
rect 27662 42406 27674 42458
rect 27726 42406 27738 42458
rect 27790 42406 27802 42458
rect 27854 42406 27866 42458
rect 27918 42406 32610 42458
rect 32662 42406 32674 42458
rect 32726 42406 32738 42458
rect 32790 42406 32802 42458
rect 32854 42406 32866 42458
rect 32918 42406 37610 42458
rect 37662 42406 37674 42458
rect 37726 42406 37738 42458
rect 37790 42406 37802 42458
rect 37854 42406 37866 42458
rect 37918 42406 42610 42458
rect 42662 42406 42674 42458
rect 42726 42406 42738 42458
rect 42790 42406 42802 42458
rect 42854 42406 42866 42458
rect 42918 42406 47610 42458
rect 47662 42406 47674 42458
rect 47726 42406 47738 42458
rect 47790 42406 47802 42458
rect 47854 42406 47866 42458
rect 47918 42406 52610 42458
rect 52662 42406 52674 42458
rect 52726 42406 52738 42458
rect 52790 42406 52802 42458
rect 52854 42406 52866 42458
rect 52918 42406 57610 42458
rect 57662 42406 57674 42458
rect 57726 42406 57738 42458
rect 57790 42406 57802 42458
rect 57854 42406 57866 42458
rect 57918 42406 58880 42458
rect 1104 42384 58880 42406
rect 58526 41964 58532 42016
rect 58584 41964 58590 42016
rect 1104 41914 58880 41936
rect 1104 41862 1950 41914
rect 2002 41862 2014 41914
rect 2066 41862 2078 41914
rect 2130 41862 2142 41914
rect 2194 41862 2206 41914
rect 2258 41862 6950 41914
rect 7002 41862 7014 41914
rect 7066 41862 7078 41914
rect 7130 41862 7142 41914
rect 7194 41862 7206 41914
rect 7258 41862 11950 41914
rect 12002 41862 12014 41914
rect 12066 41862 12078 41914
rect 12130 41862 12142 41914
rect 12194 41862 12206 41914
rect 12258 41862 16950 41914
rect 17002 41862 17014 41914
rect 17066 41862 17078 41914
rect 17130 41862 17142 41914
rect 17194 41862 17206 41914
rect 17258 41862 21950 41914
rect 22002 41862 22014 41914
rect 22066 41862 22078 41914
rect 22130 41862 22142 41914
rect 22194 41862 22206 41914
rect 22258 41862 26950 41914
rect 27002 41862 27014 41914
rect 27066 41862 27078 41914
rect 27130 41862 27142 41914
rect 27194 41862 27206 41914
rect 27258 41862 31950 41914
rect 32002 41862 32014 41914
rect 32066 41862 32078 41914
rect 32130 41862 32142 41914
rect 32194 41862 32206 41914
rect 32258 41862 36950 41914
rect 37002 41862 37014 41914
rect 37066 41862 37078 41914
rect 37130 41862 37142 41914
rect 37194 41862 37206 41914
rect 37258 41862 41950 41914
rect 42002 41862 42014 41914
rect 42066 41862 42078 41914
rect 42130 41862 42142 41914
rect 42194 41862 42206 41914
rect 42258 41862 46950 41914
rect 47002 41862 47014 41914
rect 47066 41862 47078 41914
rect 47130 41862 47142 41914
rect 47194 41862 47206 41914
rect 47258 41862 51950 41914
rect 52002 41862 52014 41914
rect 52066 41862 52078 41914
rect 52130 41862 52142 41914
rect 52194 41862 52206 41914
rect 52258 41862 56950 41914
rect 57002 41862 57014 41914
rect 57066 41862 57078 41914
rect 57130 41862 57142 41914
rect 57194 41862 57206 41914
rect 57258 41862 58880 41914
rect 1104 41840 58880 41862
rect 1104 41370 58880 41392
rect 1104 41318 2610 41370
rect 2662 41318 2674 41370
rect 2726 41318 2738 41370
rect 2790 41318 2802 41370
rect 2854 41318 2866 41370
rect 2918 41318 7610 41370
rect 7662 41318 7674 41370
rect 7726 41318 7738 41370
rect 7790 41318 7802 41370
rect 7854 41318 7866 41370
rect 7918 41318 12610 41370
rect 12662 41318 12674 41370
rect 12726 41318 12738 41370
rect 12790 41318 12802 41370
rect 12854 41318 12866 41370
rect 12918 41318 17610 41370
rect 17662 41318 17674 41370
rect 17726 41318 17738 41370
rect 17790 41318 17802 41370
rect 17854 41318 17866 41370
rect 17918 41318 22610 41370
rect 22662 41318 22674 41370
rect 22726 41318 22738 41370
rect 22790 41318 22802 41370
rect 22854 41318 22866 41370
rect 22918 41318 27610 41370
rect 27662 41318 27674 41370
rect 27726 41318 27738 41370
rect 27790 41318 27802 41370
rect 27854 41318 27866 41370
rect 27918 41318 32610 41370
rect 32662 41318 32674 41370
rect 32726 41318 32738 41370
rect 32790 41318 32802 41370
rect 32854 41318 32866 41370
rect 32918 41318 37610 41370
rect 37662 41318 37674 41370
rect 37726 41318 37738 41370
rect 37790 41318 37802 41370
rect 37854 41318 37866 41370
rect 37918 41318 42610 41370
rect 42662 41318 42674 41370
rect 42726 41318 42738 41370
rect 42790 41318 42802 41370
rect 42854 41318 42866 41370
rect 42918 41318 47610 41370
rect 47662 41318 47674 41370
rect 47726 41318 47738 41370
rect 47790 41318 47802 41370
rect 47854 41318 47866 41370
rect 47918 41318 52610 41370
rect 52662 41318 52674 41370
rect 52726 41318 52738 41370
rect 52790 41318 52802 41370
rect 52854 41318 52866 41370
rect 52918 41318 57610 41370
rect 57662 41318 57674 41370
rect 57726 41318 57738 41370
rect 57790 41318 57802 41370
rect 57854 41318 57866 41370
rect 57918 41318 58880 41370
rect 1104 41296 58880 41318
rect 58526 40876 58532 40928
rect 58584 40876 58590 40928
rect 1104 40826 58880 40848
rect 1104 40774 1950 40826
rect 2002 40774 2014 40826
rect 2066 40774 2078 40826
rect 2130 40774 2142 40826
rect 2194 40774 2206 40826
rect 2258 40774 6950 40826
rect 7002 40774 7014 40826
rect 7066 40774 7078 40826
rect 7130 40774 7142 40826
rect 7194 40774 7206 40826
rect 7258 40774 11950 40826
rect 12002 40774 12014 40826
rect 12066 40774 12078 40826
rect 12130 40774 12142 40826
rect 12194 40774 12206 40826
rect 12258 40774 16950 40826
rect 17002 40774 17014 40826
rect 17066 40774 17078 40826
rect 17130 40774 17142 40826
rect 17194 40774 17206 40826
rect 17258 40774 21950 40826
rect 22002 40774 22014 40826
rect 22066 40774 22078 40826
rect 22130 40774 22142 40826
rect 22194 40774 22206 40826
rect 22258 40774 26950 40826
rect 27002 40774 27014 40826
rect 27066 40774 27078 40826
rect 27130 40774 27142 40826
rect 27194 40774 27206 40826
rect 27258 40774 31950 40826
rect 32002 40774 32014 40826
rect 32066 40774 32078 40826
rect 32130 40774 32142 40826
rect 32194 40774 32206 40826
rect 32258 40774 36950 40826
rect 37002 40774 37014 40826
rect 37066 40774 37078 40826
rect 37130 40774 37142 40826
rect 37194 40774 37206 40826
rect 37258 40774 41950 40826
rect 42002 40774 42014 40826
rect 42066 40774 42078 40826
rect 42130 40774 42142 40826
rect 42194 40774 42206 40826
rect 42258 40774 46950 40826
rect 47002 40774 47014 40826
rect 47066 40774 47078 40826
rect 47130 40774 47142 40826
rect 47194 40774 47206 40826
rect 47258 40774 51950 40826
rect 52002 40774 52014 40826
rect 52066 40774 52078 40826
rect 52130 40774 52142 40826
rect 52194 40774 52206 40826
rect 52258 40774 56950 40826
rect 57002 40774 57014 40826
rect 57066 40774 57078 40826
rect 57130 40774 57142 40826
rect 57194 40774 57206 40826
rect 57258 40774 58880 40826
rect 1104 40752 58880 40774
rect 58526 40468 58532 40520
rect 58584 40468 58590 40520
rect 1104 40282 58880 40304
rect 1104 40230 2610 40282
rect 2662 40230 2674 40282
rect 2726 40230 2738 40282
rect 2790 40230 2802 40282
rect 2854 40230 2866 40282
rect 2918 40230 7610 40282
rect 7662 40230 7674 40282
rect 7726 40230 7738 40282
rect 7790 40230 7802 40282
rect 7854 40230 7866 40282
rect 7918 40230 12610 40282
rect 12662 40230 12674 40282
rect 12726 40230 12738 40282
rect 12790 40230 12802 40282
rect 12854 40230 12866 40282
rect 12918 40230 17610 40282
rect 17662 40230 17674 40282
rect 17726 40230 17738 40282
rect 17790 40230 17802 40282
rect 17854 40230 17866 40282
rect 17918 40230 22610 40282
rect 22662 40230 22674 40282
rect 22726 40230 22738 40282
rect 22790 40230 22802 40282
rect 22854 40230 22866 40282
rect 22918 40230 27610 40282
rect 27662 40230 27674 40282
rect 27726 40230 27738 40282
rect 27790 40230 27802 40282
rect 27854 40230 27866 40282
rect 27918 40230 32610 40282
rect 32662 40230 32674 40282
rect 32726 40230 32738 40282
rect 32790 40230 32802 40282
rect 32854 40230 32866 40282
rect 32918 40230 37610 40282
rect 37662 40230 37674 40282
rect 37726 40230 37738 40282
rect 37790 40230 37802 40282
rect 37854 40230 37866 40282
rect 37918 40230 42610 40282
rect 42662 40230 42674 40282
rect 42726 40230 42738 40282
rect 42790 40230 42802 40282
rect 42854 40230 42866 40282
rect 42918 40230 47610 40282
rect 47662 40230 47674 40282
rect 47726 40230 47738 40282
rect 47790 40230 47802 40282
rect 47854 40230 47866 40282
rect 47918 40230 52610 40282
rect 52662 40230 52674 40282
rect 52726 40230 52738 40282
rect 52790 40230 52802 40282
rect 52854 40230 52866 40282
rect 52918 40230 57610 40282
rect 57662 40230 57674 40282
rect 57726 40230 57738 40282
rect 57790 40230 57802 40282
rect 57854 40230 57866 40282
rect 57918 40230 58880 40282
rect 1104 40208 58880 40230
rect 1104 39738 58880 39760
rect 1104 39686 1950 39738
rect 2002 39686 2014 39738
rect 2066 39686 2078 39738
rect 2130 39686 2142 39738
rect 2194 39686 2206 39738
rect 2258 39686 6950 39738
rect 7002 39686 7014 39738
rect 7066 39686 7078 39738
rect 7130 39686 7142 39738
rect 7194 39686 7206 39738
rect 7258 39686 11950 39738
rect 12002 39686 12014 39738
rect 12066 39686 12078 39738
rect 12130 39686 12142 39738
rect 12194 39686 12206 39738
rect 12258 39686 16950 39738
rect 17002 39686 17014 39738
rect 17066 39686 17078 39738
rect 17130 39686 17142 39738
rect 17194 39686 17206 39738
rect 17258 39686 21950 39738
rect 22002 39686 22014 39738
rect 22066 39686 22078 39738
rect 22130 39686 22142 39738
rect 22194 39686 22206 39738
rect 22258 39686 26950 39738
rect 27002 39686 27014 39738
rect 27066 39686 27078 39738
rect 27130 39686 27142 39738
rect 27194 39686 27206 39738
rect 27258 39686 31950 39738
rect 32002 39686 32014 39738
rect 32066 39686 32078 39738
rect 32130 39686 32142 39738
rect 32194 39686 32206 39738
rect 32258 39686 36950 39738
rect 37002 39686 37014 39738
rect 37066 39686 37078 39738
rect 37130 39686 37142 39738
rect 37194 39686 37206 39738
rect 37258 39686 41950 39738
rect 42002 39686 42014 39738
rect 42066 39686 42078 39738
rect 42130 39686 42142 39738
rect 42194 39686 42206 39738
rect 42258 39686 46950 39738
rect 47002 39686 47014 39738
rect 47066 39686 47078 39738
rect 47130 39686 47142 39738
rect 47194 39686 47206 39738
rect 47258 39686 51950 39738
rect 52002 39686 52014 39738
rect 52066 39686 52078 39738
rect 52130 39686 52142 39738
rect 52194 39686 52206 39738
rect 52258 39686 56950 39738
rect 57002 39686 57014 39738
rect 57066 39686 57078 39738
rect 57130 39686 57142 39738
rect 57194 39686 57206 39738
rect 57258 39686 58880 39738
rect 1104 39664 58880 39686
rect 58526 39380 58532 39432
rect 58584 39380 58590 39432
rect 1104 39194 58880 39216
rect 1104 39142 2610 39194
rect 2662 39142 2674 39194
rect 2726 39142 2738 39194
rect 2790 39142 2802 39194
rect 2854 39142 2866 39194
rect 2918 39142 7610 39194
rect 7662 39142 7674 39194
rect 7726 39142 7738 39194
rect 7790 39142 7802 39194
rect 7854 39142 7866 39194
rect 7918 39142 12610 39194
rect 12662 39142 12674 39194
rect 12726 39142 12738 39194
rect 12790 39142 12802 39194
rect 12854 39142 12866 39194
rect 12918 39142 17610 39194
rect 17662 39142 17674 39194
rect 17726 39142 17738 39194
rect 17790 39142 17802 39194
rect 17854 39142 17866 39194
rect 17918 39142 22610 39194
rect 22662 39142 22674 39194
rect 22726 39142 22738 39194
rect 22790 39142 22802 39194
rect 22854 39142 22866 39194
rect 22918 39142 27610 39194
rect 27662 39142 27674 39194
rect 27726 39142 27738 39194
rect 27790 39142 27802 39194
rect 27854 39142 27866 39194
rect 27918 39142 32610 39194
rect 32662 39142 32674 39194
rect 32726 39142 32738 39194
rect 32790 39142 32802 39194
rect 32854 39142 32866 39194
rect 32918 39142 37610 39194
rect 37662 39142 37674 39194
rect 37726 39142 37738 39194
rect 37790 39142 37802 39194
rect 37854 39142 37866 39194
rect 37918 39142 42610 39194
rect 42662 39142 42674 39194
rect 42726 39142 42738 39194
rect 42790 39142 42802 39194
rect 42854 39142 42866 39194
rect 42918 39142 47610 39194
rect 47662 39142 47674 39194
rect 47726 39142 47738 39194
rect 47790 39142 47802 39194
rect 47854 39142 47866 39194
rect 47918 39142 52610 39194
rect 52662 39142 52674 39194
rect 52726 39142 52738 39194
rect 52790 39142 52802 39194
rect 52854 39142 52866 39194
rect 52918 39142 57610 39194
rect 57662 39142 57674 39194
rect 57726 39142 57738 39194
rect 57790 39142 57802 39194
rect 57854 39142 57866 39194
rect 57918 39142 58880 39194
rect 1104 39120 58880 39142
rect 58526 38700 58532 38752
rect 58584 38700 58590 38752
rect 1104 38650 58880 38672
rect 1104 38598 1950 38650
rect 2002 38598 2014 38650
rect 2066 38598 2078 38650
rect 2130 38598 2142 38650
rect 2194 38598 2206 38650
rect 2258 38598 6950 38650
rect 7002 38598 7014 38650
rect 7066 38598 7078 38650
rect 7130 38598 7142 38650
rect 7194 38598 7206 38650
rect 7258 38598 11950 38650
rect 12002 38598 12014 38650
rect 12066 38598 12078 38650
rect 12130 38598 12142 38650
rect 12194 38598 12206 38650
rect 12258 38598 16950 38650
rect 17002 38598 17014 38650
rect 17066 38598 17078 38650
rect 17130 38598 17142 38650
rect 17194 38598 17206 38650
rect 17258 38598 21950 38650
rect 22002 38598 22014 38650
rect 22066 38598 22078 38650
rect 22130 38598 22142 38650
rect 22194 38598 22206 38650
rect 22258 38598 26950 38650
rect 27002 38598 27014 38650
rect 27066 38598 27078 38650
rect 27130 38598 27142 38650
rect 27194 38598 27206 38650
rect 27258 38598 31950 38650
rect 32002 38598 32014 38650
rect 32066 38598 32078 38650
rect 32130 38598 32142 38650
rect 32194 38598 32206 38650
rect 32258 38598 36950 38650
rect 37002 38598 37014 38650
rect 37066 38598 37078 38650
rect 37130 38598 37142 38650
rect 37194 38598 37206 38650
rect 37258 38598 41950 38650
rect 42002 38598 42014 38650
rect 42066 38598 42078 38650
rect 42130 38598 42142 38650
rect 42194 38598 42206 38650
rect 42258 38598 46950 38650
rect 47002 38598 47014 38650
rect 47066 38598 47078 38650
rect 47130 38598 47142 38650
rect 47194 38598 47206 38650
rect 47258 38598 51950 38650
rect 52002 38598 52014 38650
rect 52066 38598 52078 38650
rect 52130 38598 52142 38650
rect 52194 38598 52206 38650
rect 52258 38598 56950 38650
rect 57002 38598 57014 38650
rect 57066 38598 57078 38650
rect 57130 38598 57142 38650
rect 57194 38598 57206 38650
rect 57258 38598 58880 38650
rect 1104 38576 58880 38598
rect 1104 38106 58880 38128
rect 1104 38054 2610 38106
rect 2662 38054 2674 38106
rect 2726 38054 2738 38106
rect 2790 38054 2802 38106
rect 2854 38054 2866 38106
rect 2918 38054 7610 38106
rect 7662 38054 7674 38106
rect 7726 38054 7738 38106
rect 7790 38054 7802 38106
rect 7854 38054 7866 38106
rect 7918 38054 12610 38106
rect 12662 38054 12674 38106
rect 12726 38054 12738 38106
rect 12790 38054 12802 38106
rect 12854 38054 12866 38106
rect 12918 38054 17610 38106
rect 17662 38054 17674 38106
rect 17726 38054 17738 38106
rect 17790 38054 17802 38106
rect 17854 38054 17866 38106
rect 17918 38054 22610 38106
rect 22662 38054 22674 38106
rect 22726 38054 22738 38106
rect 22790 38054 22802 38106
rect 22854 38054 22866 38106
rect 22918 38054 27610 38106
rect 27662 38054 27674 38106
rect 27726 38054 27738 38106
rect 27790 38054 27802 38106
rect 27854 38054 27866 38106
rect 27918 38054 32610 38106
rect 32662 38054 32674 38106
rect 32726 38054 32738 38106
rect 32790 38054 32802 38106
rect 32854 38054 32866 38106
rect 32918 38054 37610 38106
rect 37662 38054 37674 38106
rect 37726 38054 37738 38106
rect 37790 38054 37802 38106
rect 37854 38054 37866 38106
rect 37918 38054 42610 38106
rect 42662 38054 42674 38106
rect 42726 38054 42738 38106
rect 42790 38054 42802 38106
rect 42854 38054 42866 38106
rect 42918 38054 47610 38106
rect 47662 38054 47674 38106
rect 47726 38054 47738 38106
rect 47790 38054 47802 38106
rect 47854 38054 47866 38106
rect 47918 38054 52610 38106
rect 52662 38054 52674 38106
rect 52726 38054 52738 38106
rect 52790 38054 52802 38106
rect 52854 38054 52866 38106
rect 52918 38054 57610 38106
rect 57662 38054 57674 38106
rect 57726 38054 57738 38106
rect 57790 38054 57802 38106
rect 57854 38054 57866 38106
rect 57918 38054 58880 38106
rect 1104 38032 58880 38054
rect 58526 37612 58532 37664
rect 58584 37612 58590 37664
rect 1104 37562 58880 37584
rect 1104 37510 1950 37562
rect 2002 37510 2014 37562
rect 2066 37510 2078 37562
rect 2130 37510 2142 37562
rect 2194 37510 2206 37562
rect 2258 37510 6950 37562
rect 7002 37510 7014 37562
rect 7066 37510 7078 37562
rect 7130 37510 7142 37562
rect 7194 37510 7206 37562
rect 7258 37510 11950 37562
rect 12002 37510 12014 37562
rect 12066 37510 12078 37562
rect 12130 37510 12142 37562
rect 12194 37510 12206 37562
rect 12258 37510 16950 37562
rect 17002 37510 17014 37562
rect 17066 37510 17078 37562
rect 17130 37510 17142 37562
rect 17194 37510 17206 37562
rect 17258 37510 21950 37562
rect 22002 37510 22014 37562
rect 22066 37510 22078 37562
rect 22130 37510 22142 37562
rect 22194 37510 22206 37562
rect 22258 37510 26950 37562
rect 27002 37510 27014 37562
rect 27066 37510 27078 37562
rect 27130 37510 27142 37562
rect 27194 37510 27206 37562
rect 27258 37510 31950 37562
rect 32002 37510 32014 37562
rect 32066 37510 32078 37562
rect 32130 37510 32142 37562
rect 32194 37510 32206 37562
rect 32258 37510 36950 37562
rect 37002 37510 37014 37562
rect 37066 37510 37078 37562
rect 37130 37510 37142 37562
rect 37194 37510 37206 37562
rect 37258 37510 41950 37562
rect 42002 37510 42014 37562
rect 42066 37510 42078 37562
rect 42130 37510 42142 37562
rect 42194 37510 42206 37562
rect 42258 37510 46950 37562
rect 47002 37510 47014 37562
rect 47066 37510 47078 37562
rect 47130 37510 47142 37562
rect 47194 37510 47206 37562
rect 47258 37510 51950 37562
rect 52002 37510 52014 37562
rect 52066 37510 52078 37562
rect 52130 37510 52142 37562
rect 52194 37510 52206 37562
rect 52258 37510 56950 37562
rect 57002 37510 57014 37562
rect 57066 37510 57078 37562
rect 57130 37510 57142 37562
rect 57194 37510 57206 37562
rect 57258 37510 58880 37562
rect 1104 37488 58880 37510
rect 58526 37272 58532 37324
rect 58584 37272 58590 37324
rect 1104 37018 58880 37040
rect 1104 36966 2610 37018
rect 2662 36966 2674 37018
rect 2726 36966 2738 37018
rect 2790 36966 2802 37018
rect 2854 36966 2866 37018
rect 2918 36966 7610 37018
rect 7662 36966 7674 37018
rect 7726 36966 7738 37018
rect 7790 36966 7802 37018
rect 7854 36966 7866 37018
rect 7918 36966 12610 37018
rect 12662 36966 12674 37018
rect 12726 36966 12738 37018
rect 12790 36966 12802 37018
rect 12854 36966 12866 37018
rect 12918 36966 17610 37018
rect 17662 36966 17674 37018
rect 17726 36966 17738 37018
rect 17790 36966 17802 37018
rect 17854 36966 17866 37018
rect 17918 36966 22610 37018
rect 22662 36966 22674 37018
rect 22726 36966 22738 37018
rect 22790 36966 22802 37018
rect 22854 36966 22866 37018
rect 22918 36966 27610 37018
rect 27662 36966 27674 37018
rect 27726 36966 27738 37018
rect 27790 36966 27802 37018
rect 27854 36966 27866 37018
rect 27918 36966 32610 37018
rect 32662 36966 32674 37018
rect 32726 36966 32738 37018
rect 32790 36966 32802 37018
rect 32854 36966 32866 37018
rect 32918 36966 37610 37018
rect 37662 36966 37674 37018
rect 37726 36966 37738 37018
rect 37790 36966 37802 37018
rect 37854 36966 37866 37018
rect 37918 36966 42610 37018
rect 42662 36966 42674 37018
rect 42726 36966 42738 37018
rect 42790 36966 42802 37018
rect 42854 36966 42866 37018
rect 42918 36966 47610 37018
rect 47662 36966 47674 37018
rect 47726 36966 47738 37018
rect 47790 36966 47802 37018
rect 47854 36966 47866 37018
rect 47918 36966 52610 37018
rect 52662 36966 52674 37018
rect 52726 36966 52738 37018
rect 52790 36966 52802 37018
rect 52854 36966 52866 37018
rect 52918 36966 57610 37018
rect 57662 36966 57674 37018
rect 57726 36966 57738 37018
rect 57790 36966 57802 37018
rect 57854 36966 57866 37018
rect 57918 36966 58880 37018
rect 1104 36944 58880 36966
rect 1104 36474 58880 36496
rect 1104 36422 1950 36474
rect 2002 36422 2014 36474
rect 2066 36422 2078 36474
rect 2130 36422 2142 36474
rect 2194 36422 2206 36474
rect 2258 36422 6950 36474
rect 7002 36422 7014 36474
rect 7066 36422 7078 36474
rect 7130 36422 7142 36474
rect 7194 36422 7206 36474
rect 7258 36422 11950 36474
rect 12002 36422 12014 36474
rect 12066 36422 12078 36474
rect 12130 36422 12142 36474
rect 12194 36422 12206 36474
rect 12258 36422 16950 36474
rect 17002 36422 17014 36474
rect 17066 36422 17078 36474
rect 17130 36422 17142 36474
rect 17194 36422 17206 36474
rect 17258 36422 21950 36474
rect 22002 36422 22014 36474
rect 22066 36422 22078 36474
rect 22130 36422 22142 36474
rect 22194 36422 22206 36474
rect 22258 36422 26950 36474
rect 27002 36422 27014 36474
rect 27066 36422 27078 36474
rect 27130 36422 27142 36474
rect 27194 36422 27206 36474
rect 27258 36422 31950 36474
rect 32002 36422 32014 36474
rect 32066 36422 32078 36474
rect 32130 36422 32142 36474
rect 32194 36422 32206 36474
rect 32258 36422 36950 36474
rect 37002 36422 37014 36474
rect 37066 36422 37078 36474
rect 37130 36422 37142 36474
rect 37194 36422 37206 36474
rect 37258 36422 41950 36474
rect 42002 36422 42014 36474
rect 42066 36422 42078 36474
rect 42130 36422 42142 36474
rect 42194 36422 42206 36474
rect 42258 36422 46950 36474
rect 47002 36422 47014 36474
rect 47066 36422 47078 36474
rect 47130 36422 47142 36474
rect 47194 36422 47206 36474
rect 47258 36422 51950 36474
rect 52002 36422 52014 36474
rect 52066 36422 52078 36474
rect 52130 36422 52142 36474
rect 52194 36422 52206 36474
rect 52258 36422 56950 36474
rect 57002 36422 57014 36474
rect 57066 36422 57078 36474
rect 57130 36422 57142 36474
rect 57194 36422 57206 36474
rect 57258 36422 58880 36474
rect 1104 36400 58880 36422
rect 58526 36116 58532 36168
rect 58584 36116 58590 36168
rect 1104 35930 58880 35952
rect 1104 35878 2610 35930
rect 2662 35878 2674 35930
rect 2726 35878 2738 35930
rect 2790 35878 2802 35930
rect 2854 35878 2866 35930
rect 2918 35878 7610 35930
rect 7662 35878 7674 35930
rect 7726 35878 7738 35930
rect 7790 35878 7802 35930
rect 7854 35878 7866 35930
rect 7918 35878 12610 35930
rect 12662 35878 12674 35930
rect 12726 35878 12738 35930
rect 12790 35878 12802 35930
rect 12854 35878 12866 35930
rect 12918 35878 17610 35930
rect 17662 35878 17674 35930
rect 17726 35878 17738 35930
rect 17790 35878 17802 35930
rect 17854 35878 17866 35930
rect 17918 35878 22610 35930
rect 22662 35878 22674 35930
rect 22726 35878 22738 35930
rect 22790 35878 22802 35930
rect 22854 35878 22866 35930
rect 22918 35878 27610 35930
rect 27662 35878 27674 35930
rect 27726 35878 27738 35930
rect 27790 35878 27802 35930
rect 27854 35878 27866 35930
rect 27918 35878 32610 35930
rect 32662 35878 32674 35930
rect 32726 35878 32738 35930
rect 32790 35878 32802 35930
rect 32854 35878 32866 35930
rect 32918 35878 37610 35930
rect 37662 35878 37674 35930
rect 37726 35878 37738 35930
rect 37790 35878 37802 35930
rect 37854 35878 37866 35930
rect 37918 35878 42610 35930
rect 42662 35878 42674 35930
rect 42726 35878 42738 35930
rect 42790 35878 42802 35930
rect 42854 35878 42866 35930
rect 42918 35878 47610 35930
rect 47662 35878 47674 35930
rect 47726 35878 47738 35930
rect 47790 35878 47802 35930
rect 47854 35878 47866 35930
rect 47918 35878 52610 35930
rect 52662 35878 52674 35930
rect 52726 35878 52738 35930
rect 52790 35878 52802 35930
rect 52854 35878 52866 35930
rect 52918 35878 57610 35930
rect 57662 35878 57674 35930
rect 57726 35878 57738 35930
rect 57790 35878 57802 35930
rect 57854 35878 57866 35930
rect 57918 35878 58880 35930
rect 1104 35856 58880 35878
rect 58526 35436 58532 35488
rect 58584 35436 58590 35488
rect 1104 35386 58880 35408
rect 1104 35334 1950 35386
rect 2002 35334 2014 35386
rect 2066 35334 2078 35386
rect 2130 35334 2142 35386
rect 2194 35334 2206 35386
rect 2258 35334 6950 35386
rect 7002 35334 7014 35386
rect 7066 35334 7078 35386
rect 7130 35334 7142 35386
rect 7194 35334 7206 35386
rect 7258 35334 11950 35386
rect 12002 35334 12014 35386
rect 12066 35334 12078 35386
rect 12130 35334 12142 35386
rect 12194 35334 12206 35386
rect 12258 35334 16950 35386
rect 17002 35334 17014 35386
rect 17066 35334 17078 35386
rect 17130 35334 17142 35386
rect 17194 35334 17206 35386
rect 17258 35334 21950 35386
rect 22002 35334 22014 35386
rect 22066 35334 22078 35386
rect 22130 35334 22142 35386
rect 22194 35334 22206 35386
rect 22258 35334 26950 35386
rect 27002 35334 27014 35386
rect 27066 35334 27078 35386
rect 27130 35334 27142 35386
rect 27194 35334 27206 35386
rect 27258 35334 31950 35386
rect 32002 35334 32014 35386
rect 32066 35334 32078 35386
rect 32130 35334 32142 35386
rect 32194 35334 32206 35386
rect 32258 35334 36950 35386
rect 37002 35334 37014 35386
rect 37066 35334 37078 35386
rect 37130 35334 37142 35386
rect 37194 35334 37206 35386
rect 37258 35334 41950 35386
rect 42002 35334 42014 35386
rect 42066 35334 42078 35386
rect 42130 35334 42142 35386
rect 42194 35334 42206 35386
rect 42258 35334 46950 35386
rect 47002 35334 47014 35386
rect 47066 35334 47078 35386
rect 47130 35334 47142 35386
rect 47194 35334 47206 35386
rect 47258 35334 51950 35386
rect 52002 35334 52014 35386
rect 52066 35334 52078 35386
rect 52130 35334 52142 35386
rect 52194 35334 52206 35386
rect 52258 35334 56950 35386
rect 57002 35334 57014 35386
rect 57066 35334 57078 35386
rect 57130 35334 57142 35386
rect 57194 35334 57206 35386
rect 57258 35334 58880 35386
rect 1104 35312 58880 35334
rect 1104 34842 58880 34864
rect 1104 34790 2610 34842
rect 2662 34790 2674 34842
rect 2726 34790 2738 34842
rect 2790 34790 2802 34842
rect 2854 34790 2866 34842
rect 2918 34790 7610 34842
rect 7662 34790 7674 34842
rect 7726 34790 7738 34842
rect 7790 34790 7802 34842
rect 7854 34790 7866 34842
rect 7918 34790 12610 34842
rect 12662 34790 12674 34842
rect 12726 34790 12738 34842
rect 12790 34790 12802 34842
rect 12854 34790 12866 34842
rect 12918 34790 17610 34842
rect 17662 34790 17674 34842
rect 17726 34790 17738 34842
rect 17790 34790 17802 34842
rect 17854 34790 17866 34842
rect 17918 34790 22610 34842
rect 22662 34790 22674 34842
rect 22726 34790 22738 34842
rect 22790 34790 22802 34842
rect 22854 34790 22866 34842
rect 22918 34790 27610 34842
rect 27662 34790 27674 34842
rect 27726 34790 27738 34842
rect 27790 34790 27802 34842
rect 27854 34790 27866 34842
rect 27918 34790 32610 34842
rect 32662 34790 32674 34842
rect 32726 34790 32738 34842
rect 32790 34790 32802 34842
rect 32854 34790 32866 34842
rect 32918 34790 37610 34842
rect 37662 34790 37674 34842
rect 37726 34790 37738 34842
rect 37790 34790 37802 34842
rect 37854 34790 37866 34842
rect 37918 34790 42610 34842
rect 42662 34790 42674 34842
rect 42726 34790 42738 34842
rect 42790 34790 42802 34842
rect 42854 34790 42866 34842
rect 42918 34790 47610 34842
rect 47662 34790 47674 34842
rect 47726 34790 47738 34842
rect 47790 34790 47802 34842
rect 47854 34790 47866 34842
rect 47918 34790 52610 34842
rect 52662 34790 52674 34842
rect 52726 34790 52738 34842
rect 52790 34790 52802 34842
rect 52854 34790 52866 34842
rect 52918 34790 57610 34842
rect 57662 34790 57674 34842
rect 57726 34790 57738 34842
rect 57790 34790 57802 34842
rect 57854 34790 57866 34842
rect 57918 34790 58880 34842
rect 1104 34768 58880 34790
rect 58526 34348 58532 34400
rect 58584 34348 58590 34400
rect 1104 34298 58880 34320
rect 1104 34246 1950 34298
rect 2002 34246 2014 34298
rect 2066 34246 2078 34298
rect 2130 34246 2142 34298
rect 2194 34246 2206 34298
rect 2258 34246 6950 34298
rect 7002 34246 7014 34298
rect 7066 34246 7078 34298
rect 7130 34246 7142 34298
rect 7194 34246 7206 34298
rect 7258 34246 11950 34298
rect 12002 34246 12014 34298
rect 12066 34246 12078 34298
rect 12130 34246 12142 34298
rect 12194 34246 12206 34298
rect 12258 34246 16950 34298
rect 17002 34246 17014 34298
rect 17066 34246 17078 34298
rect 17130 34246 17142 34298
rect 17194 34246 17206 34298
rect 17258 34246 21950 34298
rect 22002 34246 22014 34298
rect 22066 34246 22078 34298
rect 22130 34246 22142 34298
rect 22194 34246 22206 34298
rect 22258 34246 26950 34298
rect 27002 34246 27014 34298
rect 27066 34246 27078 34298
rect 27130 34246 27142 34298
rect 27194 34246 27206 34298
rect 27258 34246 31950 34298
rect 32002 34246 32014 34298
rect 32066 34246 32078 34298
rect 32130 34246 32142 34298
rect 32194 34246 32206 34298
rect 32258 34246 36950 34298
rect 37002 34246 37014 34298
rect 37066 34246 37078 34298
rect 37130 34246 37142 34298
rect 37194 34246 37206 34298
rect 37258 34246 41950 34298
rect 42002 34246 42014 34298
rect 42066 34246 42078 34298
rect 42130 34246 42142 34298
rect 42194 34246 42206 34298
rect 42258 34246 46950 34298
rect 47002 34246 47014 34298
rect 47066 34246 47078 34298
rect 47130 34246 47142 34298
rect 47194 34246 47206 34298
rect 47258 34246 51950 34298
rect 52002 34246 52014 34298
rect 52066 34246 52078 34298
rect 52130 34246 52142 34298
rect 52194 34246 52206 34298
rect 52258 34246 56950 34298
rect 57002 34246 57014 34298
rect 57066 34246 57078 34298
rect 57130 34246 57142 34298
rect 57194 34246 57206 34298
rect 57258 34246 58880 34298
rect 1104 34224 58880 34246
rect 58526 33940 58532 33992
rect 58584 33940 58590 33992
rect 1104 33754 58880 33776
rect 1104 33702 2610 33754
rect 2662 33702 2674 33754
rect 2726 33702 2738 33754
rect 2790 33702 2802 33754
rect 2854 33702 2866 33754
rect 2918 33702 7610 33754
rect 7662 33702 7674 33754
rect 7726 33702 7738 33754
rect 7790 33702 7802 33754
rect 7854 33702 7866 33754
rect 7918 33702 12610 33754
rect 12662 33702 12674 33754
rect 12726 33702 12738 33754
rect 12790 33702 12802 33754
rect 12854 33702 12866 33754
rect 12918 33702 17610 33754
rect 17662 33702 17674 33754
rect 17726 33702 17738 33754
rect 17790 33702 17802 33754
rect 17854 33702 17866 33754
rect 17918 33702 22610 33754
rect 22662 33702 22674 33754
rect 22726 33702 22738 33754
rect 22790 33702 22802 33754
rect 22854 33702 22866 33754
rect 22918 33702 27610 33754
rect 27662 33702 27674 33754
rect 27726 33702 27738 33754
rect 27790 33702 27802 33754
rect 27854 33702 27866 33754
rect 27918 33702 32610 33754
rect 32662 33702 32674 33754
rect 32726 33702 32738 33754
rect 32790 33702 32802 33754
rect 32854 33702 32866 33754
rect 32918 33702 37610 33754
rect 37662 33702 37674 33754
rect 37726 33702 37738 33754
rect 37790 33702 37802 33754
rect 37854 33702 37866 33754
rect 37918 33702 42610 33754
rect 42662 33702 42674 33754
rect 42726 33702 42738 33754
rect 42790 33702 42802 33754
rect 42854 33702 42866 33754
rect 42918 33702 47610 33754
rect 47662 33702 47674 33754
rect 47726 33702 47738 33754
rect 47790 33702 47802 33754
rect 47854 33702 47866 33754
rect 47918 33702 52610 33754
rect 52662 33702 52674 33754
rect 52726 33702 52738 33754
rect 52790 33702 52802 33754
rect 52854 33702 52866 33754
rect 52918 33702 57610 33754
rect 57662 33702 57674 33754
rect 57726 33702 57738 33754
rect 57790 33702 57802 33754
rect 57854 33702 57866 33754
rect 57918 33702 58880 33754
rect 1104 33680 58880 33702
rect 1104 33210 58880 33232
rect 1104 33158 1950 33210
rect 2002 33158 2014 33210
rect 2066 33158 2078 33210
rect 2130 33158 2142 33210
rect 2194 33158 2206 33210
rect 2258 33158 6950 33210
rect 7002 33158 7014 33210
rect 7066 33158 7078 33210
rect 7130 33158 7142 33210
rect 7194 33158 7206 33210
rect 7258 33158 11950 33210
rect 12002 33158 12014 33210
rect 12066 33158 12078 33210
rect 12130 33158 12142 33210
rect 12194 33158 12206 33210
rect 12258 33158 16950 33210
rect 17002 33158 17014 33210
rect 17066 33158 17078 33210
rect 17130 33158 17142 33210
rect 17194 33158 17206 33210
rect 17258 33158 21950 33210
rect 22002 33158 22014 33210
rect 22066 33158 22078 33210
rect 22130 33158 22142 33210
rect 22194 33158 22206 33210
rect 22258 33158 26950 33210
rect 27002 33158 27014 33210
rect 27066 33158 27078 33210
rect 27130 33158 27142 33210
rect 27194 33158 27206 33210
rect 27258 33158 31950 33210
rect 32002 33158 32014 33210
rect 32066 33158 32078 33210
rect 32130 33158 32142 33210
rect 32194 33158 32206 33210
rect 32258 33158 36950 33210
rect 37002 33158 37014 33210
rect 37066 33158 37078 33210
rect 37130 33158 37142 33210
rect 37194 33158 37206 33210
rect 37258 33158 41950 33210
rect 42002 33158 42014 33210
rect 42066 33158 42078 33210
rect 42130 33158 42142 33210
rect 42194 33158 42206 33210
rect 42258 33158 46950 33210
rect 47002 33158 47014 33210
rect 47066 33158 47078 33210
rect 47130 33158 47142 33210
rect 47194 33158 47206 33210
rect 47258 33158 51950 33210
rect 52002 33158 52014 33210
rect 52066 33158 52078 33210
rect 52130 33158 52142 33210
rect 52194 33158 52206 33210
rect 52258 33158 56950 33210
rect 57002 33158 57014 33210
rect 57066 33158 57078 33210
rect 57130 33158 57142 33210
rect 57194 33158 57206 33210
rect 57258 33158 58880 33210
rect 1104 33136 58880 33158
rect 58526 32852 58532 32904
rect 58584 32852 58590 32904
rect 1104 32666 58880 32688
rect 1104 32614 2610 32666
rect 2662 32614 2674 32666
rect 2726 32614 2738 32666
rect 2790 32614 2802 32666
rect 2854 32614 2866 32666
rect 2918 32614 7610 32666
rect 7662 32614 7674 32666
rect 7726 32614 7738 32666
rect 7790 32614 7802 32666
rect 7854 32614 7866 32666
rect 7918 32614 12610 32666
rect 12662 32614 12674 32666
rect 12726 32614 12738 32666
rect 12790 32614 12802 32666
rect 12854 32614 12866 32666
rect 12918 32614 17610 32666
rect 17662 32614 17674 32666
rect 17726 32614 17738 32666
rect 17790 32614 17802 32666
rect 17854 32614 17866 32666
rect 17918 32614 22610 32666
rect 22662 32614 22674 32666
rect 22726 32614 22738 32666
rect 22790 32614 22802 32666
rect 22854 32614 22866 32666
rect 22918 32614 27610 32666
rect 27662 32614 27674 32666
rect 27726 32614 27738 32666
rect 27790 32614 27802 32666
rect 27854 32614 27866 32666
rect 27918 32614 32610 32666
rect 32662 32614 32674 32666
rect 32726 32614 32738 32666
rect 32790 32614 32802 32666
rect 32854 32614 32866 32666
rect 32918 32614 37610 32666
rect 37662 32614 37674 32666
rect 37726 32614 37738 32666
rect 37790 32614 37802 32666
rect 37854 32614 37866 32666
rect 37918 32614 42610 32666
rect 42662 32614 42674 32666
rect 42726 32614 42738 32666
rect 42790 32614 42802 32666
rect 42854 32614 42866 32666
rect 42918 32614 47610 32666
rect 47662 32614 47674 32666
rect 47726 32614 47738 32666
rect 47790 32614 47802 32666
rect 47854 32614 47866 32666
rect 47918 32614 52610 32666
rect 52662 32614 52674 32666
rect 52726 32614 52738 32666
rect 52790 32614 52802 32666
rect 52854 32614 52866 32666
rect 52918 32614 57610 32666
rect 57662 32614 57674 32666
rect 57726 32614 57738 32666
rect 57790 32614 57802 32666
rect 57854 32614 57866 32666
rect 57918 32614 58880 32666
rect 1104 32592 58880 32614
rect 58526 32172 58532 32224
rect 58584 32172 58590 32224
rect 1104 32122 58880 32144
rect 1104 32070 1950 32122
rect 2002 32070 2014 32122
rect 2066 32070 2078 32122
rect 2130 32070 2142 32122
rect 2194 32070 2206 32122
rect 2258 32070 6950 32122
rect 7002 32070 7014 32122
rect 7066 32070 7078 32122
rect 7130 32070 7142 32122
rect 7194 32070 7206 32122
rect 7258 32070 11950 32122
rect 12002 32070 12014 32122
rect 12066 32070 12078 32122
rect 12130 32070 12142 32122
rect 12194 32070 12206 32122
rect 12258 32070 16950 32122
rect 17002 32070 17014 32122
rect 17066 32070 17078 32122
rect 17130 32070 17142 32122
rect 17194 32070 17206 32122
rect 17258 32070 21950 32122
rect 22002 32070 22014 32122
rect 22066 32070 22078 32122
rect 22130 32070 22142 32122
rect 22194 32070 22206 32122
rect 22258 32070 26950 32122
rect 27002 32070 27014 32122
rect 27066 32070 27078 32122
rect 27130 32070 27142 32122
rect 27194 32070 27206 32122
rect 27258 32070 31950 32122
rect 32002 32070 32014 32122
rect 32066 32070 32078 32122
rect 32130 32070 32142 32122
rect 32194 32070 32206 32122
rect 32258 32070 36950 32122
rect 37002 32070 37014 32122
rect 37066 32070 37078 32122
rect 37130 32070 37142 32122
rect 37194 32070 37206 32122
rect 37258 32070 41950 32122
rect 42002 32070 42014 32122
rect 42066 32070 42078 32122
rect 42130 32070 42142 32122
rect 42194 32070 42206 32122
rect 42258 32070 46950 32122
rect 47002 32070 47014 32122
rect 47066 32070 47078 32122
rect 47130 32070 47142 32122
rect 47194 32070 47206 32122
rect 47258 32070 51950 32122
rect 52002 32070 52014 32122
rect 52066 32070 52078 32122
rect 52130 32070 52142 32122
rect 52194 32070 52206 32122
rect 52258 32070 56950 32122
rect 57002 32070 57014 32122
rect 57066 32070 57078 32122
rect 57130 32070 57142 32122
rect 57194 32070 57206 32122
rect 57258 32070 58880 32122
rect 1104 32048 58880 32070
rect 1104 31578 58880 31600
rect 1104 31526 2610 31578
rect 2662 31526 2674 31578
rect 2726 31526 2738 31578
rect 2790 31526 2802 31578
rect 2854 31526 2866 31578
rect 2918 31526 7610 31578
rect 7662 31526 7674 31578
rect 7726 31526 7738 31578
rect 7790 31526 7802 31578
rect 7854 31526 7866 31578
rect 7918 31526 12610 31578
rect 12662 31526 12674 31578
rect 12726 31526 12738 31578
rect 12790 31526 12802 31578
rect 12854 31526 12866 31578
rect 12918 31526 17610 31578
rect 17662 31526 17674 31578
rect 17726 31526 17738 31578
rect 17790 31526 17802 31578
rect 17854 31526 17866 31578
rect 17918 31526 22610 31578
rect 22662 31526 22674 31578
rect 22726 31526 22738 31578
rect 22790 31526 22802 31578
rect 22854 31526 22866 31578
rect 22918 31526 27610 31578
rect 27662 31526 27674 31578
rect 27726 31526 27738 31578
rect 27790 31526 27802 31578
rect 27854 31526 27866 31578
rect 27918 31526 32610 31578
rect 32662 31526 32674 31578
rect 32726 31526 32738 31578
rect 32790 31526 32802 31578
rect 32854 31526 32866 31578
rect 32918 31526 37610 31578
rect 37662 31526 37674 31578
rect 37726 31526 37738 31578
rect 37790 31526 37802 31578
rect 37854 31526 37866 31578
rect 37918 31526 42610 31578
rect 42662 31526 42674 31578
rect 42726 31526 42738 31578
rect 42790 31526 42802 31578
rect 42854 31526 42866 31578
rect 42918 31526 47610 31578
rect 47662 31526 47674 31578
rect 47726 31526 47738 31578
rect 47790 31526 47802 31578
rect 47854 31526 47866 31578
rect 47918 31526 52610 31578
rect 52662 31526 52674 31578
rect 52726 31526 52738 31578
rect 52790 31526 52802 31578
rect 52854 31526 52866 31578
rect 52918 31526 57610 31578
rect 57662 31526 57674 31578
rect 57726 31526 57738 31578
rect 57790 31526 57802 31578
rect 57854 31526 57866 31578
rect 57918 31526 58880 31578
rect 1104 31504 58880 31526
rect 58526 31084 58532 31136
rect 58584 31084 58590 31136
rect 1104 31034 58880 31056
rect 1104 30982 1950 31034
rect 2002 30982 2014 31034
rect 2066 30982 2078 31034
rect 2130 30982 2142 31034
rect 2194 30982 2206 31034
rect 2258 30982 6950 31034
rect 7002 30982 7014 31034
rect 7066 30982 7078 31034
rect 7130 30982 7142 31034
rect 7194 30982 7206 31034
rect 7258 30982 11950 31034
rect 12002 30982 12014 31034
rect 12066 30982 12078 31034
rect 12130 30982 12142 31034
rect 12194 30982 12206 31034
rect 12258 30982 16950 31034
rect 17002 30982 17014 31034
rect 17066 30982 17078 31034
rect 17130 30982 17142 31034
rect 17194 30982 17206 31034
rect 17258 30982 21950 31034
rect 22002 30982 22014 31034
rect 22066 30982 22078 31034
rect 22130 30982 22142 31034
rect 22194 30982 22206 31034
rect 22258 30982 26950 31034
rect 27002 30982 27014 31034
rect 27066 30982 27078 31034
rect 27130 30982 27142 31034
rect 27194 30982 27206 31034
rect 27258 30982 31950 31034
rect 32002 30982 32014 31034
rect 32066 30982 32078 31034
rect 32130 30982 32142 31034
rect 32194 30982 32206 31034
rect 32258 30982 36950 31034
rect 37002 30982 37014 31034
rect 37066 30982 37078 31034
rect 37130 30982 37142 31034
rect 37194 30982 37206 31034
rect 37258 30982 41950 31034
rect 42002 30982 42014 31034
rect 42066 30982 42078 31034
rect 42130 30982 42142 31034
rect 42194 30982 42206 31034
rect 42258 30982 46950 31034
rect 47002 30982 47014 31034
rect 47066 30982 47078 31034
rect 47130 30982 47142 31034
rect 47194 30982 47206 31034
rect 47258 30982 51950 31034
rect 52002 30982 52014 31034
rect 52066 30982 52078 31034
rect 52130 30982 52142 31034
rect 52194 30982 52206 31034
rect 52258 30982 56950 31034
rect 57002 30982 57014 31034
rect 57066 30982 57078 31034
rect 57130 30982 57142 31034
rect 57194 30982 57206 31034
rect 57258 30982 58880 31034
rect 1104 30960 58880 30982
rect 58526 30676 58532 30728
rect 58584 30676 58590 30728
rect 1104 30490 58880 30512
rect 1104 30438 2610 30490
rect 2662 30438 2674 30490
rect 2726 30438 2738 30490
rect 2790 30438 2802 30490
rect 2854 30438 2866 30490
rect 2918 30438 7610 30490
rect 7662 30438 7674 30490
rect 7726 30438 7738 30490
rect 7790 30438 7802 30490
rect 7854 30438 7866 30490
rect 7918 30438 12610 30490
rect 12662 30438 12674 30490
rect 12726 30438 12738 30490
rect 12790 30438 12802 30490
rect 12854 30438 12866 30490
rect 12918 30438 17610 30490
rect 17662 30438 17674 30490
rect 17726 30438 17738 30490
rect 17790 30438 17802 30490
rect 17854 30438 17866 30490
rect 17918 30438 22610 30490
rect 22662 30438 22674 30490
rect 22726 30438 22738 30490
rect 22790 30438 22802 30490
rect 22854 30438 22866 30490
rect 22918 30438 27610 30490
rect 27662 30438 27674 30490
rect 27726 30438 27738 30490
rect 27790 30438 27802 30490
rect 27854 30438 27866 30490
rect 27918 30438 32610 30490
rect 32662 30438 32674 30490
rect 32726 30438 32738 30490
rect 32790 30438 32802 30490
rect 32854 30438 32866 30490
rect 32918 30438 37610 30490
rect 37662 30438 37674 30490
rect 37726 30438 37738 30490
rect 37790 30438 37802 30490
rect 37854 30438 37866 30490
rect 37918 30438 42610 30490
rect 42662 30438 42674 30490
rect 42726 30438 42738 30490
rect 42790 30438 42802 30490
rect 42854 30438 42866 30490
rect 42918 30438 47610 30490
rect 47662 30438 47674 30490
rect 47726 30438 47738 30490
rect 47790 30438 47802 30490
rect 47854 30438 47866 30490
rect 47918 30438 52610 30490
rect 52662 30438 52674 30490
rect 52726 30438 52738 30490
rect 52790 30438 52802 30490
rect 52854 30438 52866 30490
rect 52918 30438 57610 30490
rect 57662 30438 57674 30490
rect 57726 30438 57738 30490
rect 57790 30438 57802 30490
rect 57854 30438 57866 30490
rect 57918 30438 58880 30490
rect 1104 30416 58880 30438
rect 1104 29946 58880 29968
rect 1104 29894 1950 29946
rect 2002 29894 2014 29946
rect 2066 29894 2078 29946
rect 2130 29894 2142 29946
rect 2194 29894 2206 29946
rect 2258 29894 6950 29946
rect 7002 29894 7014 29946
rect 7066 29894 7078 29946
rect 7130 29894 7142 29946
rect 7194 29894 7206 29946
rect 7258 29894 11950 29946
rect 12002 29894 12014 29946
rect 12066 29894 12078 29946
rect 12130 29894 12142 29946
rect 12194 29894 12206 29946
rect 12258 29894 16950 29946
rect 17002 29894 17014 29946
rect 17066 29894 17078 29946
rect 17130 29894 17142 29946
rect 17194 29894 17206 29946
rect 17258 29894 21950 29946
rect 22002 29894 22014 29946
rect 22066 29894 22078 29946
rect 22130 29894 22142 29946
rect 22194 29894 22206 29946
rect 22258 29894 26950 29946
rect 27002 29894 27014 29946
rect 27066 29894 27078 29946
rect 27130 29894 27142 29946
rect 27194 29894 27206 29946
rect 27258 29894 31950 29946
rect 32002 29894 32014 29946
rect 32066 29894 32078 29946
rect 32130 29894 32142 29946
rect 32194 29894 32206 29946
rect 32258 29894 36950 29946
rect 37002 29894 37014 29946
rect 37066 29894 37078 29946
rect 37130 29894 37142 29946
rect 37194 29894 37206 29946
rect 37258 29894 41950 29946
rect 42002 29894 42014 29946
rect 42066 29894 42078 29946
rect 42130 29894 42142 29946
rect 42194 29894 42206 29946
rect 42258 29894 46950 29946
rect 47002 29894 47014 29946
rect 47066 29894 47078 29946
rect 47130 29894 47142 29946
rect 47194 29894 47206 29946
rect 47258 29894 51950 29946
rect 52002 29894 52014 29946
rect 52066 29894 52078 29946
rect 52130 29894 52142 29946
rect 52194 29894 52206 29946
rect 52258 29894 56950 29946
rect 57002 29894 57014 29946
rect 57066 29894 57078 29946
rect 57130 29894 57142 29946
rect 57194 29894 57206 29946
rect 57258 29894 58880 29946
rect 1104 29872 58880 29894
rect 58526 29588 58532 29640
rect 58584 29588 58590 29640
rect 1104 29402 58880 29424
rect 1104 29350 2610 29402
rect 2662 29350 2674 29402
rect 2726 29350 2738 29402
rect 2790 29350 2802 29402
rect 2854 29350 2866 29402
rect 2918 29350 7610 29402
rect 7662 29350 7674 29402
rect 7726 29350 7738 29402
rect 7790 29350 7802 29402
rect 7854 29350 7866 29402
rect 7918 29350 12610 29402
rect 12662 29350 12674 29402
rect 12726 29350 12738 29402
rect 12790 29350 12802 29402
rect 12854 29350 12866 29402
rect 12918 29350 17610 29402
rect 17662 29350 17674 29402
rect 17726 29350 17738 29402
rect 17790 29350 17802 29402
rect 17854 29350 17866 29402
rect 17918 29350 22610 29402
rect 22662 29350 22674 29402
rect 22726 29350 22738 29402
rect 22790 29350 22802 29402
rect 22854 29350 22866 29402
rect 22918 29350 27610 29402
rect 27662 29350 27674 29402
rect 27726 29350 27738 29402
rect 27790 29350 27802 29402
rect 27854 29350 27866 29402
rect 27918 29350 32610 29402
rect 32662 29350 32674 29402
rect 32726 29350 32738 29402
rect 32790 29350 32802 29402
rect 32854 29350 32866 29402
rect 32918 29350 37610 29402
rect 37662 29350 37674 29402
rect 37726 29350 37738 29402
rect 37790 29350 37802 29402
rect 37854 29350 37866 29402
rect 37918 29350 42610 29402
rect 42662 29350 42674 29402
rect 42726 29350 42738 29402
rect 42790 29350 42802 29402
rect 42854 29350 42866 29402
rect 42918 29350 47610 29402
rect 47662 29350 47674 29402
rect 47726 29350 47738 29402
rect 47790 29350 47802 29402
rect 47854 29350 47866 29402
rect 47918 29350 52610 29402
rect 52662 29350 52674 29402
rect 52726 29350 52738 29402
rect 52790 29350 52802 29402
rect 52854 29350 52866 29402
rect 52918 29350 57610 29402
rect 57662 29350 57674 29402
rect 57726 29350 57738 29402
rect 57790 29350 57802 29402
rect 57854 29350 57866 29402
rect 57918 29350 58880 29402
rect 1104 29328 58880 29350
rect 58526 28976 58532 29028
rect 58584 28976 58590 29028
rect 1104 28858 58880 28880
rect 1104 28806 1950 28858
rect 2002 28806 2014 28858
rect 2066 28806 2078 28858
rect 2130 28806 2142 28858
rect 2194 28806 2206 28858
rect 2258 28806 6950 28858
rect 7002 28806 7014 28858
rect 7066 28806 7078 28858
rect 7130 28806 7142 28858
rect 7194 28806 7206 28858
rect 7258 28806 11950 28858
rect 12002 28806 12014 28858
rect 12066 28806 12078 28858
rect 12130 28806 12142 28858
rect 12194 28806 12206 28858
rect 12258 28806 16950 28858
rect 17002 28806 17014 28858
rect 17066 28806 17078 28858
rect 17130 28806 17142 28858
rect 17194 28806 17206 28858
rect 17258 28806 21950 28858
rect 22002 28806 22014 28858
rect 22066 28806 22078 28858
rect 22130 28806 22142 28858
rect 22194 28806 22206 28858
rect 22258 28806 26950 28858
rect 27002 28806 27014 28858
rect 27066 28806 27078 28858
rect 27130 28806 27142 28858
rect 27194 28806 27206 28858
rect 27258 28806 31950 28858
rect 32002 28806 32014 28858
rect 32066 28806 32078 28858
rect 32130 28806 32142 28858
rect 32194 28806 32206 28858
rect 32258 28806 36950 28858
rect 37002 28806 37014 28858
rect 37066 28806 37078 28858
rect 37130 28806 37142 28858
rect 37194 28806 37206 28858
rect 37258 28806 41950 28858
rect 42002 28806 42014 28858
rect 42066 28806 42078 28858
rect 42130 28806 42142 28858
rect 42194 28806 42206 28858
rect 42258 28806 46950 28858
rect 47002 28806 47014 28858
rect 47066 28806 47078 28858
rect 47130 28806 47142 28858
rect 47194 28806 47206 28858
rect 47258 28806 51950 28858
rect 52002 28806 52014 28858
rect 52066 28806 52078 28858
rect 52130 28806 52142 28858
rect 52194 28806 52206 28858
rect 52258 28806 56950 28858
rect 57002 28806 57014 28858
rect 57066 28806 57078 28858
rect 57130 28806 57142 28858
rect 57194 28806 57206 28858
rect 57258 28806 58880 28858
rect 1104 28784 58880 28806
rect 1104 28314 58880 28336
rect 1104 28262 2610 28314
rect 2662 28262 2674 28314
rect 2726 28262 2738 28314
rect 2790 28262 2802 28314
rect 2854 28262 2866 28314
rect 2918 28262 7610 28314
rect 7662 28262 7674 28314
rect 7726 28262 7738 28314
rect 7790 28262 7802 28314
rect 7854 28262 7866 28314
rect 7918 28262 12610 28314
rect 12662 28262 12674 28314
rect 12726 28262 12738 28314
rect 12790 28262 12802 28314
rect 12854 28262 12866 28314
rect 12918 28262 17610 28314
rect 17662 28262 17674 28314
rect 17726 28262 17738 28314
rect 17790 28262 17802 28314
rect 17854 28262 17866 28314
rect 17918 28262 22610 28314
rect 22662 28262 22674 28314
rect 22726 28262 22738 28314
rect 22790 28262 22802 28314
rect 22854 28262 22866 28314
rect 22918 28262 27610 28314
rect 27662 28262 27674 28314
rect 27726 28262 27738 28314
rect 27790 28262 27802 28314
rect 27854 28262 27866 28314
rect 27918 28262 32610 28314
rect 32662 28262 32674 28314
rect 32726 28262 32738 28314
rect 32790 28262 32802 28314
rect 32854 28262 32866 28314
rect 32918 28262 37610 28314
rect 37662 28262 37674 28314
rect 37726 28262 37738 28314
rect 37790 28262 37802 28314
rect 37854 28262 37866 28314
rect 37918 28262 42610 28314
rect 42662 28262 42674 28314
rect 42726 28262 42738 28314
rect 42790 28262 42802 28314
rect 42854 28262 42866 28314
rect 42918 28262 47610 28314
rect 47662 28262 47674 28314
rect 47726 28262 47738 28314
rect 47790 28262 47802 28314
rect 47854 28262 47866 28314
rect 47918 28262 52610 28314
rect 52662 28262 52674 28314
rect 52726 28262 52738 28314
rect 52790 28262 52802 28314
rect 52854 28262 52866 28314
rect 52918 28262 57610 28314
rect 57662 28262 57674 28314
rect 57726 28262 57738 28314
rect 57790 28262 57802 28314
rect 57854 28262 57866 28314
rect 57918 28262 58880 28314
rect 1104 28240 58880 28262
rect 58526 27820 58532 27872
rect 58584 27820 58590 27872
rect 1104 27770 58880 27792
rect 1104 27718 1950 27770
rect 2002 27718 2014 27770
rect 2066 27718 2078 27770
rect 2130 27718 2142 27770
rect 2194 27718 2206 27770
rect 2258 27718 6950 27770
rect 7002 27718 7014 27770
rect 7066 27718 7078 27770
rect 7130 27718 7142 27770
rect 7194 27718 7206 27770
rect 7258 27718 11950 27770
rect 12002 27718 12014 27770
rect 12066 27718 12078 27770
rect 12130 27718 12142 27770
rect 12194 27718 12206 27770
rect 12258 27718 16950 27770
rect 17002 27718 17014 27770
rect 17066 27718 17078 27770
rect 17130 27718 17142 27770
rect 17194 27718 17206 27770
rect 17258 27718 21950 27770
rect 22002 27718 22014 27770
rect 22066 27718 22078 27770
rect 22130 27718 22142 27770
rect 22194 27718 22206 27770
rect 22258 27718 26950 27770
rect 27002 27718 27014 27770
rect 27066 27718 27078 27770
rect 27130 27718 27142 27770
rect 27194 27718 27206 27770
rect 27258 27718 31950 27770
rect 32002 27718 32014 27770
rect 32066 27718 32078 27770
rect 32130 27718 32142 27770
rect 32194 27718 32206 27770
rect 32258 27718 36950 27770
rect 37002 27718 37014 27770
rect 37066 27718 37078 27770
rect 37130 27718 37142 27770
rect 37194 27718 37206 27770
rect 37258 27718 41950 27770
rect 42002 27718 42014 27770
rect 42066 27718 42078 27770
rect 42130 27718 42142 27770
rect 42194 27718 42206 27770
rect 42258 27718 46950 27770
rect 47002 27718 47014 27770
rect 47066 27718 47078 27770
rect 47130 27718 47142 27770
rect 47194 27718 47206 27770
rect 47258 27718 51950 27770
rect 52002 27718 52014 27770
rect 52066 27718 52078 27770
rect 52130 27718 52142 27770
rect 52194 27718 52206 27770
rect 52258 27718 56950 27770
rect 57002 27718 57014 27770
rect 57066 27718 57078 27770
rect 57130 27718 57142 27770
rect 57194 27718 57206 27770
rect 57258 27718 58880 27770
rect 1104 27696 58880 27718
rect 58526 27412 58532 27464
rect 58584 27412 58590 27464
rect 1104 27226 58880 27248
rect 1104 27174 2610 27226
rect 2662 27174 2674 27226
rect 2726 27174 2738 27226
rect 2790 27174 2802 27226
rect 2854 27174 2866 27226
rect 2918 27174 7610 27226
rect 7662 27174 7674 27226
rect 7726 27174 7738 27226
rect 7790 27174 7802 27226
rect 7854 27174 7866 27226
rect 7918 27174 12610 27226
rect 12662 27174 12674 27226
rect 12726 27174 12738 27226
rect 12790 27174 12802 27226
rect 12854 27174 12866 27226
rect 12918 27174 17610 27226
rect 17662 27174 17674 27226
rect 17726 27174 17738 27226
rect 17790 27174 17802 27226
rect 17854 27174 17866 27226
rect 17918 27174 22610 27226
rect 22662 27174 22674 27226
rect 22726 27174 22738 27226
rect 22790 27174 22802 27226
rect 22854 27174 22866 27226
rect 22918 27174 27610 27226
rect 27662 27174 27674 27226
rect 27726 27174 27738 27226
rect 27790 27174 27802 27226
rect 27854 27174 27866 27226
rect 27918 27174 32610 27226
rect 32662 27174 32674 27226
rect 32726 27174 32738 27226
rect 32790 27174 32802 27226
rect 32854 27174 32866 27226
rect 32918 27174 37610 27226
rect 37662 27174 37674 27226
rect 37726 27174 37738 27226
rect 37790 27174 37802 27226
rect 37854 27174 37866 27226
rect 37918 27174 42610 27226
rect 42662 27174 42674 27226
rect 42726 27174 42738 27226
rect 42790 27174 42802 27226
rect 42854 27174 42866 27226
rect 42918 27174 47610 27226
rect 47662 27174 47674 27226
rect 47726 27174 47738 27226
rect 47790 27174 47802 27226
rect 47854 27174 47866 27226
rect 47918 27174 52610 27226
rect 52662 27174 52674 27226
rect 52726 27174 52738 27226
rect 52790 27174 52802 27226
rect 52854 27174 52866 27226
rect 52918 27174 57610 27226
rect 57662 27174 57674 27226
rect 57726 27174 57738 27226
rect 57790 27174 57802 27226
rect 57854 27174 57866 27226
rect 57918 27174 58880 27226
rect 1104 27152 58880 27174
rect 1104 26682 58880 26704
rect 1104 26630 1950 26682
rect 2002 26630 2014 26682
rect 2066 26630 2078 26682
rect 2130 26630 2142 26682
rect 2194 26630 2206 26682
rect 2258 26630 6950 26682
rect 7002 26630 7014 26682
rect 7066 26630 7078 26682
rect 7130 26630 7142 26682
rect 7194 26630 7206 26682
rect 7258 26630 11950 26682
rect 12002 26630 12014 26682
rect 12066 26630 12078 26682
rect 12130 26630 12142 26682
rect 12194 26630 12206 26682
rect 12258 26630 16950 26682
rect 17002 26630 17014 26682
rect 17066 26630 17078 26682
rect 17130 26630 17142 26682
rect 17194 26630 17206 26682
rect 17258 26630 21950 26682
rect 22002 26630 22014 26682
rect 22066 26630 22078 26682
rect 22130 26630 22142 26682
rect 22194 26630 22206 26682
rect 22258 26630 26950 26682
rect 27002 26630 27014 26682
rect 27066 26630 27078 26682
rect 27130 26630 27142 26682
rect 27194 26630 27206 26682
rect 27258 26630 31950 26682
rect 32002 26630 32014 26682
rect 32066 26630 32078 26682
rect 32130 26630 32142 26682
rect 32194 26630 32206 26682
rect 32258 26630 36950 26682
rect 37002 26630 37014 26682
rect 37066 26630 37078 26682
rect 37130 26630 37142 26682
rect 37194 26630 37206 26682
rect 37258 26630 41950 26682
rect 42002 26630 42014 26682
rect 42066 26630 42078 26682
rect 42130 26630 42142 26682
rect 42194 26630 42206 26682
rect 42258 26630 46950 26682
rect 47002 26630 47014 26682
rect 47066 26630 47078 26682
rect 47130 26630 47142 26682
rect 47194 26630 47206 26682
rect 47258 26630 51950 26682
rect 52002 26630 52014 26682
rect 52066 26630 52078 26682
rect 52130 26630 52142 26682
rect 52194 26630 52206 26682
rect 52258 26630 56950 26682
rect 57002 26630 57014 26682
rect 57066 26630 57078 26682
rect 57130 26630 57142 26682
rect 57194 26630 57206 26682
rect 57258 26630 58880 26682
rect 1104 26608 58880 26630
rect 58342 26324 58348 26376
rect 58400 26364 58406 26376
rect 58529 26367 58587 26373
rect 58529 26364 58541 26367
rect 58400 26336 58541 26364
rect 58400 26324 58406 26336
rect 58529 26333 58541 26336
rect 58575 26333 58587 26367
rect 58529 26327 58587 26333
rect 1104 26138 58880 26160
rect 1104 26086 2610 26138
rect 2662 26086 2674 26138
rect 2726 26086 2738 26138
rect 2790 26086 2802 26138
rect 2854 26086 2866 26138
rect 2918 26086 7610 26138
rect 7662 26086 7674 26138
rect 7726 26086 7738 26138
rect 7790 26086 7802 26138
rect 7854 26086 7866 26138
rect 7918 26086 12610 26138
rect 12662 26086 12674 26138
rect 12726 26086 12738 26138
rect 12790 26086 12802 26138
rect 12854 26086 12866 26138
rect 12918 26086 17610 26138
rect 17662 26086 17674 26138
rect 17726 26086 17738 26138
rect 17790 26086 17802 26138
rect 17854 26086 17866 26138
rect 17918 26086 22610 26138
rect 22662 26086 22674 26138
rect 22726 26086 22738 26138
rect 22790 26086 22802 26138
rect 22854 26086 22866 26138
rect 22918 26086 27610 26138
rect 27662 26086 27674 26138
rect 27726 26086 27738 26138
rect 27790 26086 27802 26138
rect 27854 26086 27866 26138
rect 27918 26086 32610 26138
rect 32662 26086 32674 26138
rect 32726 26086 32738 26138
rect 32790 26086 32802 26138
rect 32854 26086 32866 26138
rect 32918 26086 37610 26138
rect 37662 26086 37674 26138
rect 37726 26086 37738 26138
rect 37790 26086 37802 26138
rect 37854 26086 37866 26138
rect 37918 26086 42610 26138
rect 42662 26086 42674 26138
rect 42726 26086 42738 26138
rect 42790 26086 42802 26138
rect 42854 26086 42866 26138
rect 42918 26086 47610 26138
rect 47662 26086 47674 26138
rect 47726 26086 47738 26138
rect 47790 26086 47802 26138
rect 47854 26086 47866 26138
rect 47918 26086 52610 26138
rect 52662 26086 52674 26138
rect 52726 26086 52738 26138
rect 52790 26086 52802 26138
rect 52854 26086 52866 26138
rect 52918 26086 57610 26138
rect 57662 26086 57674 26138
rect 57726 26086 57738 26138
rect 57790 26086 57802 26138
rect 57854 26086 57866 26138
rect 57918 26086 58880 26138
rect 1104 26064 58880 26086
rect 58526 25644 58532 25696
rect 58584 25644 58590 25696
rect 1104 25594 58880 25616
rect 1104 25542 1950 25594
rect 2002 25542 2014 25594
rect 2066 25542 2078 25594
rect 2130 25542 2142 25594
rect 2194 25542 2206 25594
rect 2258 25542 6950 25594
rect 7002 25542 7014 25594
rect 7066 25542 7078 25594
rect 7130 25542 7142 25594
rect 7194 25542 7206 25594
rect 7258 25542 11950 25594
rect 12002 25542 12014 25594
rect 12066 25542 12078 25594
rect 12130 25542 12142 25594
rect 12194 25542 12206 25594
rect 12258 25542 16950 25594
rect 17002 25542 17014 25594
rect 17066 25542 17078 25594
rect 17130 25542 17142 25594
rect 17194 25542 17206 25594
rect 17258 25542 21950 25594
rect 22002 25542 22014 25594
rect 22066 25542 22078 25594
rect 22130 25542 22142 25594
rect 22194 25542 22206 25594
rect 22258 25542 26950 25594
rect 27002 25542 27014 25594
rect 27066 25542 27078 25594
rect 27130 25542 27142 25594
rect 27194 25542 27206 25594
rect 27258 25542 31950 25594
rect 32002 25542 32014 25594
rect 32066 25542 32078 25594
rect 32130 25542 32142 25594
rect 32194 25542 32206 25594
rect 32258 25542 36950 25594
rect 37002 25542 37014 25594
rect 37066 25542 37078 25594
rect 37130 25542 37142 25594
rect 37194 25542 37206 25594
rect 37258 25542 41950 25594
rect 42002 25542 42014 25594
rect 42066 25542 42078 25594
rect 42130 25542 42142 25594
rect 42194 25542 42206 25594
rect 42258 25542 46950 25594
rect 47002 25542 47014 25594
rect 47066 25542 47078 25594
rect 47130 25542 47142 25594
rect 47194 25542 47206 25594
rect 47258 25542 51950 25594
rect 52002 25542 52014 25594
rect 52066 25542 52078 25594
rect 52130 25542 52142 25594
rect 52194 25542 52206 25594
rect 52258 25542 56950 25594
rect 57002 25542 57014 25594
rect 57066 25542 57078 25594
rect 57130 25542 57142 25594
rect 57194 25542 57206 25594
rect 57258 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 58880 25072
rect 1104 24998 2610 25050
rect 2662 24998 2674 25050
rect 2726 24998 2738 25050
rect 2790 24998 2802 25050
rect 2854 24998 2866 25050
rect 2918 24998 7610 25050
rect 7662 24998 7674 25050
rect 7726 24998 7738 25050
rect 7790 24998 7802 25050
rect 7854 24998 7866 25050
rect 7918 24998 12610 25050
rect 12662 24998 12674 25050
rect 12726 24998 12738 25050
rect 12790 24998 12802 25050
rect 12854 24998 12866 25050
rect 12918 24998 17610 25050
rect 17662 24998 17674 25050
rect 17726 24998 17738 25050
rect 17790 24998 17802 25050
rect 17854 24998 17866 25050
rect 17918 24998 22610 25050
rect 22662 24998 22674 25050
rect 22726 24998 22738 25050
rect 22790 24998 22802 25050
rect 22854 24998 22866 25050
rect 22918 24998 27610 25050
rect 27662 24998 27674 25050
rect 27726 24998 27738 25050
rect 27790 24998 27802 25050
rect 27854 24998 27866 25050
rect 27918 24998 32610 25050
rect 32662 24998 32674 25050
rect 32726 24998 32738 25050
rect 32790 24998 32802 25050
rect 32854 24998 32866 25050
rect 32918 24998 37610 25050
rect 37662 24998 37674 25050
rect 37726 24998 37738 25050
rect 37790 24998 37802 25050
rect 37854 24998 37866 25050
rect 37918 24998 42610 25050
rect 42662 24998 42674 25050
rect 42726 24998 42738 25050
rect 42790 24998 42802 25050
rect 42854 24998 42866 25050
rect 42918 24998 47610 25050
rect 47662 24998 47674 25050
rect 47726 24998 47738 25050
rect 47790 24998 47802 25050
rect 47854 24998 47866 25050
rect 47918 24998 52610 25050
rect 52662 24998 52674 25050
rect 52726 24998 52738 25050
rect 52790 24998 52802 25050
rect 52854 24998 52866 25050
rect 52918 24998 57610 25050
rect 57662 24998 57674 25050
rect 57726 24998 57738 25050
rect 57790 24998 57802 25050
rect 57854 24998 57866 25050
rect 57918 24998 58880 25050
rect 1104 24976 58880 24998
rect 58526 24556 58532 24608
rect 58584 24556 58590 24608
rect 1104 24506 58880 24528
rect 1104 24454 1950 24506
rect 2002 24454 2014 24506
rect 2066 24454 2078 24506
rect 2130 24454 2142 24506
rect 2194 24454 2206 24506
rect 2258 24454 6950 24506
rect 7002 24454 7014 24506
rect 7066 24454 7078 24506
rect 7130 24454 7142 24506
rect 7194 24454 7206 24506
rect 7258 24454 11950 24506
rect 12002 24454 12014 24506
rect 12066 24454 12078 24506
rect 12130 24454 12142 24506
rect 12194 24454 12206 24506
rect 12258 24454 16950 24506
rect 17002 24454 17014 24506
rect 17066 24454 17078 24506
rect 17130 24454 17142 24506
rect 17194 24454 17206 24506
rect 17258 24454 21950 24506
rect 22002 24454 22014 24506
rect 22066 24454 22078 24506
rect 22130 24454 22142 24506
rect 22194 24454 22206 24506
rect 22258 24454 26950 24506
rect 27002 24454 27014 24506
rect 27066 24454 27078 24506
rect 27130 24454 27142 24506
rect 27194 24454 27206 24506
rect 27258 24454 31950 24506
rect 32002 24454 32014 24506
rect 32066 24454 32078 24506
rect 32130 24454 32142 24506
rect 32194 24454 32206 24506
rect 32258 24454 36950 24506
rect 37002 24454 37014 24506
rect 37066 24454 37078 24506
rect 37130 24454 37142 24506
rect 37194 24454 37206 24506
rect 37258 24454 41950 24506
rect 42002 24454 42014 24506
rect 42066 24454 42078 24506
rect 42130 24454 42142 24506
rect 42194 24454 42206 24506
rect 42258 24454 46950 24506
rect 47002 24454 47014 24506
rect 47066 24454 47078 24506
rect 47130 24454 47142 24506
rect 47194 24454 47206 24506
rect 47258 24454 51950 24506
rect 52002 24454 52014 24506
rect 52066 24454 52078 24506
rect 52130 24454 52142 24506
rect 52194 24454 52206 24506
rect 52258 24454 56950 24506
rect 57002 24454 57014 24506
rect 57066 24454 57078 24506
rect 57130 24454 57142 24506
rect 57194 24454 57206 24506
rect 57258 24454 58880 24506
rect 1104 24432 58880 24454
rect 58526 24148 58532 24200
rect 58584 24148 58590 24200
rect 1104 23962 58880 23984
rect 1104 23910 2610 23962
rect 2662 23910 2674 23962
rect 2726 23910 2738 23962
rect 2790 23910 2802 23962
rect 2854 23910 2866 23962
rect 2918 23910 7610 23962
rect 7662 23910 7674 23962
rect 7726 23910 7738 23962
rect 7790 23910 7802 23962
rect 7854 23910 7866 23962
rect 7918 23910 12610 23962
rect 12662 23910 12674 23962
rect 12726 23910 12738 23962
rect 12790 23910 12802 23962
rect 12854 23910 12866 23962
rect 12918 23910 17610 23962
rect 17662 23910 17674 23962
rect 17726 23910 17738 23962
rect 17790 23910 17802 23962
rect 17854 23910 17866 23962
rect 17918 23910 22610 23962
rect 22662 23910 22674 23962
rect 22726 23910 22738 23962
rect 22790 23910 22802 23962
rect 22854 23910 22866 23962
rect 22918 23910 27610 23962
rect 27662 23910 27674 23962
rect 27726 23910 27738 23962
rect 27790 23910 27802 23962
rect 27854 23910 27866 23962
rect 27918 23910 32610 23962
rect 32662 23910 32674 23962
rect 32726 23910 32738 23962
rect 32790 23910 32802 23962
rect 32854 23910 32866 23962
rect 32918 23910 37610 23962
rect 37662 23910 37674 23962
rect 37726 23910 37738 23962
rect 37790 23910 37802 23962
rect 37854 23910 37866 23962
rect 37918 23910 42610 23962
rect 42662 23910 42674 23962
rect 42726 23910 42738 23962
rect 42790 23910 42802 23962
rect 42854 23910 42866 23962
rect 42918 23910 47610 23962
rect 47662 23910 47674 23962
rect 47726 23910 47738 23962
rect 47790 23910 47802 23962
rect 47854 23910 47866 23962
rect 47918 23910 52610 23962
rect 52662 23910 52674 23962
rect 52726 23910 52738 23962
rect 52790 23910 52802 23962
rect 52854 23910 52866 23962
rect 52918 23910 57610 23962
rect 57662 23910 57674 23962
rect 57726 23910 57738 23962
rect 57790 23910 57802 23962
rect 57854 23910 57866 23962
rect 57918 23910 58880 23962
rect 1104 23888 58880 23910
rect 1104 23418 58880 23440
rect 1104 23366 1950 23418
rect 2002 23366 2014 23418
rect 2066 23366 2078 23418
rect 2130 23366 2142 23418
rect 2194 23366 2206 23418
rect 2258 23366 6950 23418
rect 7002 23366 7014 23418
rect 7066 23366 7078 23418
rect 7130 23366 7142 23418
rect 7194 23366 7206 23418
rect 7258 23366 11950 23418
rect 12002 23366 12014 23418
rect 12066 23366 12078 23418
rect 12130 23366 12142 23418
rect 12194 23366 12206 23418
rect 12258 23366 16950 23418
rect 17002 23366 17014 23418
rect 17066 23366 17078 23418
rect 17130 23366 17142 23418
rect 17194 23366 17206 23418
rect 17258 23366 21950 23418
rect 22002 23366 22014 23418
rect 22066 23366 22078 23418
rect 22130 23366 22142 23418
rect 22194 23366 22206 23418
rect 22258 23366 26950 23418
rect 27002 23366 27014 23418
rect 27066 23366 27078 23418
rect 27130 23366 27142 23418
rect 27194 23366 27206 23418
rect 27258 23366 31950 23418
rect 32002 23366 32014 23418
rect 32066 23366 32078 23418
rect 32130 23366 32142 23418
rect 32194 23366 32206 23418
rect 32258 23366 36950 23418
rect 37002 23366 37014 23418
rect 37066 23366 37078 23418
rect 37130 23366 37142 23418
rect 37194 23366 37206 23418
rect 37258 23366 41950 23418
rect 42002 23366 42014 23418
rect 42066 23366 42078 23418
rect 42130 23366 42142 23418
rect 42194 23366 42206 23418
rect 42258 23366 46950 23418
rect 47002 23366 47014 23418
rect 47066 23366 47078 23418
rect 47130 23366 47142 23418
rect 47194 23366 47206 23418
rect 47258 23366 51950 23418
rect 52002 23366 52014 23418
rect 52066 23366 52078 23418
rect 52130 23366 52142 23418
rect 52194 23366 52206 23418
rect 52258 23366 56950 23418
rect 57002 23366 57014 23418
rect 57066 23366 57078 23418
rect 57130 23366 57142 23418
rect 57194 23366 57206 23418
rect 57258 23366 58880 23418
rect 1104 23344 58880 23366
rect 58526 23060 58532 23112
rect 58584 23060 58590 23112
rect 1104 22874 58880 22896
rect 1104 22822 2610 22874
rect 2662 22822 2674 22874
rect 2726 22822 2738 22874
rect 2790 22822 2802 22874
rect 2854 22822 2866 22874
rect 2918 22822 7610 22874
rect 7662 22822 7674 22874
rect 7726 22822 7738 22874
rect 7790 22822 7802 22874
rect 7854 22822 7866 22874
rect 7918 22822 12610 22874
rect 12662 22822 12674 22874
rect 12726 22822 12738 22874
rect 12790 22822 12802 22874
rect 12854 22822 12866 22874
rect 12918 22822 17610 22874
rect 17662 22822 17674 22874
rect 17726 22822 17738 22874
rect 17790 22822 17802 22874
rect 17854 22822 17866 22874
rect 17918 22822 22610 22874
rect 22662 22822 22674 22874
rect 22726 22822 22738 22874
rect 22790 22822 22802 22874
rect 22854 22822 22866 22874
rect 22918 22822 27610 22874
rect 27662 22822 27674 22874
rect 27726 22822 27738 22874
rect 27790 22822 27802 22874
rect 27854 22822 27866 22874
rect 27918 22822 32610 22874
rect 32662 22822 32674 22874
rect 32726 22822 32738 22874
rect 32790 22822 32802 22874
rect 32854 22822 32866 22874
rect 32918 22822 37610 22874
rect 37662 22822 37674 22874
rect 37726 22822 37738 22874
rect 37790 22822 37802 22874
rect 37854 22822 37866 22874
rect 37918 22822 42610 22874
rect 42662 22822 42674 22874
rect 42726 22822 42738 22874
rect 42790 22822 42802 22874
rect 42854 22822 42866 22874
rect 42918 22822 47610 22874
rect 47662 22822 47674 22874
rect 47726 22822 47738 22874
rect 47790 22822 47802 22874
rect 47854 22822 47866 22874
rect 47918 22822 52610 22874
rect 52662 22822 52674 22874
rect 52726 22822 52738 22874
rect 52790 22822 52802 22874
rect 52854 22822 52866 22874
rect 52918 22822 57610 22874
rect 57662 22822 57674 22874
rect 57726 22822 57738 22874
rect 57790 22822 57802 22874
rect 57854 22822 57866 22874
rect 57918 22822 58880 22874
rect 1104 22800 58880 22822
rect 58526 22380 58532 22432
rect 58584 22380 58590 22432
rect 1104 22330 58880 22352
rect 1104 22278 1950 22330
rect 2002 22278 2014 22330
rect 2066 22278 2078 22330
rect 2130 22278 2142 22330
rect 2194 22278 2206 22330
rect 2258 22278 6950 22330
rect 7002 22278 7014 22330
rect 7066 22278 7078 22330
rect 7130 22278 7142 22330
rect 7194 22278 7206 22330
rect 7258 22278 11950 22330
rect 12002 22278 12014 22330
rect 12066 22278 12078 22330
rect 12130 22278 12142 22330
rect 12194 22278 12206 22330
rect 12258 22278 16950 22330
rect 17002 22278 17014 22330
rect 17066 22278 17078 22330
rect 17130 22278 17142 22330
rect 17194 22278 17206 22330
rect 17258 22278 21950 22330
rect 22002 22278 22014 22330
rect 22066 22278 22078 22330
rect 22130 22278 22142 22330
rect 22194 22278 22206 22330
rect 22258 22278 26950 22330
rect 27002 22278 27014 22330
rect 27066 22278 27078 22330
rect 27130 22278 27142 22330
rect 27194 22278 27206 22330
rect 27258 22278 31950 22330
rect 32002 22278 32014 22330
rect 32066 22278 32078 22330
rect 32130 22278 32142 22330
rect 32194 22278 32206 22330
rect 32258 22278 36950 22330
rect 37002 22278 37014 22330
rect 37066 22278 37078 22330
rect 37130 22278 37142 22330
rect 37194 22278 37206 22330
rect 37258 22278 41950 22330
rect 42002 22278 42014 22330
rect 42066 22278 42078 22330
rect 42130 22278 42142 22330
rect 42194 22278 42206 22330
rect 42258 22278 46950 22330
rect 47002 22278 47014 22330
rect 47066 22278 47078 22330
rect 47130 22278 47142 22330
rect 47194 22278 47206 22330
rect 47258 22278 51950 22330
rect 52002 22278 52014 22330
rect 52066 22278 52078 22330
rect 52130 22278 52142 22330
rect 52194 22278 52206 22330
rect 52258 22278 56950 22330
rect 57002 22278 57014 22330
rect 57066 22278 57078 22330
rect 57130 22278 57142 22330
rect 57194 22278 57206 22330
rect 57258 22278 58880 22330
rect 1104 22256 58880 22278
rect 1104 21786 58880 21808
rect 1104 21734 2610 21786
rect 2662 21734 2674 21786
rect 2726 21734 2738 21786
rect 2790 21734 2802 21786
rect 2854 21734 2866 21786
rect 2918 21734 7610 21786
rect 7662 21734 7674 21786
rect 7726 21734 7738 21786
rect 7790 21734 7802 21786
rect 7854 21734 7866 21786
rect 7918 21734 12610 21786
rect 12662 21734 12674 21786
rect 12726 21734 12738 21786
rect 12790 21734 12802 21786
rect 12854 21734 12866 21786
rect 12918 21734 17610 21786
rect 17662 21734 17674 21786
rect 17726 21734 17738 21786
rect 17790 21734 17802 21786
rect 17854 21734 17866 21786
rect 17918 21734 22610 21786
rect 22662 21734 22674 21786
rect 22726 21734 22738 21786
rect 22790 21734 22802 21786
rect 22854 21734 22866 21786
rect 22918 21734 27610 21786
rect 27662 21734 27674 21786
rect 27726 21734 27738 21786
rect 27790 21734 27802 21786
rect 27854 21734 27866 21786
rect 27918 21734 32610 21786
rect 32662 21734 32674 21786
rect 32726 21734 32738 21786
rect 32790 21734 32802 21786
rect 32854 21734 32866 21786
rect 32918 21734 37610 21786
rect 37662 21734 37674 21786
rect 37726 21734 37738 21786
rect 37790 21734 37802 21786
rect 37854 21734 37866 21786
rect 37918 21734 42610 21786
rect 42662 21734 42674 21786
rect 42726 21734 42738 21786
rect 42790 21734 42802 21786
rect 42854 21734 42866 21786
rect 42918 21734 47610 21786
rect 47662 21734 47674 21786
rect 47726 21734 47738 21786
rect 47790 21734 47802 21786
rect 47854 21734 47866 21786
rect 47918 21734 52610 21786
rect 52662 21734 52674 21786
rect 52726 21734 52738 21786
rect 52790 21734 52802 21786
rect 52854 21734 52866 21786
rect 52918 21734 57610 21786
rect 57662 21734 57674 21786
rect 57726 21734 57738 21786
rect 57790 21734 57802 21786
rect 57854 21734 57866 21786
rect 57918 21734 58880 21786
rect 1104 21712 58880 21734
rect 58526 21292 58532 21344
rect 58584 21292 58590 21344
rect 1104 21242 58880 21264
rect 1104 21190 1950 21242
rect 2002 21190 2014 21242
rect 2066 21190 2078 21242
rect 2130 21190 2142 21242
rect 2194 21190 2206 21242
rect 2258 21190 6950 21242
rect 7002 21190 7014 21242
rect 7066 21190 7078 21242
rect 7130 21190 7142 21242
rect 7194 21190 7206 21242
rect 7258 21190 11950 21242
rect 12002 21190 12014 21242
rect 12066 21190 12078 21242
rect 12130 21190 12142 21242
rect 12194 21190 12206 21242
rect 12258 21190 16950 21242
rect 17002 21190 17014 21242
rect 17066 21190 17078 21242
rect 17130 21190 17142 21242
rect 17194 21190 17206 21242
rect 17258 21190 21950 21242
rect 22002 21190 22014 21242
rect 22066 21190 22078 21242
rect 22130 21190 22142 21242
rect 22194 21190 22206 21242
rect 22258 21190 26950 21242
rect 27002 21190 27014 21242
rect 27066 21190 27078 21242
rect 27130 21190 27142 21242
rect 27194 21190 27206 21242
rect 27258 21190 31950 21242
rect 32002 21190 32014 21242
rect 32066 21190 32078 21242
rect 32130 21190 32142 21242
rect 32194 21190 32206 21242
rect 32258 21190 36950 21242
rect 37002 21190 37014 21242
rect 37066 21190 37078 21242
rect 37130 21190 37142 21242
rect 37194 21190 37206 21242
rect 37258 21190 41950 21242
rect 42002 21190 42014 21242
rect 42066 21190 42078 21242
rect 42130 21190 42142 21242
rect 42194 21190 42206 21242
rect 42258 21190 46950 21242
rect 47002 21190 47014 21242
rect 47066 21190 47078 21242
rect 47130 21190 47142 21242
rect 47194 21190 47206 21242
rect 47258 21190 51950 21242
rect 52002 21190 52014 21242
rect 52066 21190 52078 21242
rect 52130 21190 52142 21242
rect 52194 21190 52206 21242
rect 52258 21190 56950 21242
rect 57002 21190 57014 21242
rect 57066 21190 57078 21242
rect 57130 21190 57142 21242
rect 57194 21190 57206 21242
rect 57258 21190 58880 21242
rect 1104 21168 58880 21190
rect 58526 20884 58532 20936
rect 58584 20884 58590 20936
rect 1104 20698 58880 20720
rect 1104 20646 2610 20698
rect 2662 20646 2674 20698
rect 2726 20646 2738 20698
rect 2790 20646 2802 20698
rect 2854 20646 2866 20698
rect 2918 20646 7610 20698
rect 7662 20646 7674 20698
rect 7726 20646 7738 20698
rect 7790 20646 7802 20698
rect 7854 20646 7866 20698
rect 7918 20646 12610 20698
rect 12662 20646 12674 20698
rect 12726 20646 12738 20698
rect 12790 20646 12802 20698
rect 12854 20646 12866 20698
rect 12918 20646 17610 20698
rect 17662 20646 17674 20698
rect 17726 20646 17738 20698
rect 17790 20646 17802 20698
rect 17854 20646 17866 20698
rect 17918 20646 22610 20698
rect 22662 20646 22674 20698
rect 22726 20646 22738 20698
rect 22790 20646 22802 20698
rect 22854 20646 22866 20698
rect 22918 20646 27610 20698
rect 27662 20646 27674 20698
rect 27726 20646 27738 20698
rect 27790 20646 27802 20698
rect 27854 20646 27866 20698
rect 27918 20646 32610 20698
rect 32662 20646 32674 20698
rect 32726 20646 32738 20698
rect 32790 20646 32802 20698
rect 32854 20646 32866 20698
rect 32918 20646 37610 20698
rect 37662 20646 37674 20698
rect 37726 20646 37738 20698
rect 37790 20646 37802 20698
rect 37854 20646 37866 20698
rect 37918 20646 42610 20698
rect 42662 20646 42674 20698
rect 42726 20646 42738 20698
rect 42790 20646 42802 20698
rect 42854 20646 42866 20698
rect 42918 20646 47610 20698
rect 47662 20646 47674 20698
rect 47726 20646 47738 20698
rect 47790 20646 47802 20698
rect 47854 20646 47866 20698
rect 47918 20646 52610 20698
rect 52662 20646 52674 20698
rect 52726 20646 52738 20698
rect 52790 20646 52802 20698
rect 52854 20646 52866 20698
rect 52918 20646 57610 20698
rect 57662 20646 57674 20698
rect 57726 20646 57738 20698
rect 57790 20646 57802 20698
rect 57854 20646 57866 20698
rect 57918 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 1950 20154
rect 2002 20102 2014 20154
rect 2066 20102 2078 20154
rect 2130 20102 2142 20154
rect 2194 20102 2206 20154
rect 2258 20102 6950 20154
rect 7002 20102 7014 20154
rect 7066 20102 7078 20154
rect 7130 20102 7142 20154
rect 7194 20102 7206 20154
rect 7258 20102 11950 20154
rect 12002 20102 12014 20154
rect 12066 20102 12078 20154
rect 12130 20102 12142 20154
rect 12194 20102 12206 20154
rect 12258 20102 16950 20154
rect 17002 20102 17014 20154
rect 17066 20102 17078 20154
rect 17130 20102 17142 20154
rect 17194 20102 17206 20154
rect 17258 20102 21950 20154
rect 22002 20102 22014 20154
rect 22066 20102 22078 20154
rect 22130 20102 22142 20154
rect 22194 20102 22206 20154
rect 22258 20102 26950 20154
rect 27002 20102 27014 20154
rect 27066 20102 27078 20154
rect 27130 20102 27142 20154
rect 27194 20102 27206 20154
rect 27258 20102 31950 20154
rect 32002 20102 32014 20154
rect 32066 20102 32078 20154
rect 32130 20102 32142 20154
rect 32194 20102 32206 20154
rect 32258 20102 36950 20154
rect 37002 20102 37014 20154
rect 37066 20102 37078 20154
rect 37130 20102 37142 20154
rect 37194 20102 37206 20154
rect 37258 20102 41950 20154
rect 42002 20102 42014 20154
rect 42066 20102 42078 20154
rect 42130 20102 42142 20154
rect 42194 20102 42206 20154
rect 42258 20102 46950 20154
rect 47002 20102 47014 20154
rect 47066 20102 47078 20154
rect 47130 20102 47142 20154
rect 47194 20102 47206 20154
rect 47258 20102 51950 20154
rect 52002 20102 52014 20154
rect 52066 20102 52078 20154
rect 52130 20102 52142 20154
rect 52194 20102 52206 20154
rect 52258 20102 56950 20154
rect 57002 20102 57014 20154
rect 57066 20102 57078 20154
rect 57130 20102 57142 20154
rect 57194 20102 57206 20154
rect 57258 20102 58880 20154
rect 1104 20080 58880 20102
rect 58526 19796 58532 19848
rect 58584 19796 58590 19848
rect 1104 19610 58880 19632
rect 1104 19558 2610 19610
rect 2662 19558 2674 19610
rect 2726 19558 2738 19610
rect 2790 19558 2802 19610
rect 2854 19558 2866 19610
rect 2918 19558 7610 19610
rect 7662 19558 7674 19610
rect 7726 19558 7738 19610
rect 7790 19558 7802 19610
rect 7854 19558 7866 19610
rect 7918 19558 12610 19610
rect 12662 19558 12674 19610
rect 12726 19558 12738 19610
rect 12790 19558 12802 19610
rect 12854 19558 12866 19610
rect 12918 19558 17610 19610
rect 17662 19558 17674 19610
rect 17726 19558 17738 19610
rect 17790 19558 17802 19610
rect 17854 19558 17866 19610
rect 17918 19558 22610 19610
rect 22662 19558 22674 19610
rect 22726 19558 22738 19610
rect 22790 19558 22802 19610
rect 22854 19558 22866 19610
rect 22918 19558 27610 19610
rect 27662 19558 27674 19610
rect 27726 19558 27738 19610
rect 27790 19558 27802 19610
rect 27854 19558 27866 19610
rect 27918 19558 32610 19610
rect 32662 19558 32674 19610
rect 32726 19558 32738 19610
rect 32790 19558 32802 19610
rect 32854 19558 32866 19610
rect 32918 19558 37610 19610
rect 37662 19558 37674 19610
rect 37726 19558 37738 19610
rect 37790 19558 37802 19610
rect 37854 19558 37866 19610
rect 37918 19558 42610 19610
rect 42662 19558 42674 19610
rect 42726 19558 42738 19610
rect 42790 19558 42802 19610
rect 42854 19558 42866 19610
rect 42918 19558 47610 19610
rect 47662 19558 47674 19610
rect 47726 19558 47738 19610
rect 47790 19558 47802 19610
rect 47854 19558 47866 19610
rect 47918 19558 52610 19610
rect 52662 19558 52674 19610
rect 52726 19558 52738 19610
rect 52790 19558 52802 19610
rect 52854 19558 52866 19610
rect 52918 19558 57610 19610
rect 57662 19558 57674 19610
rect 57726 19558 57738 19610
rect 57790 19558 57802 19610
rect 57854 19558 57866 19610
rect 57918 19558 58880 19610
rect 1104 19536 58880 19558
rect 58526 19116 58532 19168
rect 58584 19116 58590 19168
rect 1104 19066 58880 19088
rect 1104 19014 1950 19066
rect 2002 19014 2014 19066
rect 2066 19014 2078 19066
rect 2130 19014 2142 19066
rect 2194 19014 2206 19066
rect 2258 19014 6950 19066
rect 7002 19014 7014 19066
rect 7066 19014 7078 19066
rect 7130 19014 7142 19066
rect 7194 19014 7206 19066
rect 7258 19014 11950 19066
rect 12002 19014 12014 19066
rect 12066 19014 12078 19066
rect 12130 19014 12142 19066
rect 12194 19014 12206 19066
rect 12258 19014 16950 19066
rect 17002 19014 17014 19066
rect 17066 19014 17078 19066
rect 17130 19014 17142 19066
rect 17194 19014 17206 19066
rect 17258 19014 21950 19066
rect 22002 19014 22014 19066
rect 22066 19014 22078 19066
rect 22130 19014 22142 19066
rect 22194 19014 22206 19066
rect 22258 19014 26950 19066
rect 27002 19014 27014 19066
rect 27066 19014 27078 19066
rect 27130 19014 27142 19066
rect 27194 19014 27206 19066
rect 27258 19014 31950 19066
rect 32002 19014 32014 19066
rect 32066 19014 32078 19066
rect 32130 19014 32142 19066
rect 32194 19014 32206 19066
rect 32258 19014 36950 19066
rect 37002 19014 37014 19066
rect 37066 19014 37078 19066
rect 37130 19014 37142 19066
rect 37194 19014 37206 19066
rect 37258 19014 41950 19066
rect 42002 19014 42014 19066
rect 42066 19014 42078 19066
rect 42130 19014 42142 19066
rect 42194 19014 42206 19066
rect 42258 19014 46950 19066
rect 47002 19014 47014 19066
rect 47066 19014 47078 19066
rect 47130 19014 47142 19066
rect 47194 19014 47206 19066
rect 47258 19014 51950 19066
rect 52002 19014 52014 19066
rect 52066 19014 52078 19066
rect 52130 19014 52142 19066
rect 52194 19014 52206 19066
rect 52258 19014 56950 19066
rect 57002 19014 57014 19066
rect 57066 19014 57078 19066
rect 57130 19014 57142 19066
rect 57194 19014 57206 19066
rect 57258 19014 58880 19066
rect 1104 18992 58880 19014
rect 1104 18522 58880 18544
rect 1104 18470 2610 18522
rect 2662 18470 2674 18522
rect 2726 18470 2738 18522
rect 2790 18470 2802 18522
rect 2854 18470 2866 18522
rect 2918 18470 7610 18522
rect 7662 18470 7674 18522
rect 7726 18470 7738 18522
rect 7790 18470 7802 18522
rect 7854 18470 7866 18522
rect 7918 18470 12610 18522
rect 12662 18470 12674 18522
rect 12726 18470 12738 18522
rect 12790 18470 12802 18522
rect 12854 18470 12866 18522
rect 12918 18470 17610 18522
rect 17662 18470 17674 18522
rect 17726 18470 17738 18522
rect 17790 18470 17802 18522
rect 17854 18470 17866 18522
rect 17918 18470 22610 18522
rect 22662 18470 22674 18522
rect 22726 18470 22738 18522
rect 22790 18470 22802 18522
rect 22854 18470 22866 18522
rect 22918 18470 27610 18522
rect 27662 18470 27674 18522
rect 27726 18470 27738 18522
rect 27790 18470 27802 18522
rect 27854 18470 27866 18522
rect 27918 18470 32610 18522
rect 32662 18470 32674 18522
rect 32726 18470 32738 18522
rect 32790 18470 32802 18522
rect 32854 18470 32866 18522
rect 32918 18470 37610 18522
rect 37662 18470 37674 18522
rect 37726 18470 37738 18522
rect 37790 18470 37802 18522
rect 37854 18470 37866 18522
rect 37918 18470 42610 18522
rect 42662 18470 42674 18522
rect 42726 18470 42738 18522
rect 42790 18470 42802 18522
rect 42854 18470 42866 18522
rect 42918 18470 47610 18522
rect 47662 18470 47674 18522
rect 47726 18470 47738 18522
rect 47790 18470 47802 18522
rect 47854 18470 47866 18522
rect 47918 18470 52610 18522
rect 52662 18470 52674 18522
rect 52726 18470 52738 18522
rect 52790 18470 52802 18522
rect 52854 18470 52866 18522
rect 52918 18470 57610 18522
rect 57662 18470 57674 18522
rect 57726 18470 57738 18522
rect 57790 18470 57802 18522
rect 57854 18470 57866 18522
rect 57918 18470 58880 18522
rect 1104 18448 58880 18470
rect 58526 18028 58532 18080
rect 58584 18028 58590 18080
rect 1104 17978 58880 18000
rect 1104 17926 1950 17978
rect 2002 17926 2014 17978
rect 2066 17926 2078 17978
rect 2130 17926 2142 17978
rect 2194 17926 2206 17978
rect 2258 17926 6950 17978
rect 7002 17926 7014 17978
rect 7066 17926 7078 17978
rect 7130 17926 7142 17978
rect 7194 17926 7206 17978
rect 7258 17926 11950 17978
rect 12002 17926 12014 17978
rect 12066 17926 12078 17978
rect 12130 17926 12142 17978
rect 12194 17926 12206 17978
rect 12258 17926 16950 17978
rect 17002 17926 17014 17978
rect 17066 17926 17078 17978
rect 17130 17926 17142 17978
rect 17194 17926 17206 17978
rect 17258 17926 21950 17978
rect 22002 17926 22014 17978
rect 22066 17926 22078 17978
rect 22130 17926 22142 17978
rect 22194 17926 22206 17978
rect 22258 17926 26950 17978
rect 27002 17926 27014 17978
rect 27066 17926 27078 17978
rect 27130 17926 27142 17978
rect 27194 17926 27206 17978
rect 27258 17926 31950 17978
rect 32002 17926 32014 17978
rect 32066 17926 32078 17978
rect 32130 17926 32142 17978
rect 32194 17926 32206 17978
rect 32258 17926 36950 17978
rect 37002 17926 37014 17978
rect 37066 17926 37078 17978
rect 37130 17926 37142 17978
rect 37194 17926 37206 17978
rect 37258 17926 41950 17978
rect 42002 17926 42014 17978
rect 42066 17926 42078 17978
rect 42130 17926 42142 17978
rect 42194 17926 42206 17978
rect 42258 17926 46950 17978
rect 47002 17926 47014 17978
rect 47066 17926 47078 17978
rect 47130 17926 47142 17978
rect 47194 17926 47206 17978
rect 47258 17926 51950 17978
rect 52002 17926 52014 17978
rect 52066 17926 52078 17978
rect 52130 17926 52142 17978
rect 52194 17926 52206 17978
rect 52258 17926 56950 17978
rect 57002 17926 57014 17978
rect 57066 17926 57078 17978
rect 57130 17926 57142 17978
rect 57194 17926 57206 17978
rect 57258 17926 58880 17978
rect 1104 17904 58880 17926
rect 58526 17620 58532 17672
rect 58584 17620 58590 17672
rect 1104 17434 58880 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 22610 17434
rect 22662 17382 22674 17434
rect 22726 17382 22738 17434
rect 22790 17382 22802 17434
rect 22854 17382 22866 17434
rect 22918 17382 27610 17434
rect 27662 17382 27674 17434
rect 27726 17382 27738 17434
rect 27790 17382 27802 17434
rect 27854 17382 27866 17434
rect 27918 17382 32610 17434
rect 32662 17382 32674 17434
rect 32726 17382 32738 17434
rect 32790 17382 32802 17434
rect 32854 17382 32866 17434
rect 32918 17382 37610 17434
rect 37662 17382 37674 17434
rect 37726 17382 37738 17434
rect 37790 17382 37802 17434
rect 37854 17382 37866 17434
rect 37918 17382 42610 17434
rect 42662 17382 42674 17434
rect 42726 17382 42738 17434
rect 42790 17382 42802 17434
rect 42854 17382 42866 17434
rect 42918 17382 47610 17434
rect 47662 17382 47674 17434
rect 47726 17382 47738 17434
rect 47790 17382 47802 17434
rect 47854 17382 47866 17434
rect 47918 17382 52610 17434
rect 52662 17382 52674 17434
rect 52726 17382 52738 17434
rect 52790 17382 52802 17434
rect 52854 17382 52866 17434
rect 52918 17382 57610 17434
rect 57662 17382 57674 17434
rect 57726 17382 57738 17434
rect 57790 17382 57802 17434
rect 57854 17382 57866 17434
rect 57918 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 21950 16890
rect 22002 16838 22014 16890
rect 22066 16838 22078 16890
rect 22130 16838 22142 16890
rect 22194 16838 22206 16890
rect 22258 16838 26950 16890
rect 27002 16838 27014 16890
rect 27066 16838 27078 16890
rect 27130 16838 27142 16890
rect 27194 16838 27206 16890
rect 27258 16838 31950 16890
rect 32002 16838 32014 16890
rect 32066 16838 32078 16890
rect 32130 16838 32142 16890
rect 32194 16838 32206 16890
rect 32258 16838 36950 16890
rect 37002 16838 37014 16890
rect 37066 16838 37078 16890
rect 37130 16838 37142 16890
rect 37194 16838 37206 16890
rect 37258 16838 41950 16890
rect 42002 16838 42014 16890
rect 42066 16838 42078 16890
rect 42130 16838 42142 16890
rect 42194 16838 42206 16890
rect 42258 16838 46950 16890
rect 47002 16838 47014 16890
rect 47066 16838 47078 16890
rect 47130 16838 47142 16890
rect 47194 16838 47206 16890
rect 47258 16838 51950 16890
rect 52002 16838 52014 16890
rect 52066 16838 52078 16890
rect 52130 16838 52142 16890
rect 52194 16838 52206 16890
rect 52258 16838 56950 16890
rect 57002 16838 57014 16890
rect 57066 16838 57078 16890
rect 57130 16838 57142 16890
rect 57194 16838 57206 16890
rect 57258 16838 58880 16890
rect 1104 16816 58880 16838
rect 57974 16600 57980 16652
rect 58032 16640 58038 16652
rect 58529 16643 58587 16649
rect 58529 16640 58541 16643
rect 58032 16612 58541 16640
rect 58032 16600 58038 16612
rect 58529 16609 58541 16612
rect 58575 16609 58587 16643
rect 58529 16603 58587 16609
rect 1104 16346 58880 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 22610 16346
rect 22662 16294 22674 16346
rect 22726 16294 22738 16346
rect 22790 16294 22802 16346
rect 22854 16294 22866 16346
rect 22918 16294 27610 16346
rect 27662 16294 27674 16346
rect 27726 16294 27738 16346
rect 27790 16294 27802 16346
rect 27854 16294 27866 16346
rect 27918 16294 32610 16346
rect 32662 16294 32674 16346
rect 32726 16294 32738 16346
rect 32790 16294 32802 16346
rect 32854 16294 32866 16346
rect 32918 16294 37610 16346
rect 37662 16294 37674 16346
rect 37726 16294 37738 16346
rect 37790 16294 37802 16346
rect 37854 16294 37866 16346
rect 37918 16294 42610 16346
rect 42662 16294 42674 16346
rect 42726 16294 42738 16346
rect 42790 16294 42802 16346
rect 42854 16294 42866 16346
rect 42918 16294 47610 16346
rect 47662 16294 47674 16346
rect 47726 16294 47738 16346
rect 47790 16294 47802 16346
rect 47854 16294 47866 16346
rect 47918 16294 52610 16346
rect 52662 16294 52674 16346
rect 52726 16294 52738 16346
rect 52790 16294 52802 16346
rect 52854 16294 52866 16346
rect 52918 16294 57610 16346
rect 57662 16294 57674 16346
rect 57726 16294 57738 16346
rect 57790 16294 57802 16346
rect 57854 16294 57866 16346
rect 57918 16294 58880 16346
rect 1104 16272 58880 16294
rect 58526 15852 58532 15904
rect 58584 15852 58590 15904
rect 1104 15802 58880 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 21950 15802
rect 22002 15750 22014 15802
rect 22066 15750 22078 15802
rect 22130 15750 22142 15802
rect 22194 15750 22206 15802
rect 22258 15750 26950 15802
rect 27002 15750 27014 15802
rect 27066 15750 27078 15802
rect 27130 15750 27142 15802
rect 27194 15750 27206 15802
rect 27258 15750 31950 15802
rect 32002 15750 32014 15802
rect 32066 15750 32078 15802
rect 32130 15750 32142 15802
rect 32194 15750 32206 15802
rect 32258 15750 36950 15802
rect 37002 15750 37014 15802
rect 37066 15750 37078 15802
rect 37130 15750 37142 15802
rect 37194 15750 37206 15802
rect 37258 15750 41950 15802
rect 42002 15750 42014 15802
rect 42066 15750 42078 15802
rect 42130 15750 42142 15802
rect 42194 15750 42206 15802
rect 42258 15750 46950 15802
rect 47002 15750 47014 15802
rect 47066 15750 47078 15802
rect 47130 15750 47142 15802
rect 47194 15750 47206 15802
rect 47258 15750 51950 15802
rect 52002 15750 52014 15802
rect 52066 15750 52078 15802
rect 52130 15750 52142 15802
rect 52194 15750 52206 15802
rect 52258 15750 56950 15802
rect 57002 15750 57014 15802
rect 57066 15750 57078 15802
rect 57130 15750 57142 15802
rect 57194 15750 57206 15802
rect 57258 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 22610 15258
rect 22662 15206 22674 15258
rect 22726 15206 22738 15258
rect 22790 15206 22802 15258
rect 22854 15206 22866 15258
rect 22918 15206 27610 15258
rect 27662 15206 27674 15258
rect 27726 15206 27738 15258
rect 27790 15206 27802 15258
rect 27854 15206 27866 15258
rect 27918 15206 32610 15258
rect 32662 15206 32674 15258
rect 32726 15206 32738 15258
rect 32790 15206 32802 15258
rect 32854 15206 32866 15258
rect 32918 15206 37610 15258
rect 37662 15206 37674 15258
rect 37726 15206 37738 15258
rect 37790 15206 37802 15258
rect 37854 15206 37866 15258
rect 37918 15206 42610 15258
rect 42662 15206 42674 15258
rect 42726 15206 42738 15258
rect 42790 15206 42802 15258
rect 42854 15206 42866 15258
rect 42918 15206 47610 15258
rect 47662 15206 47674 15258
rect 47726 15206 47738 15258
rect 47790 15206 47802 15258
rect 47854 15206 47866 15258
rect 47918 15206 52610 15258
rect 52662 15206 52674 15258
rect 52726 15206 52738 15258
rect 52790 15206 52802 15258
rect 52854 15206 52866 15258
rect 52918 15206 57610 15258
rect 57662 15206 57674 15258
rect 57726 15206 57738 15258
rect 57790 15206 57802 15258
rect 57854 15206 57866 15258
rect 57918 15206 58880 15258
rect 1104 15184 58880 15206
rect 58526 14764 58532 14816
rect 58584 14764 58590 14816
rect 1104 14714 58880 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 21950 14714
rect 22002 14662 22014 14714
rect 22066 14662 22078 14714
rect 22130 14662 22142 14714
rect 22194 14662 22206 14714
rect 22258 14662 26950 14714
rect 27002 14662 27014 14714
rect 27066 14662 27078 14714
rect 27130 14662 27142 14714
rect 27194 14662 27206 14714
rect 27258 14662 31950 14714
rect 32002 14662 32014 14714
rect 32066 14662 32078 14714
rect 32130 14662 32142 14714
rect 32194 14662 32206 14714
rect 32258 14662 36950 14714
rect 37002 14662 37014 14714
rect 37066 14662 37078 14714
rect 37130 14662 37142 14714
rect 37194 14662 37206 14714
rect 37258 14662 41950 14714
rect 42002 14662 42014 14714
rect 42066 14662 42078 14714
rect 42130 14662 42142 14714
rect 42194 14662 42206 14714
rect 42258 14662 46950 14714
rect 47002 14662 47014 14714
rect 47066 14662 47078 14714
rect 47130 14662 47142 14714
rect 47194 14662 47206 14714
rect 47258 14662 51950 14714
rect 52002 14662 52014 14714
rect 52066 14662 52078 14714
rect 52130 14662 52142 14714
rect 52194 14662 52206 14714
rect 52258 14662 56950 14714
rect 57002 14662 57014 14714
rect 57066 14662 57078 14714
rect 57130 14662 57142 14714
rect 57194 14662 57206 14714
rect 57258 14662 58880 14714
rect 1104 14640 58880 14662
rect 58526 14356 58532 14408
rect 58584 14356 58590 14408
rect 1104 14170 58880 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 22610 14170
rect 22662 14118 22674 14170
rect 22726 14118 22738 14170
rect 22790 14118 22802 14170
rect 22854 14118 22866 14170
rect 22918 14118 27610 14170
rect 27662 14118 27674 14170
rect 27726 14118 27738 14170
rect 27790 14118 27802 14170
rect 27854 14118 27866 14170
rect 27918 14118 32610 14170
rect 32662 14118 32674 14170
rect 32726 14118 32738 14170
rect 32790 14118 32802 14170
rect 32854 14118 32866 14170
rect 32918 14118 37610 14170
rect 37662 14118 37674 14170
rect 37726 14118 37738 14170
rect 37790 14118 37802 14170
rect 37854 14118 37866 14170
rect 37918 14118 42610 14170
rect 42662 14118 42674 14170
rect 42726 14118 42738 14170
rect 42790 14118 42802 14170
rect 42854 14118 42866 14170
rect 42918 14118 47610 14170
rect 47662 14118 47674 14170
rect 47726 14118 47738 14170
rect 47790 14118 47802 14170
rect 47854 14118 47866 14170
rect 47918 14118 52610 14170
rect 52662 14118 52674 14170
rect 52726 14118 52738 14170
rect 52790 14118 52802 14170
rect 52854 14118 52866 14170
rect 52918 14118 57610 14170
rect 57662 14118 57674 14170
rect 57726 14118 57738 14170
rect 57790 14118 57802 14170
rect 57854 14118 57866 14170
rect 57918 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 21950 13626
rect 22002 13574 22014 13626
rect 22066 13574 22078 13626
rect 22130 13574 22142 13626
rect 22194 13574 22206 13626
rect 22258 13574 26950 13626
rect 27002 13574 27014 13626
rect 27066 13574 27078 13626
rect 27130 13574 27142 13626
rect 27194 13574 27206 13626
rect 27258 13574 31950 13626
rect 32002 13574 32014 13626
rect 32066 13574 32078 13626
rect 32130 13574 32142 13626
rect 32194 13574 32206 13626
rect 32258 13574 36950 13626
rect 37002 13574 37014 13626
rect 37066 13574 37078 13626
rect 37130 13574 37142 13626
rect 37194 13574 37206 13626
rect 37258 13574 41950 13626
rect 42002 13574 42014 13626
rect 42066 13574 42078 13626
rect 42130 13574 42142 13626
rect 42194 13574 42206 13626
rect 42258 13574 46950 13626
rect 47002 13574 47014 13626
rect 47066 13574 47078 13626
rect 47130 13574 47142 13626
rect 47194 13574 47206 13626
rect 47258 13574 51950 13626
rect 52002 13574 52014 13626
rect 52066 13574 52078 13626
rect 52130 13574 52142 13626
rect 52194 13574 52206 13626
rect 52258 13574 56950 13626
rect 57002 13574 57014 13626
rect 57066 13574 57078 13626
rect 57130 13574 57142 13626
rect 57194 13574 57206 13626
rect 57258 13574 58880 13626
rect 1104 13552 58880 13574
rect 58526 13268 58532 13320
rect 58584 13268 58590 13320
rect 1104 13082 58880 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 22610 13082
rect 22662 13030 22674 13082
rect 22726 13030 22738 13082
rect 22790 13030 22802 13082
rect 22854 13030 22866 13082
rect 22918 13030 27610 13082
rect 27662 13030 27674 13082
rect 27726 13030 27738 13082
rect 27790 13030 27802 13082
rect 27854 13030 27866 13082
rect 27918 13030 32610 13082
rect 32662 13030 32674 13082
rect 32726 13030 32738 13082
rect 32790 13030 32802 13082
rect 32854 13030 32866 13082
rect 32918 13030 37610 13082
rect 37662 13030 37674 13082
rect 37726 13030 37738 13082
rect 37790 13030 37802 13082
rect 37854 13030 37866 13082
rect 37918 13030 42610 13082
rect 42662 13030 42674 13082
rect 42726 13030 42738 13082
rect 42790 13030 42802 13082
rect 42854 13030 42866 13082
rect 42918 13030 47610 13082
rect 47662 13030 47674 13082
rect 47726 13030 47738 13082
rect 47790 13030 47802 13082
rect 47854 13030 47866 13082
rect 47918 13030 52610 13082
rect 52662 13030 52674 13082
rect 52726 13030 52738 13082
rect 52790 13030 52802 13082
rect 52854 13030 52866 13082
rect 52918 13030 57610 13082
rect 57662 13030 57674 13082
rect 57726 13030 57738 13082
rect 57790 13030 57802 13082
rect 57854 13030 57866 13082
rect 57918 13030 58880 13082
rect 1104 13008 58880 13030
rect 58526 12588 58532 12640
rect 58584 12588 58590 12640
rect 1104 12538 58880 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 21950 12538
rect 22002 12486 22014 12538
rect 22066 12486 22078 12538
rect 22130 12486 22142 12538
rect 22194 12486 22206 12538
rect 22258 12486 26950 12538
rect 27002 12486 27014 12538
rect 27066 12486 27078 12538
rect 27130 12486 27142 12538
rect 27194 12486 27206 12538
rect 27258 12486 31950 12538
rect 32002 12486 32014 12538
rect 32066 12486 32078 12538
rect 32130 12486 32142 12538
rect 32194 12486 32206 12538
rect 32258 12486 36950 12538
rect 37002 12486 37014 12538
rect 37066 12486 37078 12538
rect 37130 12486 37142 12538
rect 37194 12486 37206 12538
rect 37258 12486 41950 12538
rect 42002 12486 42014 12538
rect 42066 12486 42078 12538
rect 42130 12486 42142 12538
rect 42194 12486 42206 12538
rect 42258 12486 46950 12538
rect 47002 12486 47014 12538
rect 47066 12486 47078 12538
rect 47130 12486 47142 12538
rect 47194 12486 47206 12538
rect 47258 12486 51950 12538
rect 52002 12486 52014 12538
rect 52066 12486 52078 12538
rect 52130 12486 52142 12538
rect 52194 12486 52206 12538
rect 52258 12486 56950 12538
rect 57002 12486 57014 12538
rect 57066 12486 57078 12538
rect 57130 12486 57142 12538
rect 57194 12486 57206 12538
rect 57258 12486 58880 12538
rect 1104 12464 58880 12486
rect 1104 11994 58880 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 22610 11994
rect 22662 11942 22674 11994
rect 22726 11942 22738 11994
rect 22790 11942 22802 11994
rect 22854 11942 22866 11994
rect 22918 11942 27610 11994
rect 27662 11942 27674 11994
rect 27726 11942 27738 11994
rect 27790 11942 27802 11994
rect 27854 11942 27866 11994
rect 27918 11942 32610 11994
rect 32662 11942 32674 11994
rect 32726 11942 32738 11994
rect 32790 11942 32802 11994
rect 32854 11942 32866 11994
rect 32918 11942 37610 11994
rect 37662 11942 37674 11994
rect 37726 11942 37738 11994
rect 37790 11942 37802 11994
rect 37854 11942 37866 11994
rect 37918 11942 42610 11994
rect 42662 11942 42674 11994
rect 42726 11942 42738 11994
rect 42790 11942 42802 11994
rect 42854 11942 42866 11994
rect 42918 11942 47610 11994
rect 47662 11942 47674 11994
rect 47726 11942 47738 11994
rect 47790 11942 47802 11994
rect 47854 11942 47866 11994
rect 47918 11942 52610 11994
rect 52662 11942 52674 11994
rect 52726 11942 52738 11994
rect 52790 11942 52802 11994
rect 52854 11942 52866 11994
rect 52918 11942 57610 11994
rect 57662 11942 57674 11994
rect 57726 11942 57738 11994
rect 57790 11942 57802 11994
rect 57854 11942 57866 11994
rect 57918 11942 58880 11994
rect 1104 11920 58880 11942
rect 58526 11500 58532 11552
rect 58584 11500 58590 11552
rect 1104 11450 58880 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 21950 11450
rect 22002 11398 22014 11450
rect 22066 11398 22078 11450
rect 22130 11398 22142 11450
rect 22194 11398 22206 11450
rect 22258 11398 26950 11450
rect 27002 11398 27014 11450
rect 27066 11398 27078 11450
rect 27130 11398 27142 11450
rect 27194 11398 27206 11450
rect 27258 11398 31950 11450
rect 32002 11398 32014 11450
rect 32066 11398 32078 11450
rect 32130 11398 32142 11450
rect 32194 11398 32206 11450
rect 32258 11398 36950 11450
rect 37002 11398 37014 11450
rect 37066 11398 37078 11450
rect 37130 11398 37142 11450
rect 37194 11398 37206 11450
rect 37258 11398 41950 11450
rect 42002 11398 42014 11450
rect 42066 11398 42078 11450
rect 42130 11398 42142 11450
rect 42194 11398 42206 11450
rect 42258 11398 46950 11450
rect 47002 11398 47014 11450
rect 47066 11398 47078 11450
rect 47130 11398 47142 11450
rect 47194 11398 47206 11450
rect 47258 11398 51950 11450
rect 52002 11398 52014 11450
rect 52066 11398 52078 11450
rect 52130 11398 52142 11450
rect 52194 11398 52206 11450
rect 52258 11398 56950 11450
rect 57002 11398 57014 11450
rect 57066 11398 57078 11450
rect 57130 11398 57142 11450
rect 57194 11398 57206 11450
rect 57258 11398 58880 11450
rect 1104 11376 58880 11398
rect 58526 11092 58532 11144
rect 58584 11092 58590 11144
rect 1104 10906 58880 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 22610 10906
rect 22662 10854 22674 10906
rect 22726 10854 22738 10906
rect 22790 10854 22802 10906
rect 22854 10854 22866 10906
rect 22918 10854 27610 10906
rect 27662 10854 27674 10906
rect 27726 10854 27738 10906
rect 27790 10854 27802 10906
rect 27854 10854 27866 10906
rect 27918 10854 32610 10906
rect 32662 10854 32674 10906
rect 32726 10854 32738 10906
rect 32790 10854 32802 10906
rect 32854 10854 32866 10906
rect 32918 10854 37610 10906
rect 37662 10854 37674 10906
rect 37726 10854 37738 10906
rect 37790 10854 37802 10906
rect 37854 10854 37866 10906
rect 37918 10854 42610 10906
rect 42662 10854 42674 10906
rect 42726 10854 42738 10906
rect 42790 10854 42802 10906
rect 42854 10854 42866 10906
rect 42918 10854 47610 10906
rect 47662 10854 47674 10906
rect 47726 10854 47738 10906
rect 47790 10854 47802 10906
rect 47854 10854 47866 10906
rect 47918 10854 52610 10906
rect 52662 10854 52674 10906
rect 52726 10854 52738 10906
rect 52790 10854 52802 10906
rect 52854 10854 52866 10906
rect 52918 10854 57610 10906
rect 57662 10854 57674 10906
rect 57726 10854 57738 10906
rect 57790 10854 57802 10906
rect 57854 10854 57866 10906
rect 57918 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 21950 10362
rect 22002 10310 22014 10362
rect 22066 10310 22078 10362
rect 22130 10310 22142 10362
rect 22194 10310 22206 10362
rect 22258 10310 26950 10362
rect 27002 10310 27014 10362
rect 27066 10310 27078 10362
rect 27130 10310 27142 10362
rect 27194 10310 27206 10362
rect 27258 10310 31950 10362
rect 32002 10310 32014 10362
rect 32066 10310 32078 10362
rect 32130 10310 32142 10362
rect 32194 10310 32206 10362
rect 32258 10310 36950 10362
rect 37002 10310 37014 10362
rect 37066 10310 37078 10362
rect 37130 10310 37142 10362
rect 37194 10310 37206 10362
rect 37258 10310 41950 10362
rect 42002 10310 42014 10362
rect 42066 10310 42078 10362
rect 42130 10310 42142 10362
rect 42194 10310 42206 10362
rect 42258 10310 46950 10362
rect 47002 10310 47014 10362
rect 47066 10310 47078 10362
rect 47130 10310 47142 10362
rect 47194 10310 47206 10362
rect 47258 10310 51950 10362
rect 52002 10310 52014 10362
rect 52066 10310 52078 10362
rect 52130 10310 52142 10362
rect 52194 10310 52206 10362
rect 52258 10310 56950 10362
rect 57002 10310 57014 10362
rect 57066 10310 57078 10362
rect 57130 10310 57142 10362
rect 57194 10310 57206 10362
rect 57258 10310 58880 10362
rect 1104 10288 58880 10310
rect 58526 10004 58532 10056
rect 58584 10004 58590 10056
rect 1104 9818 58880 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 22610 9818
rect 22662 9766 22674 9818
rect 22726 9766 22738 9818
rect 22790 9766 22802 9818
rect 22854 9766 22866 9818
rect 22918 9766 27610 9818
rect 27662 9766 27674 9818
rect 27726 9766 27738 9818
rect 27790 9766 27802 9818
rect 27854 9766 27866 9818
rect 27918 9766 32610 9818
rect 32662 9766 32674 9818
rect 32726 9766 32738 9818
rect 32790 9766 32802 9818
rect 32854 9766 32866 9818
rect 32918 9766 37610 9818
rect 37662 9766 37674 9818
rect 37726 9766 37738 9818
rect 37790 9766 37802 9818
rect 37854 9766 37866 9818
rect 37918 9766 42610 9818
rect 42662 9766 42674 9818
rect 42726 9766 42738 9818
rect 42790 9766 42802 9818
rect 42854 9766 42866 9818
rect 42918 9766 47610 9818
rect 47662 9766 47674 9818
rect 47726 9766 47738 9818
rect 47790 9766 47802 9818
rect 47854 9766 47866 9818
rect 47918 9766 52610 9818
rect 52662 9766 52674 9818
rect 52726 9766 52738 9818
rect 52790 9766 52802 9818
rect 52854 9766 52866 9818
rect 52918 9766 57610 9818
rect 57662 9766 57674 9818
rect 57726 9766 57738 9818
rect 57790 9766 57802 9818
rect 57854 9766 57866 9818
rect 57918 9766 58880 9818
rect 1104 9744 58880 9766
rect 58526 9324 58532 9376
rect 58584 9324 58590 9376
rect 1104 9274 58880 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 21950 9274
rect 22002 9222 22014 9274
rect 22066 9222 22078 9274
rect 22130 9222 22142 9274
rect 22194 9222 22206 9274
rect 22258 9222 26950 9274
rect 27002 9222 27014 9274
rect 27066 9222 27078 9274
rect 27130 9222 27142 9274
rect 27194 9222 27206 9274
rect 27258 9222 31950 9274
rect 32002 9222 32014 9274
rect 32066 9222 32078 9274
rect 32130 9222 32142 9274
rect 32194 9222 32206 9274
rect 32258 9222 36950 9274
rect 37002 9222 37014 9274
rect 37066 9222 37078 9274
rect 37130 9222 37142 9274
rect 37194 9222 37206 9274
rect 37258 9222 41950 9274
rect 42002 9222 42014 9274
rect 42066 9222 42078 9274
rect 42130 9222 42142 9274
rect 42194 9222 42206 9274
rect 42258 9222 46950 9274
rect 47002 9222 47014 9274
rect 47066 9222 47078 9274
rect 47130 9222 47142 9274
rect 47194 9222 47206 9274
rect 47258 9222 51950 9274
rect 52002 9222 52014 9274
rect 52066 9222 52078 9274
rect 52130 9222 52142 9274
rect 52194 9222 52206 9274
rect 52258 9222 56950 9274
rect 57002 9222 57014 9274
rect 57066 9222 57078 9274
rect 57130 9222 57142 9274
rect 57194 9222 57206 9274
rect 57258 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 22610 8730
rect 22662 8678 22674 8730
rect 22726 8678 22738 8730
rect 22790 8678 22802 8730
rect 22854 8678 22866 8730
rect 22918 8678 27610 8730
rect 27662 8678 27674 8730
rect 27726 8678 27738 8730
rect 27790 8678 27802 8730
rect 27854 8678 27866 8730
rect 27918 8678 32610 8730
rect 32662 8678 32674 8730
rect 32726 8678 32738 8730
rect 32790 8678 32802 8730
rect 32854 8678 32866 8730
rect 32918 8678 37610 8730
rect 37662 8678 37674 8730
rect 37726 8678 37738 8730
rect 37790 8678 37802 8730
rect 37854 8678 37866 8730
rect 37918 8678 42610 8730
rect 42662 8678 42674 8730
rect 42726 8678 42738 8730
rect 42790 8678 42802 8730
rect 42854 8678 42866 8730
rect 42918 8678 47610 8730
rect 47662 8678 47674 8730
rect 47726 8678 47738 8730
rect 47790 8678 47802 8730
rect 47854 8678 47866 8730
rect 47918 8678 52610 8730
rect 52662 8678 52674 8730
rect 52726 8678 52738 8730
rect 52790 8678 52802 8730
rect 52854 8678 52866 8730
rect 52918 8678 57610 8730
rect 57662 8678 57674 8730
rect 57726 8678 57738 8730
rect 57790 8678 57802 8730
rect 57854 8678 57866 8730
rect 57918 8678 58880 8730
rect 1104 8656 58880 8678
rect 58526 8304 58532 8356
rect 58584 8304 58590 8356
rect 1104 8186 58880 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 21950 8186
rect 22002 8134 22014 8186
rect 22066 8134 22078 8186
rect 22130 8134 22142 8186
rect 22194 8134 22206 8186
rect 22258 8134 26950 8186
rect 27002 8134 27014 8186
rect 27066 8134 27078 8186
rect 27130 8134 27142 8186
rect 27194 8134 27206 8186
rect 27258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 36950 8186
rect 37002 8134 37014 8186
rect 37066 8134 37078 8186
rect 37130 8134 37142 8186
rect 37194 8134 37206 8186
rect 37258 8134 41950 8186
rect 42002 8134 42014 8186
rect 42066 8134 42078 8186
rect 42130 8134 42142 8186
rect 42194 8134 42206 8186
rect 42258 8134 46950 8186
rect 47002 8134 47014 8186
rect 47066 8134 47078 8186
rect 47130 8134 47142 8186
rect 47194 8134 47206 8186
rect 47258 8134 51950 8186
rect 52002 8134 52014 8186
rect 52066 8134 52078 8186
rect 52130 8134 52142 8186
rect 52194 8134 52206 8186
rect 52258 8134 56950 8186
rect 57002 8134 57014 8186
rect 57066 8134 57078 8186
rect 57130 8134 57142 8186
rect 57194 8134 57206 8186
rect 57258 8134 58880 8186
rect 1104 8112 58880 8134
rect 58526 7828 58532 7880
rect 58584 7828 58590 7880
rect 1104 7642 58880 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 22610 7642
rect 22662 7590 22674 7642
rect 22726 7590 22738 7642
rect 22790 7590 22802 7642
rect 22854 7590 22866 7642
rect 22918 7590 27610 7642
rect 27662 7590 27674 7642
rect 27726 7590 27738 7642
rect 27790 7590 27802 7642
rect 27854 7590 27866 7642
rect 27918 7590 32610 7642
rect 32662 7590 32674 7642
rect 32726 7590 32738 7642
rect 32790 7590 32802 7642
rect 32854 7590 32866 7642
rect 32918 7590 37610 7642
rect 37662 7590 37674 7642
rect 37726 7590 37738 7642
rect 37790 7590 37802 7642
rect 37854 7590 37866 7642
rect 37918 7590 42610 7642
rect 42662 7590 42674 7642
rect 42726 7590 42738 7642
rect 42790 7590 42802 7642
rect 42854 7590 42866 7642
rect 42918 7590 47610 7642
rect 47662 7590 47674 7642
rect 47726 7590 47738 7642
rect 47790 7590 47802 7642
rect 47854 7590 47866 7642
rect 47918 7590 52610 7642
rect 52662 7590 52674 7642
rect 52726 7590 52738 7642
rect 52790 7590 52802 7642
rect 52854 7590 52866 7642
rect 52918 7590 57610 7642
rect 57662 7590 57674 7642
rect 57726 7590 57738 7642
rect 57790 7590 57802 7642
rect 57854 7590 57866 7642
rect 57918 7590 58880 7642
rect 1104 7568 58880 7590
rect 1104 7098 58880 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 21950 7098
rect 22002 7046 22014 7098
rect 22066 7046 22078 7098
rect 22130 7046 22142 7098
rect 22194 7046 22206 7098
rect 22258 7046 26950 7098
rect 27002 7046 27014 7098
rect 27066 7046 27078 7098
rect 27130 7046 27142 7098
rect 27194 7046 27206 7098
rect 27258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 36950 7098
rect 37002 7046 37014 7098
rect 37066 7046 37078 7098
rect 37130 7046 37142 7098
rect 37194 7046 37206 7098
rect 37258 7046 41950 7098
rect 42002 7046 42014 7098
rect 42066 7046 42078 7098
rect 42130 7046 42142 7098
rect 42194 7046 42206 7098
rect 42258 7046 46950 7098
rect 47002 7046 47014 7098
rect 47066 7046 47078 7098
rect 47130 7046 47142 7098
rect 47194 7046 47206 7098
rect 47258 7046 51950 7098
rect 52002 7046 52014 7098
rect 52066 7046 52078 7098
rect 52130 7046 52142 7098
rect 52194 7046 52206 7098
rect 52258 7046 56950 7098
rect 57002 7046 57014 7098
rect 57066 7046 57078 7098
rect 57130 7046 57142 7098
rect 57194 7046 57206 7098
rect 57258 7046 58880 7098
rect 1104 7024 58880 7046
rect 58526 6740 58532 6792
rect 58584 6740 58590 6792
rect 1104 6554 58880 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 22610 6554
rect 22662 6502 22674 6554
rect 22726 6502 22738 6554
rect 22790 6502 22802 6554
rect 22854 6502 22866 6554
rect 22918 6502 27610 6554
rect 27662 6502 27674 6554
rect 27726 6502 27738 6554
rect 27790 6502 27802 6554
rect 27854 6502 27866 6554
rect 27918 6502 32610 6554
rect 32662 6502 32674 6554
rect 32726 6502 32738 6554
rect 32790 6502 32802 6554
rect 32854 6502 32866 6554
rect 32918 6502 37610 6554
rect 37662 6502 37674 6554
rect 37726 6502 37738 6554
rect 37790 6502 37802 6554
rect 37854 6502 37866 6554
rect 37918 6502 42610 6554
rect 42662 6502 42674 6554
rect 42726 6502 42738 6554
rect 42790 6502 42802 6554
rect 42854 6502 42866 6554
rect 42918 6502 47610 6554
rect 47662 6502 47674 6554
rect 47726 6502 47738 6554
rect 47790 6502 47802 6554
rect 47854 6502 47866 6554
rect 47918 6502 52610 6554
rect 52662 6502 52674 6554
rect 52726 6502 52738 6554
rect 52790 6502 52802 6554
rect 52854 6502 52866 6554
rect 52918 6502 57610 6554
rect 57662 6502 57674 6554
rect 57726 6502 57738 6554
rect 57790 6502 57802 6554
rect 57854 6502 57866 6554
rect 57918 6502 58880 6554
rect 1104 6480 58880 6502
rect 58526 6060 58532 6112
rect 58584 6060 58590 6112
rect 1104 6010 58880 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 21950 6010
rect 22002 5958 22014 6010
rect 22066 5958 22078 6010
rect 22130 5958 22142 6010
rect 22194 5958 22206 6010
rect 22258 5958 26950 6010
rect 27002 5958 27014 6010
rect 27066 5958 27078 6010
rect 27130 5958 27142 6010
rect 27194 5958 27206 6010
rect 27258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 36950 6010
rect 37002 5958 37014 6010
rect 37066 5958 37078 6010
rect 37130 5958 37142 6010
rect 37194 5958 37206 6010
rect 37258 5958 41950 6010
rect 42002 5958 42014 6010
rect 42066 5958 42078 6010
rect 42130 5958 42142 6010
rect 42194 5958 42206 6010
rect 42258 5958 46950 6010
rect 47002 5958 47014 6010
rect 47066 5958 47078 6010
rect 47130 5958 47142 6010
rect 47194 5958 47206 6010
rect 47258 5958 51950 6010
rect 52002 5958 52014 6010
rect 52066 5958 52078 6010
rect 52130 5958 52142 6010
rect 52194 5958 52206 6010
rect 52258 5958 56950 6010
rect 57002 5958 57014 6010
rect 57066 5958 57078 6010
rect 57130 5958 57142 6010
rect 57194 5958 57206 6010
rect 57258 5958 58880 6010
rect 1104 5936 58880 5958
rect 1104 5466 58880 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 22610 5466
rect 22662 5414 22674 5466
rect 22726 5414 22738 5466
rect 22790 5414 22802 5466
rect 22854 5414 22866 5466
rect 22918 5414 27610 5466
rect 27662 5414 27674 5466
rect 27726 5414 27738 5466
rect 27790 5414 27802 5466
rect 27854 5414 27866 5466
rect 27918 5414 32610 5466
rect 32662 5414 32674 5466
rect 32726 5414 32738 5466
rect 32790 5414 32802 5466
rect 32854 5414 32866 5466
rect 32918 5414 37610 5466
rect 37662 5414 37674 5466
rect 37726 5414 37738 5466
rect 37790 5414 37802 5466
rect 37854 5414 37866 5466
rect 37918 5414 42610 5466
rect 42662 5414 42674 5466
rect 42726 5414 42738 5466
rect 42790 5414 42802 5466
rect 42854 5414 42866 5466
rect 42918 5414 47610 5466
rect 47662 5414 47674 5466
rect 47726 5414 47738 5466
rect 47790 5414 47802 5466
rect 47854 5414 47866 5466
rect 47918 5414 52610 5466
rect 52662 5414 52674 5466
rect 52726 5414 52738 5466
rect 52790 5414 52802 5466
rect 52854 5414 52866 5466
rect 52918 5414 57610 5466
rect 57662 5414 57674 5466
rect 57726 5414 57738 5466
rect 57790 5414 57802 5466
rect 57854 5414 57866 5466
rect 57918 5414 58880 5466
rect 1104 5392 58880 5414
rect 58526 4972 58532 5024
rect 58584 4972 58590 5024
rect 1104 4922 58880 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 21950 4922
rect 22002 4870 22014 4922
rect 22066 4870 22078 4922
rect 22130 4870 22142 4922
rect 22194 4870 22206 4922
rect 22258 4870 26950 4922
rect 27002 4870 27014 4922
rect 27066 4870 27078 4922
rect 27130 4870 27142 4922
rect 27194 4870 27206 4922
rect 27258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 36950 4922
rect 37002 4870 37014 4922
rect 37066 4870 37078 4922
rect 37130 4870 37142 4922
rect 37194 4870 37206 4922
rect 37258 4870 41950 4922
rect 42002 4870 42014 4922
rect 42066 4870 42078 4922
rect 42130 4870 42142 4922
rect 42194 4870 42206 4922
rect 42258 4870 46950 4922
rect 47002 4870 47014 4922
rect 47066 4870 47078 4922
rect 47130 4870 47142 4922
rect 47194 4870 47206 4922
rect 47258 4870 51950 4922
rect 52002 4870 52014 4922
rect 52066 4870 52078 4922
rect 52130 4870 52142 4922
rect 52194 4870 52206 4922
rect 52258 4870 56950 4922
rect 57002 4870 57014 4922
rect 57066 4870 57078 4922
rect 57130 4870 57142 4922
rect 57194 4870 57206 4922
rect 57258 4870 58880 4922
rect 1104 4848 58880 4870
rect 58526 4564 58532 4616
rect 58584 4564 58590 4616
rect 1104 4378 58880 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 22610 4378
rect 22662 4326 22674 4378
rect 22726 4326 22738 4378
rect 22790 4326 22802 4378
rect 22854 4326 22866 4378
rect 22918 4326 27610 4378
rect 27662 4326 27674 4378
rect 27726 4326 27738 4378
rect 27790 4326 27802 4378
rect 27854 4326 27866 4378
rect 27918 4326 32610 4378
rect 32662 4326 32674 4378
rect 32726 4326 32738 4378
rect 32790 4326 32802 4378
rect 32854 4326 32866 4378
rect 32918 4326 37610 4378
rect 37662 4326 37674 4378
rect 37726 4326 37738 4378
rect 37790 4326 37802 4378
rect 37854 4326 37866 4378
rect 37918 4326 42610 4378
rect 42662 4326 42674 4378
rect 42726 4326 42738 4378
rect 42790 4326 42802 4378
rect 42854 4326 42866 4378
rect 42918 4326 47610 4378
rect 47662 4326 47674 4378
rect 47726 4326 47738 4378
rect 47790 4326 47802 4378
rect 47854 4326 47866 4378
rect 47918 4326 52610 4378
rect 52662 4326 52674 4378
rect 52726 4326 52738 4378
rect 52790 4326 52802 4378
rect 52854 4326 52866 4378
rect 52918 4326 57610 4378
rect 57662 4326 57674 4378
rect 57726 4326 57738 4378
rect 57790 4326 57802 4378
rect 57854 4326 57866 4378
rect 57918 4326 58880 4378
rect 1104 4304 58880 4326
rect 1104 3834 58880 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 21950 3834
rect 22002 3782 22014 3834
rect 22066 3782 22078 3834
rect 22130 3782 22142 3834
rect 22194 3782 22206 3834
rect 22258 3782 26950 3834
rect 27002 3782 27014 3834
rect 27066 3782 27078 3834
rect 27130 3782 27142 3834
rect 27194 3782 27206 3834
rect 27258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 36950 3834
rect 37002 3782 37014 3834
rect 37066 3782 37078 3834
rect 37130 3782 37142 3834
rect 37194 3782 37206 3834
rect 37258 3782 41950 3834
rect 42002 3782 42014 3834
rect 42066 3782 42078 3834
rect 42130 3782 42142 3834
rect 42194 3782 42206 3834
rect 42258 3782 46950 3834
rect 47002 3782 47014 3834
rect 47066 3782 47078 3834
rect 47130 3782 47142 3834
rect 47194 3782 47206 3834
rect 47258 3782 51950 3834
rect 52002 3782 52014 3834
rect 52066 3782 52078 3834
rect 52130 3782 52142 3834
rect 52194 3782 52206 3834
rect 52258 3782 56950 3834
rect 57002 3782 57014 3834
rect 57066 3782 57078 3834
rect 57130 3782 57142 3834
rect 57194 3782 57206 3834
rect 57258 3782 58880 3834
rect 1104 3760 58880 3782
rect 1104 3290 58880 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 22610 3290
rect 22662 3238 22674 3290
rect 22726 3238 22738 3290
rect 22790 3238 22802 3290
rect 22854 3238 22866 3290
rect 22918 3238 27610 3290
rect 27662 3238 27674 3290
rect 27726 3238 27738 3290
rect 27790 3238 27802 3290
rect 27854 3238 27866 3290
rect 27918 3238 32610 3290
rect 32662 3238 32674 3290
rect 32726 3238 32738 3290
rect 32790 3238 32802 3290
rect 32854 3238 32866 3290
rect 32918 3238 37610 3290
rect 37662 3238 37674 3290
rect 37726 3238 37738 3290
rect 37790 3238 37802 3290
rect 37854 3238 37866 3290
rect 37918 3238 42610 3290
rect 42662 3238 42674 3290
rect 42726 3238 42738 3290
rect 42790 3238 42802 3290
rect 42854 3238 42866 3290
rect 42918 3238 47610 3290
rect 47662 3238 47674 3290
rect 47726 3238 47738 3290
rect 47790 3238 47802 3290
rect 47854 3238 47866 3290
rect 47918 3238 52610 3290
rect 52662 3238 52674 3290
rect 52726 3238 52738 3290
rect 52790 3238 52802 3290
rect 52854 3238 52866 3290
rect 52918 3238 57610 3290
rect 57662 3238 57674 3290
rect 57726 3238 57738 3290
rect 57790 3238 57802 3290
rect 57854 3238 57866 3290
rect 57918 3238 58880 3290
rect 1104 3216 58880 3238
rect 1104 2746 58880 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 21950 2746
rect 22002 2694 22014 2746
rect 22066 2694 22078 2746
rect 22130 2694 22142 2746
rect 22194 2694 22206 2746
rect 22258 2694 26950 2746
rect 27002 2694 27014 2746
rect 27066 2694 27078 2746
rect 27130 2694 27142 2746
rect 27194 2694 27206 2746
rect 27258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 36950 2746
rect 37002 2694 37014 2746
rect 37066 2694 37078 2746
rect 37130 2694 37142 2746
rect 37194 2694 37206 2746
rect 37258 2694 41950 2746
rect 42002 2694 42014 2746
rect 42066 2694 42078 2746
rect 42130 2694 42142 2746
rect 42194 2694 42206 2746
rect 42258 2694 46950 2746
rect 47002 2694 47014 2746
rect 47066 2694 47078 2746
rect 47130 2694 47142 2746
rect 47194 2694 47206 2746
rect 47258 2694 51950 2746
rect 52002 2694 52014 2746
rect 52066 2694 52078 2746
rect 52130 2694 52142 2746
rect 52194 2694 52206 2746
rect 52258 2694 56950 2746
rect 57002 2694 57014 2746
rect 57066 2694 57078 2746
rect 57130 2694 57142 2746
rect 57194 2694 57206 2746
rect 57258 2694 58880 2746
rect 1104 2672 58880 2694
rect 1104 2202 58880 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 22610 2202
rect 22662 2150 22674 2202
rect 22726 2150 22738 2202
rect 22790 2150 22802 2202
rect 22854 2150 22866 2202
rect 22918 2150 27610 2202
rect 27662 2150 27674 2202
rect 27726 2150 27738 2202
rect 27790 2150 27802 2202
rect 27854 2150 27866 2202
rect 27918 2150 32610 2202
rect 32662 2150 32674 2202
rect 32726 2150 32738 2202
rect 32790 2150 32802 2202
rect 32854 2150 32866 2202
rect 32918 2150 37610 2202
rect 37662 2150 37674 2202
rect 37726 2150 37738 2202
rect 37790 2150 37802 2202
rect 37854 2150 37866 2202
rect 37918 2150 42610 2202
rect 42662 2150 42674 2202
rect 42726 2150 42738 2202
rect 42790 2150 42802 2202
rect 42854 2150 42866 2202
rect 42918 2150 47610 2202
rect 47662 2150 47674 2202
rect 47726 2150 47738 2202
rect 47790 2150 47802 2202
rect 47854 2150 47866 2202
rect 47918 2150 52610 2202
rect 52662 2150 52674 2202
rect 52726 2150 52738 2202
rect 52790 2150 52802 2202
rect 52854 2150 52866 2202
rect 52918 2150 57610 2202
rect 57662 2150 57674 2202
rect 57726 2150 57738 2202
rect 57790 2150 57802 2202
rect 57854 2150 57866 2202
rect 57918 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 2610 57638 2662 57690
rect 2674 57638 2726 57690
rect 2738 57638 2790 57690
rect 2802 57638 2854 57690
rect 2866 57638 2918 57690
rect 7610 57638 7662 57690
rect 7674 57638 7726 57690
rect 7738 57638 7790 57690
rect 7802 57638 7854 57690
rect 7866 57638 7918 57690
rect 12610 57638 12662 57690
rect 12674 57638 12726 57690
rect 12738 57638 12790 57690
rect 12802 57638 12854 57690
rect 12866 57638 12918 57690
rect 17610 57638 17662 57690
rect 17674 57638 17726 57690
rect 17738 57638 17790 57690
rect 17802 57638 17854 57690
rect 17866 57638 17918 57690
rect 22610 57638 22662 57690
rect 22674 57638 22726 57690
rect 22738 57638 22790 57690
rect 22802 57638 22854 57690
rect 22866 57638 22918 57690
rect 27610 57638 27662 57690
rect 27674 57638 27726 57690
rect 27738 57638 27790 57690
rect 27802 57638 27854 57690
rect 27866 57638 27918 57690
rect 32610 57638 32662 57690
rect 32674 57638 32726 57690
rect 32738 57638 32790 57690
rect 32802 57638 32854 57690
rect 32866 57638 32918 57690
rect 37610 57638 37662 57690
rect 37674 57638 37726 57690
rect 37738 57638 37790 57690
rect 37802 57638 37854 57690
rect 37866 57638 37918 57690
rect 42610 57638 42662 57690
rect 42674 57638 42726 57690
rect 42738 57638 42790 57690
rect 42802 57638 42854 57690
rect 42866 57638 42918 57690
rect 47610 57638 47662 57690
rect 47674 57638 47726 57690
rect 47738 57638 47790 57690
rect 47802 57638 47854 57690
rect 47866 57638 47918 57690
rect 52610 57638 52662 57690
rect 52674 57638 52726 57690
rect 52738 57638 52790 57690
rect 52802 57638 52854 57690
rect 52866 57638 52918 57690
rect 57610 57638 57662 57690
rect 57674 57638 57726 57690
rect 57738 57638 57790 57690
rect 57802 57638 57854 57690
rect 57866 57638 57918 57690
rect 1950 57094 2002 57146
rect 2014 57094 2066 57146
rect 2078 57094 2130 57146
rect 2142 57094 2194 57146
rect 2206 57094 2258 57146
rect 6950 57094 7002 57146
rect 7014 57094 7066 57146
rect 7078 57094 7130 57146
rect 7142 57094 7194 57146
rect 7206 57094 7258 57146
rect 11950 57094 12002 57146
rect 12014 57094 12066 57146
rect 12078 57094 12130 57146
rect 12142 57094 12194 57146
rect 12206 57094 12258 57146
rect 16950 57094 17002 57146
rect 17014 57094 17066 57146
rect 17078 57094 17130 57146
rect 17142 57094 17194 57146
rect 17206 57094 17258 57146
rect 21950 57094 22002 57146
rect 22014 57094 22066 57146
rect 22078 57094 22130 57146
rect 22142 57094 22194 57146
rect 22206 57094 22258 57146
rect 26950 57094 27002 57146
rect 27014 57094 27066 57146
rect 27078 57094 27130 57146
rect 27142 57094 27194 57146
rect 27206 57094 27258 57146
rect 31950 57094 32002 57146
rect 32014 57094 32066 57146
rect 32078 57094 32130 57146
rect 32142 57094 32194 57146
rect 32206 57094 32258 57146
rect 36950 57094 37002 57146
rect 37014 57094 37066 57146
rect 37078 57094 37130 57146
rect 37142 57094 37194 57146
rect 37206 57094 37258 57146
rect 41950 57094 42002 57146
rect 42014 57094 42066 57146
rect 42078 57094 42130 57146
rect 42142 57094 42194 57146
rect 42206 57094 42258 57146
rect 46950 57094 47002 57146
rect 47014 57094 47066 57146
rect 47078 57094 47130 57146
rect 47142 57094 47194 57146
rect 47206 57094 47258 57146
rect 51950 57094 52002 57146
rect 52014 57094 52066 57146
rect 52078 57094 52130 57146
rect 52142 57094 52194 57146
rect 52206 57094 52258 57146
rect 56950 57094 57002 57146
rect 57014 57094 57066 57146
rect 57078 57094 57130 57146
rect 57142 57094 57194 57146
rect 57206 57094 57258 57146
rect 2610 56550 2662 56602
rect 2674 56550 2726 56602
rect 2738 56550 2790 56602
rect 2802 56550 2854 56602
rect 2866 56550 2918 56602
rect 7610 56550 7662 56602
rect 7674 56550 7726 56602
rect 7738 56550 7790 56602
rect 7802 56550 7854 56602
rect 7866 56550 7918 56602
rect 12610 56550 12662 56602
rect 12674 56550 12726 56602
rect 12738 56550 12790 56602
rect 12802 56550 12854 56602
rect 12866 56550 12918 56602
rect 17610 56550 17662 56602
rect 17674 56550 17726 56602
rect 17738 56550 17790 56602
rect 17802 56550 17854 56602
rect 17866 56550 17918 56602
rect 22610 56550 22662 56602
rect 22674 56550 22726 56602
rect 22738 56550 22790 56602
rect 22802 56550 22854 56602
rect 22866 56550 22918 56602
rect 27610 56550 27662 56602
rect 27674 56550 27726 56602
rect 27738 56550 27790 56602
rect 27802 56550 27854 56602
rect 27866 56550 27918 56602
rect 32610 56550 32662 56602
rect 32674 56550 32726 56602
rect 32738 56550 32790 56602
rect 32802 56550 32854 56602
rect 32866 56550 32918 56602
rect 37610 56550 37662 56602
rect 37674 56550 37726 56602
rect 37738 56550 37790 56602
rect 37802 56550 37854 56602
rect 37866 56550 37918 56602
rect 42610 56550 42662 56602
rect 42674 56550 42726 56602
rect 42738 56550 42790 56602
rect 42802 56550 42854 56602
rect 42866 56550 42918 56602
rect 47610 56550 47662 56602
rect 47674 56550 47726 56602
rect 47738 56550 47790 56602
rect 47802 56550 47854 56602
rect 47866 56550 47918 56602
rect 52610 56550 52662 56602
rect 52674 56550 52726 56602
rect 52738 56550 52790 56602
rect 52802 56550 52854 56602
rect 52866 56550 52918 56602
rect 57610 56550 57662 56602
rect 57674 56550 57726 56602
rect 57738 56550 57790 56602
rect 57802 56550 57854 56602
rect 57866 56550 57918 56602
rect 1950 56006 2002 56058
rect 2014 56006 2066 56058
rect 2078 56006 2130 56058
rect 2142 56006 2194 56058
rect 2206 56006 2258 56058
rect 6950 56006 7002 56058
rect 7014 56006 7066 56058
rect 7078 56006 7130 56058
rect 7142 56006 7194 56058
rect 7206 56006 7258 56058
rect 11950 56006 12002 56058
rect 12014 56006 12066 56058
rect 12078 56006 12130 56058
rect 12142 56006 12194 56058
rect 12206 56006 12258 56058
rect 16950 56006 17002 56058
rect 17014 56006 17066 56058
rect 17078 56006 17130 56058
rect 17142 56006 17194 56058
rect 17206 56006 17258 56058
rect 21950 56006 22002 56058
rect 22014 56006 22066 56058
rect 22078 56006 22130 56058
rect 22142 56006 22194 56058
rect 22206 56006 22258 56058
rect 26950 56006 27002 56058
rect 27014 56006 27066 56058
rect 27078 56006 27130 56058
rect 27142 56006 27194 56058
rect 27206 56006 27258 56058
rect 31950 56006 32002 56058
rect 32014 56006 32066 56058
rect 32078 56006 32130 56058
rect 32142 56006 32194 56058
rect 32206 56006 32258 56058
rect 36950 56006 37002 56058
rect 37014 56006 37066 56058
rect 37078 56006 37130 56058
rect 37142 56006 37194 56058
rect 37206 56006 37258 56058
rect 41950 56006 42002 56058
rect 42014 56006 42066 56058
rect 42078 56006 42130 56058
rect 42142 56006 42194 56058
rect 42206 56006 42258 56058
rect 46950 56006 47002 56058
rect 47014 56006 47066 56058
rect 47078 56006 47130 56058
rect 47142 56006 47194 56058
rect 47206 56006 47258 56058
rect 51950 56006 52002 56058
rect 52014 56006 52066 56058
rect 52078 56006 52130 56058
rect 52142 56006 52194 56058
rect 52206 56006 52258 56058
rect 56950 56006 57002 56058
rect 57014 56006 57066 56058
rect 57078 56006 57130 56058
rect 57142 56006 57194 56058
rect 57206 56006 57258 56058
rect 58532 55743 58584 55752
rect 58532 55709 58541 55743
rect 58541 55709 58575 55743
rect 58575 55709 58584 55743
rect 58532 55700 58584 55709
rect 2610 55462 2662 55514
rect 2674 55462 2726 55514
rect 2738 55462 2790 55514
rect 2802 55462 2854 55514
rect 2866 55462 2918 55514
rect 7610 55462 7662 55514
rect 7674 55462 7726 55514
rect 7738 55462 7790 55514
rect 7802 55462 7854 55514
rect 7866 55462 7918 55514
rect 12610 55462 12662 55514
rect 12674 55462 12726 55514
rect 12738 55462 12790 55514
rect 12802 55462 12854 55514
rect 12866 55462 12918 55514
rect 17610 55462 17662 55514
rect 17674 55462 17726 55514
rect 17738 55462 17790 55514
rect 17802 55462 17854 55514
rect 17866 55462 17918 55514
rect 22610 55462 22662 55514
rect 22674 55462 22726 55514
rect 22738 55462 22790 55514
rect 22802 55462 22854 55514
rect 22866 55462 22918 55514
rect 27610 55462 27662 55514
rect 27674 55462 27726 55514
rect 27738 55462 27790 55514
rect 27802 55462 27854 55514
rect 27866 55462 27918 55514
rect 32610 55462 32662 55514
rect 32674 55462 32726 55514
rect 32738 55462 32790 55514
rect 32802 55462 32854 55514
rect 32866 55462 32918 55514
rect 37610 55462 37662 55514
rect 37674 55462 37726 55514
rect 37738 55462 37790 55514
rect 37802 55462 37854 55514
rect 37866 55462 37918 55514
rect 42610 55462 42662 55514
rect 42674 55462 42726 55514
rect 42738 55462 42790 55514
rect 42802 55462 42854 55514
rect 42866 55462 42918 55514
rect 47610 55462 47662 55514
rect 47674 55462 47726 55514
rect 47738 55462 47790 55514
rect 47802 55462 47854 55514
rect 47866 55462 47918 55514
rect 52610 55462 52662 55514
rect 52674 55462 52726 55514
rect 52738 55462 52790 55514
rect 52802 55462 52854 55514
rect 52866 55462 52918 55514
rect 57610 55462 57662 55514
rect 57674 55462 57726 55514
rect 57738 55462 57790 55514
rect 57802 55462 57854 55514
rect 57866 55462 57918 55514
rect 58532 55063 58584 55072
rect 58532 55029 58541 55063
rect 58541 55029 58575 55063
rect 58575 55029 58584 55063
rect 58532 55020 58584 55029
rect 1950 54918 2002 54970
rect 2014 54918 2066 54970
rect 2078 54918 2130 54970
rect 2142 54918 2194 54970
rect 2206 54918 2258 54970
rect 6950 54918 7002 54970
rect 7014 54918 7066 54970
rect 7078 54918 7130 54970
rect 7142 54918 7194 54970
rect 7206 54918 7258 54970
rect 11950 54918 12002 54970
rect 12014 54918 12066 54970
rect 12078 54918 12130 54970
rect 12142 54918 12194 54970
rect 12206 54918 12258 54970
rect 16950 54918 17002 54970
rect 17014 54918 17066 54970
rect 17078 54918 17130 54970
rect 17142 54918 17194 54970
rect 17206 54918 17258 54970
rect 21950 54918 22002 54970
rect 22014 54918 22066 54970
rect 22078 54918 22130 54970
rect 22142 54918 22194 54970
rect 22206 54918 22258 54970
rect 26950 54918 27002 54970
rect 27014 54918 27066 54970
rect 27078 54918 27130 54970
rect 27142 54918 27194 54970
rect 27206 54918 27258 54970
rect 31950 54918 32002 54970
rect 32014 54918 32066 54970
rect 32078 54918 32130 54970
rect 32142 54918 32194 54970
rect 32206 54918 32258 54970
rect 36950 54918 37002 54970
rect 37014 54918 37066 54970
rect 37078 54918 37130 54970
rect 37142 54918 37194 54970
rect 37206 54918 37258 54970
rect 41950 54918 42002 54970
rect 42014 54918 42066 54970
rect 42078 54918 42130 54970
rect 42142 54918 42194 54970
rect 42206 54918 42258 54970
rect 46950 54918 47002 54970
rect 47014 54918 47066 54970
rect 47078 54918 47130 54970
rect 47142 54918 47194 54970
rect 47206 54918 47258 54970
rect 51950 54918 52002 54970
rect 52014 54918 52066 54970
rect 52078 54918 52130 54970
rect 52142 54918 52194 54970
rect 52206 54918 52258 54970
rect 56950 54918 57002 54970
rect 57014 54918 57066 54970
rect 57078 54918 57130 54970
rect 57142 54918 57194 54970
rect 57206 54918 57258 54970
rect 2610 54374 2662 54426
rect 2674 54374 2726 54426
rect 2738 54374 2790 54426
rect 2802 54374 2854 54426
rect 2866 54374 2918 54426
rect 7610 54374 7662 54426
rect 7674 54374 7726 54426
rect 7738 54374 7790 54426
rect 7802 54374 7854 54426
rect 7866 54374 7918 54426
rect 12610 54374 12662 54426
rect 12674 54374 12726 54426
rect 12738 54374 12790 54426
rect 12802 54374 12854 54426
rect 12866 54374 12918 54426
rect 17610 54374 17662 54426
rect 17674 54374 17726 54426
rect 17738 54374 17790 54426
rect 17802 54374 17854 54426
rect 17866 54374 17918 54426
rect 22610 54374 22662 54426
rect 22674 54374 22726 54426
rect 22738 54374 22790 54426
rect 22802 54374 22854 54426
rect 22866 54374 22918 54426
rect 27610 54374 27662 54426
rect 27674 54374 27726 54426
rect 27738 54374 27790 54426
rect 27802 54374 27854 54426
rect 27866 54374 27918 54426
rect 32610 54374 32662 54426
rect 32674 54374 32726 54426
rect 32738 54374 32790 54426
rect 32802 54374 32854 54426
rect 32866 54374 32918 54426
rect 37610 54374 37662 54426
rect 37674 54374 37726 54426
rect 37738 54374 37790 54426
rect 37802 54374 37854 54426
rect 37866 54374 37918 54426
rect 42610 54374 42662 54426
rect 42674 54374 42726 54426
rect 42738 54374 42790 54426
rect 42802 54374 42854 54426
rect 42866 54374 42918 54426
rect 47610 54374 47662 54426
rect 47674 54374 47726 54426
rect 47738 54374 47790 54426
rect 47802 54374 47854 54426
rect 47866 54374 47918 54426
rect 52610 54374 52662 54426
rect 52674 54374 52726 54426
rect 52738 54374 52790 54426
rect 52802 54374 52854 54426
rect 52866 54374 52918 54426
rect 57610 54374 57662 54426
rect 57674 54374 57726 54426
rect 57738 54374 57790 54426
rect 57802 54374 57854 54426
rect 57866 54374 57918 54426
rect 58532 53975 58584 53984
rect 58532 53941 58541 53975
rect 58541 53941 58575 53975
rect 58575 53941 58584 53975
rect 58532 53932 58584 53941
rect 1950 53830 2002 53882
rect 2014 53830 2066 53882
rect 2078 53830 2130 53882
rect 2142 53830 2194 53882
rect 2206 53830 2258 53882
rect 6950 53830 7002 53882
rect 7014 53830 7066 53882
rect 7078 53830 7130 53882
rect 7142 53830 7194 53882
rect 7206 53830 7258 53882
rect 11950 53830 12002 53882
rect 12014 53830 12066 53882
rect 12078 53830 12130 53882
rect 12142 53830 12194 53882
rect 12206 53830 12258 53882
rect 16950 53830 17002 53882
rect 17014 53830 17066 53882
rect 17078 53830 17130 53882
rect 17142 53830 17194 53882
rect 17206 53830 17258 53882
rect 21950 53830 22002 53882
rect 22014 53830 22066 53882
rect 22078 53830 22130 53882
rect 22142 53830 22194 53882
rect 22206 53830 22258 53882
rect 26950 53830 27002 53882
rect 27014 53830 27066 53882
rect 27078 53830 27130 53882
rect 27142 53830 27194 53882
rect 27206 53830 27258 53882
rect 31950 53830 32002 53882
rect 32014 53830 32066 53882
rect 32078 53830 32130 53882
rect 32142 53830 32194 53882
rect 32206 53830 32258 53882
rect 36950 53830 37002 53882
rect 37014 53830 37066 53882
rect 37078 53830 37130 53882
rect 37142 53830 37194 53882
rect 37206 53830 37258 53882
rect 41950 53830 42002 53882
rect 42014 53830 42066 53882
rect 42078 53830 42130 53882
rect 42142 53830 42194 53882
rect 42206 53830 42258 53882
rect 46950 53830 47002 53882
rect 47014 53830 47066 53882
rect 47078 53830 47130 53882
rect 47142 53830 47194 53882
rect 47206 53830 47258 53882
rect 51950 53830 52002 53882
rect 52014 53830 52066 53882
rect 52078 53830 52130 53882
rect 52142 53830 52194 53882
rect 52206 53830 52258 53882
rect 56950 53830 57002 53882
rect 57014 53830 57066 53882
rect 57078 53830 57130 53882
rect 57142 53830 57194 53882
rect 57206 53830 57258 53882
rect 58532 53567 58584 53576
rect 58532 53533 58541 53567
rect 58541 53533 58575 53567
rect 58575 53533 58584 53567
rect 58532 53524 58584 53533
rect 2610 53286 2662 53338
rect 2674 53286 2726 53338
rect 2738 53286 2790 53338
rect 2802 53286 2854 53338
rect 2866 53286 2918 53338
rect 7610 53286 7662 53338
rect 7674 53286 7726 53338
rect 7738 53286 7790 53338
rect 7802 53286 7854 53338
rect 7866 53286 7918 53338
rect 12610 53286 12662 53338
rect 12674 53286 12726 53338
rect 12738 53286 12790 53338
rect 12802 53286 12854 53338
rect 12866 53286 12918 53338
rect 17610 53286 17662 53338
rect 17674 53286 17726 53338
rect 17738 53286 17790 53338
rect 17802 53286 17854 53338
rect 17866 53286 17918 53338
rect 22610 53286 22662 53338
rect 22674 53286 22726 53338
rect 22738 53286 22790 53338
rect 22802 53286 22854 53338
rect 22866 53286 22918 53338
rect 27610 53286 27662 53338
rect 27674 53286 27726 53338
rect 27738 53286 27790 53338
rect 27802 53286 27854 53338
rect 27866 53286 27918 53338
rect 32610 53286 32662 53338
rect 32674 53286 32726 53338
rect 32738 53286 32790 53338
rect 32802 53286 32854 53338
rect 32866 53286 32918 53338
rect 37610 53286 37662 53338
rect 37674 53286 37726 53338
rect 37738 53286 37790 53338
rect 37802 53286 37854 53338
rect 37866 53286 37918 53338
rect 42610 53286 42662 53338
rect 42674 53286 42726 53338
rect 42738 53286 42790 53338
rect 42802 53286 42854 53338
rect 42866 53286 42918 53338
rect 47610 53286 47662 53338
rect 47674 53286 47726 53338
rect 47738 53286 47790 53338
rect 47802 53286 47854 53338
rect 47866 53286 47918 53338
rect 52610 53286 52662 53338
rect 52674 53286 52726 53338
rect 52738 53286 52790 53338
rect 52802 53286 52854 53338
rect 52866 53286 52918 53338
rect 57610 53286 57662 53338
rect 57674 53286 57726 53338
rect 57738 53286 57790 53338
rect 57802 53286 57854 53338
rect 57866 53286 57918 53338
rect 1950 52742 2002 52794
rect 2014 52742 2066 52794
rect 2078 52742 2130 52794
rect 2142 52742 2194 52794
rect 2206 52742 2258 52794
rect 6950 52742 7002 52794
rect 7014 52742 7066 52794
rect 7078 52742 7130 52794
rect 7142 52742 7194 52794
rect 7206 52742 7258 52794
rect 11950 52742 12002 52794
rect 12014 52742 12066 52794
rect 12078 52742 12130 52794
rect 12142 52742 12194 52794
rect 12206 52742 12258 52794
rect 16950 52742 17002 52794
rect 17014 52742 17066 52794
rect 17078 52742 17130 52794
rect 17142 52742 17194 52794
rect 17206 52742 17258 52794
rect 21950 52742 22002 52794
rect 22014 52742 22066 52794
rect 22078 52742 22130 52794
rect 22142 52742 22194 52794
rect 22206 52742 22258 52794
rect 26950 52742 27002 52794
rect 27014 52742 27066 52794
rect 27078 52742 27130 52794
rect 27142 52742 27194 52794
rect 27206 52742 27258 52794
rect 31950 52742 32002 52794
rect 32014 52742 32066 52794
rect 32078 52742 32130 52794
rect 32142 52742 32194 52794
rect 32206 52742 32258 52794
rect 36950 52742 37002 52794
rect 37014 52742 37066 52794
rect 37078 52742 37130 52794
rect 37142 52742 37194 52794
rect 37206 52742 37258 52794
rect 41950 52742 42002 52794
rect 42014 52742 42066 52794
rect 42078 52742 42130 52794
rect 42142 52742 42194 52794
rect 42206 52742 42258 52794
rect 46950 52742 47002 52794
rect 47014 52742 47066 52794
rect 47078 52742 47130 52794
rect 47142 52742 47194 52794
rect 47206 52742 47258 52794
rect 51950 52742 52002 52794
rect 52014 52742 52066 52794
rect 52078 52742 52130 52794
rect 52142 52742 52194 52794
rect 52206 52742 52258 52794
rect 56950 52742 57002 52794
rect 57014 52742 57066 52794
rect 57078 52742 57130 52794
rect 57142 52742 57194 52794
rect 57206 52742 57258 52794
rect 58532 52479 58584 52488
rect 58532 52445 58541 52479
rect 58541 52445 58575 52479
rect 58575 52445 58584 52479
rect 58532 52436 58584 52445
rect 2610 52198 2662 52250
rect 2674 52198 2726 52250
rect 2738 52198 2790 52250
rect 2802 52198 2854 52250
rect 2866 52198 2918 52250
rect 7610 52198 7662 52250
rect 7674 52198 7726 52250
rect 7738 52198 7790 52250
rect 7802 52198 7854 52250
rect 7866 52198 7918 52250
rect 12610 52198 12662 52250
rect 12674 52198 12726 52250
rect 12738 52198 12790 52250
rect 12802 52198 12854 52250
rect 12866 52198 12918 52250
rect 17610 52198 17662 52250
rect 17674 52198 17726 52250
rect 17738 52198 17790 52250
rect 17802 52198 17854 52250
rect 17866 52198 17918 52250
rect 22610 52198 22662 52250
rect 22674 52198 22726 52250
rect 22738 52198 22790 52250
rect 22802 52198 22854 52250
rect 22866 52198 22918 52250
rect 27610 52198 27662 52250
rect 27674 52198 27726 52250
rect 27738 52198 27790 52250
rect 27802 52198 27854 52250
rect 27866 52198 27918 52250
rect 32610 52198 32662 52250
rect 32674 52198 32726 52250
rect 32738 52198 32790 52250
rect 32802 52198 32854 52250
rect 32866 52198 32918 52250
rect 37610 52198 37662 52250
rect 37674 52198 37726 52250
rect 37738 52198 37790 52250
rect 37802 52198 37854 52250
rect 37866 52198 37918 52250
rect 42610 52198 42662 52250
rect 42674 52198 42726 52250
rect 42738 52198 42790 52250
rect 42802 52198 42854 52250
rect 42866 52198 42918 52250
rect 47610 52198 47662 52250
rect 47674 52198 47726 52250
rect 47738 52198 47790 52250
rect 47802 52198 47854 52250
rect 47866 52198 47918 52250
rect 52610 52198 52662 52250
rect 52674 52198 52726 52250
rect 52738 52198 52790 52250
rect 52802 52198 52854 52250
rect 52866 52198 52918 52250
rect 57610 52198 57662 52250
rect 57674 52198 57726 52250
rect 57738 52198 57790 52250
rect 57802 52198 57854 52250
rect 57866 52198 57918 52250
rect 58532 51799 58584 51808
rect 58532 51765 58541 51799
rect 58541 51765 58575 51799
rect 58575 51765 58584 51799
rect 58532 51756 58584 51765
rect 1950 51654 2002 51706
rect 2014 51654 2066 51706
rect 2078 51654 2130 51706
rect 2142 51654 2194 51706
rect 2206 51654 2258 51706
rect 6950 51654 7002 51706
rect 7014 51654 7066 51706
rect 7078 51654 7130 51706
rect 7142 51654 7194 51706
rect 7206 51654 7258 51706
rect 11950 51654 12002 51706
rect 12014 51654 12066 51706
rect 12078 51654 12130 51706
rect 12142 51654 12194 51706
rect 12206 51654 12258 51706
rect 16950 51654 17002 51706
rect 17014 51654 17066 51706
rect 17078 51654 17130 51706
rect 17142 51654 17194 51706
rect 17206 51654 17258 51706
rect 21950 51654 22002 51706
rect 22014 51654 22066 51706
rect 22078 51654 22130 51706
rect 22142 51654 22194 51706
rect 22206 51654 22258 51706
rect 26950 51654 27002 51706
rect 27014 51654 27066 51706
rect 27078 51654 27130 51706
rect 27142 51654 27194 51706
rect 27206 51654 27258 51706
rect 31950 51654 32002 51706
rect 32014 51654 32066 51706
rect 32078 51654 32130 51706
rect 32142 51654 32194 51706
rect 32206 51654 32258 51706
rect 36950 51654 37002 51706
rect 37014 51654 37066 51706
rect 37078 51654 37130 51706
rect 37142 51654 37194 51706
rect 37206 51654 37258 51706
rect 41950 51654 42002 51706
rect 42014 51654 42066 51706
rect 42078 51654 42130 51706
rect 42142 51654 42194 51706
rect 42206 51654 42258 51706
rect 46950 51654 47002 51706
rect 47014 51654 47066 51706
rect 47078 51654 47130 51706
rect 47142 51654 47194 51706
rect 47206 51654 47258 51706
rect 51950 51654 52002 51706
rect 52014 51654 52066 51706
rect 52078 51654 52130 51706
rect 52142 51654 52194 51706
rect 52206 51654 52258 51706
rect 56950 51654 57002 51706
rect 57014 51654 57066 51706
rect 57078 51654 57130 51706
rect 57142 51654 57194 51706
rect 57206 51654 57258 51706
rect 2610 51110 2662 51162
rect 2674 51110 2726 51162
rect 2738 51110 2790 51162
rect 2802 51110 2854 51162
rect 2866 51110 2918 51162
rect 7610 51110 7662 51162
rect 7674 51110 7726 51162
rect 7738 51110 7790 51162
rect 7802 51110 7854 51162
rect 7866 51110 7918 51162
rect 12610 51110 12662 51162
rect 12674 51110 12726 51162
rect 12738 51110 12790 51162
rect 12802 51110 12854 51162
rect 12866 51110 12918 51162
rect 17610 51110 17662 51162
rect 17674 51110 17726 51162
rect 17738 51110 17790 51162
rect 17802 51110 17854 51162
rect 17866 51110 17918 51162
rect 22610 51110 22662 51162
rect 22674 51110 22726 51162
rect 22738 51110 22790 51162
rect 22802 51110 22854 51162
rect 22866 51110 22918 51162
rect 27610 51110 27662 51162
rect 27674 51110 27726 51162
rect 27738 51110 27790 51162
rect 27802 51110 27854 51162
rect 27866 51110 27918 51162
rect 32610 51110 32662 51162
rect 32674 51110 32726 51162
rect 32738 51110 32790 51162
rect 32802 51110 32854 51162
rect 32866 51110 32918 51162
rect 37610 51110 37662 51162
rect 37674 51110 37726 51162
rect 37738 51110 37790 51162
rect 37802 51110 37854 51162
rect 37866 51110 37918 51162
rect 42610 51110 42662 51162
rect 42674 51110 42726 51162
rect 42738 51110 42790 51162
rect 42802 51110 42854 51162
rect 42866 51110 42918 51162
rect 47610 51110 47662 51162
rect 47674 51110 47726 51162
rect 47738 51110 47790 51162
rect 47802 51110 47854 51162
rect 47866 51110 47918 51162
rect 52610 51110 52662 51162
rect 52674 51110 52726 51162
rect 52738 51110 52790 51162
rect 52802 51110 52854 51162
rect 52866 51110 52918 51162
rect 57610 51110 57662 51162
rect 57674 51110 57726 51162
rect 57738 51110 57790 51162
rect 57802 51110 57854 51162
rect 57866 51110 57918 51162
rect 58532 50711 58584 50720
rect 58532 50677 58541 50711
rect 58541 50677 58575 50711
rect 58575 50677 58584 50711
rect 58532 50668 58584 50677
rect 1950 50566 2002 50618
rect 2014 50566 2066 50618
rect 2078 50566 2130 50618
rect 2142 50566 2194 50618
rect 2206 50566 2258 50618
rect 6950 50566 7002 50618
rect 7014 50566 7066 50618
rect 7078 50566 7130 50618
rect 7142 50566 7194 50618
rect 7206 50566 7258 50618
rect 11950 50566 12002 50618
rect 12014 50566 12066 50618
rect 12078 50566 12130 50618
rect 12142 50566 12194 50618
rect 12206 50566 12258 50618
rect 16950 50566 17002 50618
rect 17014 50566 17066 50618
rect 17078 50566 17130 50618
rect 17142 50566 17194 50618
rect 17206 50566 17258 50618
rect 21950 50566 22002 50618
rect 22014 50566 22066 50618
rect 22078 50566 22130 50618
rect 22142 50566 22194 50618
rect 22206 50566 22258 50618
rect 26950 50566 27002 50618
rect 27014 50566 27066 50618
rect 27078 50566 27130 50618
rect 27142 50566 27194 50618
rect 27206 50566 27258 50618
rect 31950 50566 32002 50618
rect 32014 50566 32066 50618
rect 32078 50566 32130 50618
rect 32142 50566 32194 50618
rect 32206 50566 32258 50618
rect 36950 50566 37002 50618
rect 37014 50566 37066 50618
rect 37078 50566 37130 50618
rect 37142 50566 37194 50618
rect 37206 50566 37258 50618
rect 41950 50566 42002 50618
rect 42014 50566 42066 50618
rect 42078 50566 42130 50618
rect 42142 50566 42194 50618
rect 42206 50566 42258 50618
rect 46950 50566 47002 50618
rect 47014 50566 47066 50618
rect 47078 50566 47130 50618
rect 47142 50566 47194 50618
rect 47206 50566 47258 50618
rect 51950 50566 52002 50618
rect 52014 50566 52066 50618
rect 52078 50566 52130 50618
rect 52142 50566 52194 50618
rect 52206 50566 52258 50618
rect 56950 50566 57002 50618
rect 57014 50566 57066 50618
rect 57078 50566 57130 50618
rect 57142 50566 57194 50618
rect 57206 50566 57258 50618
rect 58532 50303 58584 50312
rect 58532 50269 58541 50303
rect 58541 50269 58575 50303
rect 58575 50269 58584 50303
rect 58532 50260 58584 50269
rect 2610 50022 2662 50074
rect 2674 50022 2726 50074
rect 2738 50022 2790 50074
rect 2802 50022 2854 50074
rect 2866 50022 2918 50074
rect 7610 50022 7662 50074
rect 7674 50022 7726 50074
rect 7738 50022 7790 50074
rect 7802 50022 7854 50074
rect 7866 50022 7918 50074
rect 12610 50022 12662 50074
rect 12674 50022 12726 50074
rect 12738 50022 12790 50074
rect 12802 50022 12854 50074
rect 12866 50022 12918 50074
rect 17610 50022 17662 50074
rect 17674 50022 17726 50074
rect 17738 50022 17790 50074
rect 17802 50022 17854 50074
rect 17866 50022 17918 50074
rect 22610 50022 22662 50074
rect 22674 50022 22726 50074
rect 22738 50022 22790 50074
rect 22802 50022 22854 50074
rect 22866 50022 22918 50074
rect 27610 50022 27662 50074
rect 27674 50022 27726 50074
rect 27738 50022 27790 50074
rect 27802 50022 27854 50074
rect 27866 50022 27918 50074
rect 32610 50022 32662 50074
rect 32674 50022 32726 50074
rect 32738 50022 32790 50074
rect 32802 50022 32854 50074
rect 32866 50022 32918 50074
rect 37610 50022 37662 50074
rect 37674 50022 37726 50074
rect 37738 50022 37790 50074
rect 37802 50022 37854 50074
rect 37866 50022 37918 50074
rect 42610 50022 42662 50074
rect 42674 50022 42726 50074
rect 42738 50022 42790 50074
rect 42802 50022 42854 50074
rect 42866 50022 42918 50074
rect 47610 50022 47662 50074
rect 47674 50022 47726 50074
rect 47738 50022 47790 50074
rect 47802 50022 47854 50074
rect 47866 50022 47918 50074
rect 52610 50022 52662 50074
rect 52674 50022 52726 50074
rect 52738 50022 52790 50074
rect 52802 50022 52854 50074
rect 52866 50022 52918 50074
rect 57610 50022 57662 50074
rect 57674 50022 57726 50074
rect 57738 50022 57790 50074
rect 57802 50022 57854 50074
rect 57866 50022 57918 50074
rect 1950 49478 2002 49530
rect 2014 49478 2066 49530
rect 2078 49478 2130 49530
rect 2142 49478 2194 49530
rect 2206 49478 2258 49530
rect 6950 49478 7002 49530
rect 7014 49478 7066 49530
rect 7078 49478 7130 49530
rect 7142 49478 7194 49530
rect 7206 49478 7258 49530
rect 11950 49478 12002 49530
rect 12014 49478 12066 49530
rect 12078 49478 12130 49530
rect 12142 49478 12194 49530
rect 12206 49478 12258 49530
rect 16950 49478 17002 49530
rect 17014 49478 17066 49530
rect 17078 49478 17130 49530
rect 17142 49478 17194 49530
rect 17206 49478 17258 49530
rect 21950 49478 22002 49530
rect 22014 49478 22066 49530
rect 22078 49478 22130 49530
rect 22142 49478 22194 49530
rect 22206 49478 22258 49530
rect 26950 49478 27002 49530
rect 27014 49478 27066 49530
rect 27078 49478 27130 49530
rect 27142 49478 27194 49530
rect 27206 49478 27258 49530
rect 31950 49478 32002 49530
rect 32014 49478 32066 49530
rect 32078 49478 32130 49530
rect 32142 49478 32194 49530
rect 32206 49478 32258 49530
rect 36950 49478 37002 49530
rect 37014 49478 37066 49530
rect 37078 49478 37130 49530
rect 37142 49478 37194 49530
rect 37206 49478 37258 49530
rect 41950 49478 42002 49530
rect 42014 49478 42066 49530
rect 42078 49478 42130 49530
rect 42142 49478 42194 49530
rect 42206 49478 42258 49530
rect 46950 49478 47002 49530
rect 47014 49478 47066 49530
rect 47078 49478 47130 49530
rect 47142 49478 47194 49530
rect 47206 49478 47258 49530
rect 51950 49478 52002 49530
rect 52014 49478 52066 49530
rect 52078 49478 52130 49530
rect 52142 49478 52194 49530
rect 52206 49478 52258 49530
rect 56950 49478 57002 49530
rect 57014 49478 57066 49530
rect 57078 49478 57130 49530
rect 57142 49478 57194 49530
rect 57206 49478 57258 49530
rect 58532 49215 58584 49224
rect 58532 49181 58541 49215
rect 58541 49181 58575 49215
rect 58575 49181 58584 49215
rect 58532 49172 58584 49181
rect 2610 48934 2662 48986
rect 2674 48934 2726 48986
rect 2738 48934 2790 48986
rect 2802 48934 2854 48986
rect 2866 48934 2918 48986
rect 7610 48934 7662 48986
rect 7674 48934 7726 48986
rect 7738 48934 7790 48986
rect 7802 48934 7854 48986
rect 7866 48934 7918 48986
rect 12610 48934 12662 48986
rect 12674 48934 12726 48986
rect 12738 48934 12790 48986
rect 12802 48934 12854 48986
rect 12866 48934 12918 48986
rect 17610 48934 17662 48986
rect 17674 48934 17726 48986
rect 17738 48934 17790 48986
rect 17802 48934 17854 48986
rect 17866 48934 17918 48986
rect 22610 48934 22662 48986
rect 22674 48934 22726 48986
rect 22738 48934 22790 48986
rect 22802 48934 22854 48986
rect 22866 48934 22918 48986
rect 27610 48934 27662 48986
rect 27674 48934 27726 48986
rect 27738 48934 27790 48986
rect 27802 48934 27854 48986
rect 27866 48934 27918 48986
rect 32610 48934 32662 48986
rect 32674 48934 32726 48986
rect 32738 48934 32790 48986
rect 32802 48934 32854 48986
rect 32866 48934 32918 48986
rect 37610 48934 37662 48986
rect 37674 48934 37726 48986
rect 37738 48934 37790 48986
rect 37802 48934 37854 48986
rect 37866 48934 37918 48986
rect 42610 48934 42662 48986
rect 42674 48934 42726 48986
rect 42738 48934 42790 48986
rect 42802 48934 42854 48986
rect 42866 48934 42918 48986
rect 47610 48934 47662 48986
rect 47674 48934 47726 48986
rect 47738 48934 47790 48986
rect 47802 48934 47854 48986
rect 47866 48934 47918 48986
rect 52610 48934 52662 48986
rect 52674 48934 52726 48986
rect 52738 48934 52790 48986
rect 52802 48934 52854 48986
rect 52866 48934 52918 48986
rect 57610 48934 57662 48986
rect 57674 48934 57726 48986
rect 57738 48934 57790 48986
rect 57802 48934 57854 48986
rect 57866 48934 57918 48986
rect 58532 48535 58584 48544
rect 58532 48501 58541 48535
rect 58541 48501 58575 48535
rect 58575 48501 58584 48535
rect 58532 48492 58584 48501
rect 1950 48390 2002 48442
rect 2014 48390 2066 48442
rect 2078 48390 2130 48442
rect 2142 48390 2194 48442
rect 2206 48390 2258 48442
rect 6950 48390 7002 48442
rect 7014 48390 7066 48442
rect 7078 48390 7130 48442
rect 7142 48390 7194 48442
rect 7206 48390 7258 48442
rect 11950 48390 12002 48442
rect 12014 48390 12066 48442
rect 12078 48390 12130 48442
rect 12142 48390 12194 48442
rect 12206 48390 12258 48442
rect 16950 48390 17002 48442
rect 17014 48390 17066 48442
rect 17078 48390 17130 48442
rect 17142 48390 17194 48442
rect 17206 48390 17258 48442
rect 21950 48390 22002 48442
rect 22014 48390 22066 48442
rect 22078 48390 22130 48442
rect 22142 48390 22194 48442
rect 22206 48390 22258 48442
rect 26950 48390 27002 48442
rect 27014 48390 27066 48442
rect 27078 48390 27130 48442
rect 27142 48390 27194 48442
rect 27206 48390 27258 48442
rect 31950 48390 32002 48442
rect 32014 48390 32066 48442
rect 32078 48390 32130 48442
rect 32142 48390 32194 48442
rect 32206 48390 32258 48442
rect 36950 48390 37002 48442
rect 37014 48390 37066 48442
rect 37078 48390 37130 48442
rect 37142 48390 37194 48442
rect 37206 48390 37258 48442
rect 41950 48390 42002 48442
rect 42014 48390 42066 48442
rect 42078 48390 42130 48442
rect 42142 48390 42194 48442
rect 42206 48390 42258 48442
rect 46950 48390 47002 48442
rect 47014 48390 47066 48442
rect 47078 48390 47130 48442
rect 47142 48390 47194 48442
rect 47206 48390 47258 48442
rect 51950 48390 52002 48442
rect 52014 48390 52066 48442
rect 52078 48390 52130 48442
rect 52142 48390 52194 48442
rect 52206 48390 52258 48442
rect 56950 48390 57002 48442
rect 57014 48390 57066 48442
rect 57078 48390 57130 48442
rect 57142 48390 57194 48442
rect 57206 48390 57258 48442
rect 2610 47846 2662 47898
rect 2674 47846 2726 47898
rect 2738 47846 2790 47898
rect 2802 47846 2854 47898
rect 2866 47846 2918 47898
rect 7610 47846 7662 47898
rect 7674 47846 7726 47898
rect 7738 47846 7790 47898
rect 7802 47846 7854 47898
rect 7866 47846 7918 47898
rect 12610 47846 12662 47898
rect 12674 47846 12726 47898
rect 12738 47846 12790 47898
rect 12802 47846 12854 47898
rect 12866 47846 12918 47898
rect 17610 47846 17662 47898
rect 17674 47846 17726 47898
rect 17738 47846 17790 47898
rect 17802 47846 17854 47898
rect 17866 47846 17918 47898
rect 22610 47846 22662 47898
rect 22674 47846 22726 47898
rect 22738 47846 22790 47898
rect 22802 47846 22854 47898
rect 22866 47846 22918 47898
rect 27610 47846 27662 47898
rect 27674 47846 27726 47898
rect 27738 47846 27790 47898
rect 27802 47846 27854 47898
rect 27866 47846 27918 47898
rect 32610 47846 32662 47898
rect 32674 47846 32726 47898
rect 32738 47846 32790 47898
rect 32802 47846 32854 47898
rect 32866 47846 32918 47898
rect 37610 47846 37662 47898
rect 37674 47846 37726 47898
rect 37738 47846 37790 47898
rect 37802 47846 37854 47898
rect 37866 47846 37918 47898
rect 42610 47846 42662 47898
rect 42674 47846 42726 47898
rect 42738 47846 42790 47898
rect 42802 47846 42854 47898
rect 42866 47846 42918 47898
rect 47610 47846 47662 47898
rect 47674 47846 47726 47898
rect 47738 47846 47790 47898
rect 47802 47846 47854 47898
rect 47866 47846 47918 47898
rect 52610 47846 52662 47898
rect 52674 47846 52726 47898
rect 52738 47846 52790 47898
rect 52802 47846 52854 47898
rect 52866 47846 52918 47898
rect 57610 47846 57662 47898
rect 57674 47846 57726 47898
rect 57738 47846 57790 47898
rect 57802 47846 57854 47898
rect 57866 47846 57918 47898
rect 58532 47447 58584 47456
rect 58532 47413 58541 47447
rect 58541 47413 58575 47447
rect 58575 47413 58584 47447
rect 58532 47404 58584 47413
rect 1950 47302 2002 47354
rect 2014 47302 2066 47354
rect 2078 47302 2130 47354
rect 2142 47302 2194 47354
rect 2206 47302 2258 47354
rect 6950 47302 7002 47354
rect 7014 47302 7066 47354
rect 7078 47302 7130 47354
rect 7142 47302 7194 47354
rect 7206 47302 7258 47354
rect 11950 47302 12002 47354
rect 12014 47302 12066 47354
rect 12078 47302 12130 47354
rect 12142 47302 12194 47354
rect 12206 47302 12258 47354
rect 16950 47302 17002 47354
rect 17014 47302 17066 47354
rect 17078 47302 17130 47354
rect 17142 47302 17194 47354
rect 17206 47302 17258 47354
rect 21950 47302 22002 47354
rect 22014 47302 22066 47354
rect 22078 47302 22130 47354
rect 22142 47302 22194 47354
rect 22206 47302 22258 47354
rect 26950 47302 27002 47354
rect 27014 47302 27066 47354
rect 27078 47302 27130 47354
rect 27142 47302 27194 47354
rect 27206 47302 27258 47354
rect 31950 47302 32002 47354
rect 32014 47302 32066 47354
rect 32078 47302 32130 47354
rect 32142 47302 32194 47354
rect 32206 47302 32258 47354
rect 36950 47302 37002 47354
rect 37014 47302 37066 47354
rect 37078 47302 37130 47354
rect 37142 47302 37194 47354
rect 37206 47302 37258 47354
rect 41950 47302 42002 47354
rect 42014 47302 42066 47354
rect 42078 47302 42130 47354
rect 42142 47302 42194 47354
rect 42206 47302 42258 47354
rect 46950 47302 47002 47354
rect 47014 47302 47066 47354
rect 47078 47302 47130 47354
rect 47142 47302 47194 47354
rect 47206 47302 47258 47354
rect 51950 47302 52002 47354
rect 52014 47302 52066 47354
rect 52078 47302 52130 47354
rect 52142 47302 52194 47354
rect 52206 47302 52258 47354
rect 56950 47302 57002 47354
rect 57014 47302 57066 47354
rect 57078 47302 57130 47354
rect 57142 47302 57194 47354
rect 57206 47302 57258 47354
rect 58532 47039 58584 47048
rect 58532 47005 58541 47039
rect 58541 47005 58575 47039
rect 58575 47005 58584 47039
rect 58532 46996 58584 47005
rect 2610 46758 2662 46810
rect 2674 46758 2726 46810
rect 2738 46758 2790 46810
rect 2802 46758 2854 46810
rect 2866 46758 2918 46810
rect 7610 46758 7662 46810
rect 7674 46758 7726 46810
rect 7738 46758 7790 46810
rect 7802 46758 7854 46810
rect 7866 46758 7918 46810
rect 12610 46758 12662 46810
rect 12674 46758 12726 46810
rect 12738 46758 12790 46810
rect 12802 46758 12854 46810
rect 12866 46758 12918 46810
rect 17610 46758 17662 46810
rect 17674 46758 17726 46810
rect 17738 46758 17790 46810
rect 17802 46758 17854 46810
rect 17866 46758 17918 46810
rect 22610 46758 22662 46810
rect 22674 46758 22726 46810
rect 22738 46758 22790 46810
rect 22802 46758 22854 46810
rect 22866 46758 22918 46810
rect 27610 46758 27662 46810
rect 27674 46758 27726 46810
rect 27738 46758 27790 46810
rect 27802 46758 27854 46810
rect 27866 46758 27918 46810
rect 32610 46758 32662 46810
rect 32674 46758 32726 46810
rect 32738 46758 32790 46810
rect 32802 46758 32854 46810
rect 32866 46758 32918 46810
rect 37610 46758 37662 46810
rect 37674 46758 37726 46810
rect 37738 46758 37790 46810
rect 37802 46758 37854 46810
rect 37866 46758 37918 46810
rect 42610 46758 42662 46810
rect 42674 46758 42726 46810
rect 42738 46758 42790 46810
rect 42802 46758 42854 46810
rect 42866 46758 42918 46810
rect 47610 46758 47662 46810
rect 47674 46758 47726 46810
rect 47738 46758 47790 46810
rect 47802 46758 47854 46810
rect 47866 46758 47918 46810
rect 52610 46758 52662 46810
rect 52674 46758 52726 46810
rect 52738 46758 52790 46810
rect 52802 46758 52854 46810
rect 52866 46758 52918 46810
rect 57610 46758 57662 46810
rect 57674 46758 57726 46810
rect 57738 46758 57790 46810
rect 57802 46758 57854 46810
rect 57866 46758 57918 46810
rect 1950 46214 2002 46266
rect 2014 46214 2066 46266
rect 2078 46214 2130 46266
rect 2142 46214 2194 46266
rect 2206 46214 2258 46266
rect 6950 46214 7002 46266
rect 7014 46214 7066 46266
rect 7078 46214 7130 46266
rect 7142 46214 7194 46266
rect 7206 46214 7258 46266
rect 11950 46214 12002 46266
rect 12014 46214 12066 46266
rect 12078 46214 12130 46266
rect 12142 46214 12194 46266
rect 12206 46214 12258 46266
rect 16950 46214 17002 46266
rect 17014 46214 17066 46266
rect 17078 46214 17130 46266
rect 17142 46214 17194 46266
rect 17206 46214 17258 46266
rect 21950 46214 22002 46266
rect 22014 46214 22066 46266
rect 22078 46214 22130 46266
rect 22142 46214 22194 46266
rect 22206 46214 22258 46266
rect 26950 46214 27002 46266
rect 27014 46214 27066 46266
rect 27078 46214 27130 46266
rect 27142 46214 27194 46266
rect 27206 46214 27258 46266
rect 31950 46214 32002 46266
rect 32014 46214 32066 46266
rect 32078 46214 32130 46266
rect 32142 46214 32194 46266
rect 32206 46214 32258 46266
rect 36950 46214 37002 46266
rect 37014 46214 37066 46266
rect 37078 46214 37130 46266
rect 37142 46214 37194 46266
rect 37206 46214 37258 46266
rect 41950 46214 42002 46266
rect 42014 46214 42066 46266
rect 42078 46214 42130 46266
rect 42142 46214 42194 46266
rect 42206 46214 42258 46266
rect 46950 46214 47002 46266
rect 47014 46214 47066 46266
rect 47078 46214 47130 46266
rect 47142 46214 47194 46266
rect 47206 46214 47258 46266
rect 51950 46214 52002 46266
rect 52014 46214 52066 46266
rect 52078 46214 52130 46266
rect 52142 46214 52194 46266
rect 52206 46214 52258 46266
rect 56950 46214 57002 46266
rect 57014 46214 57066 46266
rect 57078 46214 57130 46266
rect 57142 46214 57194 46266
rect 57206 46214 57258 46266
rect 58532 45951 58584 45960
rect 58532 45917 58541 45951
rect 58541 45917 58575 45951
rect 58575 45917 58584 45951
rect 58532 45908 58584 45917
rect 2610 45670 2662 45722
rect 2674 45670 2726 45722
rect 2738 45670 2790 45722
rect 2802 45670 2854 45722
rect 2866 45670 2918 45722
rect 7610 45670 7662 45722
rect 7674 45670 7726 45722
rect 7738 45670 7790 45722
rect 7802 45670 7854 45722
rect 7866 45670 7918 45722
rect 12610 45670 12662 45722
rect 12674 45670 12726 45722
rect 12738 45670 12790 45722
rect 12802 45670 12854 45722
rect 12866 45670 12918 45722
rect 17610 45670 17662 45722
rect 17674 45670 17726 45722
rect 17738 45670 17790 45722
rect 17802 45670 17854 45722
rect 17866 45670 17918 45722
rect 22610 45670 22662 45722
rect 22674 45670 22726 45722
rect 22738 45670 22790 45722
rect 22802 45670 22854 45722
rect 22866 45670 22918 45722
rect 27610 45670 27662 45722
rect 27674 45670 27726 45722
rect 27738 45670 27790 45722
rect 27802 45670 27854 45722
rect 27866 45670 27918 45722
rect 32610 45670 32662 45722
rect 32674 45670 32726 45722
rect 32738 45670 32790 45722
rect 32802 45670 32854 45722
rect 32866 45670 32918 45722
rect 37610 45670 37662 45722
rect 37674 45670 37726 45722
rect 37738 45670 37790 45722
rect 37802 45670 37854 45722
rect 37866 45670 37918 45722
rect 42610 45670 42662 45722
rect 42674 45670 42726 45722
rect 42738 45670 42790 45722
rect 42802 45670 42854 45722
rect 42866 45670 42918 45722
rect 47610 45670 47662 45722
rect 47674 45670 47726 45722
rect 47738 45670 47790 45722
rect 47802 45670 47854 45722
rect 47866 45670 47918 45722
rect 52610 45670 52662 45722
rect 52674 45670 52726 45722
rect 52738 45670 52790 45722
rect 52802 45670 52854 45722
rect 52866 45670 52918 45722
rect 57610 45670 57662 45722
rect 57674 45670 57726 45722
rect 57738 45670 57790 45722
rect 57802 45670 57854 45722
rect 57866 45670 57918 45722
rect 58532 45271 58584 45280
rect 58532 45237 58541 45271
rect 58541 45237 58575 45271
rect 58575 45237 58584 45271
rect 58532 45228 58584 45237
rect 1950 45126 2002 45178
rect 2014 45126 2066 45178
rect 2078 45126 2130 45178
rect 2142 45126 2194 45178
rect 2206 45126 2258 45178
rect 6950 45126 7002 45178
rect 7014 45126 7066 45178
rect 7078 45126 7130 45178
rect 7142 45126 7194 45178
rect 7206 45126 7258 45178
rect 11950 45126 12002 45178
rect 12014 45126 12066 45178
rect 12078 45126 12130 45178
rect 12142 45126 12194 45178
rect 12206 45126 12258 45178
rect 16950 45126 17002 45178
rect 17014 45126 17066 45178
rect 17078 45126 17130 45178
rect 17142 45126 17194 45178
rect 17206 45126 17258 45178
rect 21950 45126 22002 45178
rect 22014 45126 22066 45178
rect 22078 45126 22130 45178
rect 22142 45126 22194 45178
rect 22206 45126 22258 45178
rect 26950 45126 27002 45178
rect 27014 45126 27066 45178
rect 27078 45126 27130 45178
rect 27142 45126 27194 45178
rect 27206 45126 27258 45178
rect 31950 45126 32002 45178
rect 32014 45126 32066 45178
rect 32078 45126 32130 45178
rect 32142 45126 32194 45178
rect 32206 45126 32258 45178
rect 36950 45126 37002 45178
rect 37014 45126 37066 45178
rect 37078 45126 37130 45178
rect 37142 45126 37194 45178
rect 37206 45126 37258 45178
rect 41950 45126 42002 45178
rect 42014 45126 42066 45178
rect 42078 45126 42130 45178
rect 42142 45126 42194 45178
rect 42206 45126 42258 45178
rect 46950 45126 47002 45178
rect 47014 45126 47066 45178
rect 47078 45126 47130 45178
rect 47142 45126 47194 45178
rect 47206 45126 47258 45178
rect 51950 45126 52002 45178
rect 52014 45126 52066 45178
rect 52078 45126 52130 45178
rect 52142 45126 52194 45178
rect 52206 45126 52258 45178
rect 56950 45126 57002 45178
rect 57014 45126 57066 45178
rect 57078 45126 57130 45178
rect 57142 45126 57194 45178
rect 57206 45126 57258 45178
rect 2610 44582 2662 44634
rect 2674 44582 2726 44634
rect 2738 44582 2790 44634
rect 2802 44582 2854 44634
rect 2866 44582 2918 44634
rect 7610 44582 7662 44634
rect 7674 44582 7726 44634
rect 7738 44582 7790 44634
rect 7802 44582 7854 44634
rect 7866 44582 7918 44634
rect 12610 44582 12662 44634
rect 12674 44582 12726 44634
rect 12738 44582 12790 44634
rect 12802 44582 12854 44634
rect 12866 44582 12918 44634
rect 17610 44582 17662 44634
rect 17674 44582 17726 44634
rect 17738 44582 17790 44634
rect 17802 44582 17854 44634
rect 17866 44582 17918 44634
rect 22610 44582 22662 44634
rect 22674 44582 22726 44634
rect 22738 44582 22790 44634
rect 22802 44582 22854 44634
rect 22866 44582 22918 44634
rect 27610 44582 27662 44634
rect 27674 44582 27726 44634
rect 27738 44582 27790 44634
rect 27802 44582 27854 44634
rect 27866 44582 27918 44634
rect 32610 44582 32662 44634
rect 32674 44582 32726 44634
rect 32738 44582 32790 44634
rect 32802 44582 32854 44634
rect 32866 44582 32918 44634
rect 37610 44582 37662 44634
rect 37674 44582 37726 44634
rect 37738 44582 37790 44634
rect 37802 44582 37854 44634
rect 37866 44582 37918 44634
rect 42610 44582 42662 44634
rect 42674 44582 42726 44634
rect 42738 44582 42790 44634
rect 42802 44582 42854 44634
rect 42866 44582 42918 44634
rect 47610 44582 47662 44634
rect 47674 44582 47726 44634
rect 47738 44582 47790 44634
rect 47802 44582 47854 44634
rect 47866 44582 47918 44634
rect 52610 44582 52662 44634
rect 52674 44582 52726 44634
rect 52738 44582 52790 44634
rect 52802 44582 52854 44634
rect 52866 44582 52918 44634
rect 57610 44582 57662 44634
rect 57674 44582 57726 44634
rect 57738 44582 57790 44634
rect 57802 44582 57854 44634
rect 57866 44582 57918 44634
rect 58532 44183 58584 44192
rect 58532 44149 58541 44183
rect 58541 44149 58575 44183
rect 58575 44149 58584 44183
rect 58532 44140 58584 44149
rect 1950 44038 2002 44090
rect 2014 44038 2066 44090
rect 2078 44038 2130 44090
rect 2142 44038 2194 44090
rect 2206 44038 2258 44090
rect 6950 44038 7002 44090
rect 7014 44038 7066 44090
rect 7078 44038 7130 44090
rect 7142 44038 7194 44090
rect 7206 44038 7258 44090
rect 11950 44038 12002 44090
rect 12014 44038 12066 44090
rect 12078 44038 12130 44090
rect 12142 44038 12194 44090
rect 12206 44038 12258 44090
rect 16950 44038 17002 44090
rect 17014 44038 17066 44090
rect 17078 44038 17130 44090
rect 17142 44038 17194 44090
rect 17206 44038 17258 44090
rect 21950 44038 22002 44090
rect 22014 44038 22066 44090
rect 22078 44038 22130 44090
rect 22142 44038 22194 44090
rect 22206 44038 22258 44090
rect 26950 44038 27002 44090
rect 27014 44038 27066 44090
rect 27078 44038 27130 44090
rect 27142 44038 27194 44090
rect 27206 44038 27258 44090
rect 31950 44038 32002 44090
rect 32014 44038 32066 44090
rect 32078 44038 32130 44090
rect 32142 44038 32194 44090
rect 32206 44038 32258 44090
rect 36950 44038 37002 44090
rect 37014 44038 37066 44090
rect 37078 44038 37130 44090
rect 37142 44038 37194 44090
rect 37206 44038 37258 44090
rect 41950 44038 42002 44090
rect 42014 44038 42066 44090
rect 42078 44038 42130 44090
rect 42142 44038 42194 44090
rect 42206 44038 42258 44090
rect 46950 44038 47002 44090
rect 47014 44038 47066 44090
rect 47078 44038 47130 44090
rect 47142 44038 47194 44090
rect 47206 44038 47258 44090
rect 51950 44038 52002 44090
rect 52014 44038 52066 44090
rect 52078 44038 52130 44090
rect 52142 44038 52194 44090
rect 52206 44038 52258 44090
rect 56950 44038 57002 44090
rect 57014 44038 57066 44090
rect 57078 44038 57130 44090
rect 57142 44038 57194 44090
rect 57206 44038 57258 44090
rect 58532 43775 58584 43784
rect 58532 43741 58541 43775
rect 58541 43741 58575 43775
rect 58575 43741 58584 43775
rect 58532 43732 58584 43741
rect 2610 43494 2662 43546
rect 2674 43494 2726 43546
rect 2738 43494 2790 43546
rect 2802 43494 2854 43546
rect 2866 43494 2918 43546
rect 7610 43494 7662 43546
rect 7674 43494 7726 43546
rect 7738 43494 7790 43546
rect 7802 43494 7854 43546
rect 7866 43494 7918 43546
rect 12610 43494 12662 43546
rect 12674 43494 12726 43546
rect 12738 43494 12790 43546
rect 12802 43494 12854 43546
rect 12866 43494 12918 43546
rect 17610 43494 17662 43546
rect 17674 43494 17726 43546
rect 17738 43494 17790 43546
rect 17802 43494 17854 43546
rect 17866 43494 17918 43546
rect 22610 43494 22662 43546
rect 22674 43494 22726 43546
rect 22738 43494 22790 43546
rect 22802 43494 22854 43546
rect 22866 43494 22918 43546
rect 27610 43494 27662 43546
rect 27674 43494 27726 43546
rect 27738 43494 27790 43546
rect 27802 43494 27854 43546
rect 27866 43494 27918 43546
rect 32610 43494 32662 43546
rect 32674 43494 32726 43546
rect 32738 43494 32790 43546
rect 32802 43494 32854 43546
rect 32866 43494 32918 43546
rect 37610 43494 37662 43546
rect 37674 43494 37726 43546
rect 37738 43494 37790 43546
rect 37802 43494 37854 43546
rect 37866 43494 37918 43546
rect 42610 43494 42662 43546
rect 42674 43494 42726 43546
rect 42738 43494 42790 43546
rect 42802 43494 42854 43546
rect 42866 43494 42918 43546
rect 47610 43494 47662 43546
rect 47674 43494 47726 43546
rect 47738 43494 47790 43546
rect 47802 43494 47854 43546
rect 47866 43494 47918 43546
rect 52610 43494 52662 43546
rect 52674 43494 52726 43546
rect 52738 43494 52790 43546
rect 52802 43494 52854 43546
rect 52866 43494 52918 43546
rect 57610 43494 57662 43546
rect 57674 43494 57726 43546
rect 57738 43494 57790 43546
rect 57802 43494 57854 43546
rect 57866 43494 57918 43546
rect 1950 42950 2002 43002
rect 2014 42950 2066 43002
rect 2078 42950 2130 43002
rect 2142 42950 2194 43002
rect 2206 42950 2258 43002
rect 6950 42950 7002 43002
rect 7014 42950 7066 43002
rect 7078 42950 7130 43002
rect 7142 42950 7194 43002
rect 7206 42950 7258 43002
rect 11950 42950 12002 43002
rect 12014 42950 12066 43002
rect 12078 42950 12130 43002
rect 12142 42950 12194 43002
rect 12206 42950 12258 43002
rect 16950 42950 17002 43002
rect 17014 42950 17066 43002
rect 17078 42950 17130 43002
rect 17142 42950 17194 43002
rect 17206 42950 17258 43002
rect 21950 42950 22002 43002
rect 22014 42950 22066 43002
rect 22078 42950 22130 43002
rect 22142 42950 22194 43002
rect 22206 42950 22258 43002
rect 26950 42950 27002 43002
rect 27014 42950 27066 43002
rect 27078 42950 27130 43002
rect 27142 42950 27194 43002
rect 27206 42950 27258 43002
rect 31950 42950 32002 43002
rect 32014 42950 32066 43002
rect 32078 42950 32130 43002
rect 32142 42950 32194 43002
rect 32206 42950 32258 43002
rect 36950 42950 37002 43002
rect 37014 42950 37066 43002
rect 37078 42950 37130 43002
rect 37142 42950 37194 43002
rect 37206 42950 37258 43002
rect 41950 42950 42002 43002
rect 42014 42950 42066 43002
rect 42078 42950 42130 43002
rect 42142 42950 42194 43002
rect 42206 42950 42258 43002
rect 46950 42950 47002 43002
rect 47014 42950 47066 43002
rect 47078 42950 47130 43002
rect 47142 42950 47194 43002
rect 47206 42950 47258 43002
rect 51950 42950 52002 43002
rect 52014 42950 52066 43002
rect 52078 42950 52130 43002
rect 52142 42950 52194 43002
rect 52206 42950 52258 43002
rect 56950 42950 57002 43002
rect 57014 42950 57066 43002
rect 57078 42950 57130 43002
rect 57142 42950 57194 43002
rect 57206 42950 57258 43002
rect 58532 42687 58584 42696
rect 58532 42653 58541 42687
rect 58541 42653 58575 42687
rect 58575 42653 58584 42687
rect 58532 42644 58584 42653
rect 2610 42406 2662 42458
rect 2674 42406 2726 42458
rect 2738 42406 2790 42458
rect 2802 42406 2854 42458
rect 2866 42406 2918 42458
rect 7610 42406 7662 42458
rect 7674 42406 7726 42458
rect 7738 42406 7790 42458
rect 7802 42406 7854 42458
rect 7866 42406 7918 42458
rect 12610 42406 12662 42458
rect 12674 42406 12726 42458
rect 12738 42406 12790 42458
rect 12802 42406 12854 42458
rect 12866 42406 12918 42458
rect 17610 42406 17662 42458
rect 17674 42406 17726 42458
rect 17738 42406 17790 42458
rect 17802 42406 17854 42458
rect 17866 42406 17918 42458
rect 22610 42406 22662 42458
rect 22674 42406 22726 42458
rect 22738 42406 22790 42458
rect 22802 42406 22854 42458
rect 22866 42406 22918 42458
rect 27610 42406 27662 42458
rect 27674 42406 27726 42458
rect 27738 42406 27790 42458
rect 27802 42406 27854 42458
rect 27866 42406 27918 42458
rect 32610 42406 32662 42458
rect 32674 42406 32726 42458
rect 32738 42406 32790 42458
rect 32802 42406 32854 42458
rect 32866 42406 32918 42458
rect 37610 42406 37662 42458
rect 37674 42406 37726 42458
rect 37738 42406 37790 42458
rect 37802 42406 37854 42458
rect 37866 42406 37918 42458
rect 42610 42406 42662 42458
rect 42674 42406 42726 42458
rect 42738 42406 42790 42458
rect 42802 42406 42854 42458
rect 42866 42406 42918 42458
rect 47610 42406 47662 42458
rect 47674 42406 47726 42458
rect 47738 42406 47790 42458
rect 47802 42406 47854 42458
rect 47866 42406 47918 42458
rect 52610 42406 52662 42458
rect 52674 42406 52726 42458
rect 52738 42406 52790 42458
rect 52802 42406 52854 42458
rect 52866 42406 52918 42458
rect 57610 42406 57662 42458
rect 57674 42406 57726 42458
rect 57738 42406 57790 42458
rect 57802 42406 57854 42458
rect 57866 42406 57918 42458
rect 58532 42007 58584 42016
rect 58532 41973 58541 42007
rect 58541 41973 58575 42007
rect 58575 41973 58584 42007
rect 58532 41964 58584 41973
rect 1950 41862 2002 41914
rect 2014 41862 2066 41914
rect 2078 41862 2130 41914
rect 2142 41862 2194 41914
rect 2206 41862 2258 41914
rect 6950 41862 7002 41914
rect 7014 41862 7066 41914
rect 7078 41862 7130 41914
rect 7142 41862 7194 41914
rect 7206 41862 7258 41914
rect 11950 41862 12002 41914
rect 12014 41862 12066 41914
rect 12078 41862 12130 41914
rect 12142 41862 12194 41914
rect 12206 41862 12258 41914
rect 16950 41862 17002 41914
rect 17014 41862 17066 41914
rect 17078 41862 17130 41914
rect 17142 41862 17194 41914
rect 17206 41862 17258 41914
rect 21950 41862 22002 41914
rect 22014 41862 22066 41914
rect 22078 41862 22130 41914
rect 22142 41862 22194 41914
rect 22206 41862 22258 41914
rect 26950 41862 27002 41914
rect 27014 41862 27066 41914
rect 27078 41862 27130 41914
rect 27142 41862 27194 41914
rect 27206 41862 27258 41914
rect 31950 41862 32002 41914
rect 32014 41862 32066 41914
rect 32078 41862 32130 41914
rect 32142 41862 32194 41914
rect 32206 41862 32258 41914
rect 36950 41862 37002 41914
rect 37014 41862 37066 41914
rect 37078 41862 37130 41914
rect 37142 41862 37194 41914
rect 37206 41862 37258 41914
rect 41950 41862 42002 41914
rect 42014 41862 42066 41914
rect 42078 41862 42130 41914
rect 42142 41862 42194 41914
rect 42206 41862 42258 41914
rect 46950 41862 47002 41914
rect 47014 41862 47066 41914
rect 47078 41862 47130 41914
rect 47142 41862 47194 41914
rect 47206 41862 47258 41914
rect 51950 41862 52002 41914
rect 52014 41862 52066 41914
rect 52078 41862 52130 41914
rect 52142 41862 52194 41914
rect 52206 41862 52258 41914
rect 56950 41862 57002 41914
rect 57014 41862 57066 41914
rect 57078 41862 57130 41914
rect 57142 41862 57194 41914
rect 57206 41862 57258 41914
rect 2610 41318 2662 41370
rect 2674 41318 2726 41370
rect 2738 41318 2790 41370
rect 2802 41318 2854 41370
rect 2866 41318 2918 41370
rect 7610 41318 7662 41370
rect 7674 41318 7726 41370
rect 7738 41318 7790 41370
rect 7802 41318 7854 41370
rect 7866 41318 7918 41370
rect 12610 41318 12662 41370
rect 12674 41318 12726 41370
rect 12738 41318 12790 41370
rect 12802 41318 12854 41370
rect 12866 41318 12918 41370
rect 17610 41318 17662 41370
rect 17674 41318 17726 41370
rect 17738 41318 17790 41370
rect 17802 41318 17854 41370
rect 17866 41318 17918 41370
rect 22610 41318 22662 41370
rect 22674 41318 22726 41370
rect 22738 41318 22790 41370
rect 22802 41318 22854 41370
rect 22866 41318 22918 41370
rect 27610 41318 27662 41370
rect 27674 41318 27726 41370
rect 27738 41318 27790 41370
rect 27802 41318 27854 41370
rect 27866 41318 27918 41370
rect 32610 41318 32662 41370
rect 32674 41318 32726 41370
rect 32738 41318 32790 41370
rect 32802 41318 32854 41370
rect 32866 41318 32918 41370
rect 37610 41318 37662 41370
rect 37674 41318 37726 41370
rect 37738 41318 37790 41370
rect 37802 41318 37854 41370
rect 37866 41318 37918 41370
rect 42610 41318 42662 41370
rect 42674 41318 42726 41370
rect 42738 41318 42790 41370
rect 42802 41318 42854 41370
rect 42866 41318 42918 41370
rect 47610 41318 47662 41370
rect 47674 41318 47726 41370
rect 47738 41318 47790 41370
rect 47802 41318 47854 41370
rect 47866 41318 47918 41370
rect 52610 41318 52662 41370
rect 52674 41318 52726 41370
rect 52738 41318 52790 41370
rect 52802 41318 52854 41370
rect 52866 41318 52918 41370
rect 57610 41318 57662 41370
rect 57674 41318 57726 41370
rect 57738 41318 57790 41370
rect 57802 41318 57854 41370
rect 57866 41318 57918 41370
rect 58532 40919 58584 40928
rect 58532 40885 58541 40919
rect 58541 40885 58575 40919
rect 58575 40885 58584 40919
rect 58532 40876 58584 40885
rect 1950 40774 2002 40826
rect 2014 40774 2066 40826
rect 2078 40774 2130 40826
rect 2142 40774 2194 40826
rect 2206 40774 2258 40826
rect 6950 40774 7002 40826
rect 7014 40774 7066 40826
rect 7078 40774 7130 40826
rect 7142 40774 7194 40826
rect 7206 40774 7258 40826
rect 11950 40774 12002 40826
rect 12014 40774 12066 40826
rect 12078 40774 12130 40826
rect 12142 40774 12194 40826
rect 12206 40774 12258 40826
rect 16950 40774 17002 40826
rect 17014 40774 17066 40826
rect 17078 40774 17130 40826
rect 17142 40774 17194 40826
rect 17206 40774 17258 40826
rect 21950 40774 22002 40826
rect 22014 40774 22066 40826
rect 22078 40774 22130 40826
rect 22142 40774 22194 40826
rect 22206 40774 22258 40826
rect 26950 40774 27002 40826
rect 27014 40774 27066 40826
rect 27078 40774 27130 40826
rect 27142 40774 27194 40826
rect 27206 40774 27258 40826
rect 31950 40774 32002 40826
rect 32014 40774 32066 40826
rect 32078 40774 32130 40826
rect 32142 40774 32194 40826
rect 32206 40774 32258 40826
rect 36950 40774 37002 40826
rect 37014 40774 37066 40826
rect 37078 40774 37130 40826
rect 37142 40774 37194 40826
rect 37206 40774 37258 40826
rect 41950 40774 42002 40826
rect 42014 40774 42066 40826
rect 42078 40774 42130 40826
rect 42142 40774 42194 40826
rect 42206 40774 42258 40826
rect 46950 40774 47002 40826
rect 47014 40774 47066 40826
rect 47078 40774 47130 40826
rect 47142 40774 47194 40826
rect 47206 40774 47258 40826
rect 51950 40774 52002 40826
rect 52014 40774 52066 40826
rect 52078 40774 52130 40826
rect 52142 40774 52194 40826
rect 52206 40774 52258 40826
rect 56950 40774 57002 40826
rect 57014 40774 57066 40826
rect 57078 40774 57130 40826
rect 57142 40774 57194 40826
rect 57206 40774 57258 40826
rect 58532 40511 58584 40520
rect 58532 40477 58541 40511
rect 58541 40477 58575 40511
rect 58575 40477 58584 40511
rect 58532 40468 58584 40477
rect 2610 40230 2662 40282
rect 2674 40230 2726 40282
rect 2738 40230 2790 40282
rect 2802 40230 2854 40282
rect 2866 40230 2918 40282
rect 7610 40230 7662 40282
rect 7674 40230 7726 40282
rect 7738 40230 7790 40282
rect 7802 40230 7854 40282
rect 7866 40230 7918 40282
rect 12610 40230 12662 40282
rect 12674 40230 12726 40282
rect 12738 40230 12790 40282
rect 12802 40230 12854 40282
rect 12866 40230 12918 40282
rect 17610 40230 17662 40282
rect 17674 40230 17726 40282
rect 17738 40230 17790 40282
rect 17802 40230 17854 40282
rect 17866 40230 17918 40282
rect 22610 40230 22662 40282
rect 22674 40230 22726 40282
rect 22738 40230 22790 40282
rect 22802 40230 22854 40282
rect 22866 40230 22918 40282
rect 27610 40230 27662 40282
rect 27674 40230 27726 40282
rect 27738 40230 27790 40282
rect 27802 40230 27854 40282
rect 27866 40230 27918 40282
rect 32610 40230 32662 40282
rect 32674 40230 32726 40282
rect 32738 40230 32790 40282
rect 32802 40230 32854 40282
rect 32866 40230 32918 40282
rect 37610 40230 37662 40282
rect 37674 40230 37726 40282
rect 37738 40230 37790 40282
rect 37802 40230 37854 40282
rect 37866 40230 37918 40282
rect 42610 40230 42662 40282
rect 42674 40230 42726 40282
rect 42738 40230 42790 40282
rect 42802 40230 42854 40282
rect 42866 40230 42918 40282
rect 47610 40230 47662 40282
rect 47674 40230 47726 40282
rect 47738 40230 47790 40282
rect 47802 40230 47854 40282
rect 47866 40230 47918 40282
rect 52610 40230 52662 40282
rect 52674 40230 52726 40282
rect 52738 40230 52790 40282
rect 52802 40230 52854 40282
rect 52866 40230 52918 40282
rect 57610 40230 57662 40282
rect 57674 40230 57726 40282
rect 57738 40230 57790 40282
rect 57802 40230 57854 40282
rect 57866 40230 57918 40282
rect 1950 39686 2002 39738
rect 2014 39686 2066 39738
rect 2078 39686 2130 39738
rect 2142 39686 2194 39738
rect 2206 39686 2258 39738
rect 6950 39686 7002 39738
rect 7014 39686 7066 39738
rect 7078 39686 7130 39738
rect 7142 39686 7194 39738
rect 7206 39686 7258 39738
rect 11950 39686 12002 39738
rect 12014 39686 12066 39738
rect 12078 39686 12130 39738
rect 12142 39686 12194 39738
rect 12206 39686 12258 39738
rect 16950 39686 17002 39738
rect 17014 39686 17066 39738
rect 17078 39686 17130 39738
rect 17142 39686 17194 39738
rect 17206 39686 17258 39738
rect 21950 39686 22002 39738
rect 22014 39686 22066 39738
rect 22078 39686 22130 39738
rect 22142 39686 22194 39738
rect 22206 39686 22258 39738
rect 26950 39686 27002 39738
rect 27014 39686 27066 39738
rect 27078 39686 27130 39738
rect 27142 39686 27194 39738
rect 27206 39686 27258 39738
rect 31950 39686 32002 39738
rect 32014 39686 32066 39738
rect 32078 39686 32130 39738
rect 32142 39686 32194 39738
rect 32206 39686 32258 39738
rect 36950 39686 37002 39738
rect 37014 39686 37066 39738
rect 37078 39686 37130 39738
rect 37142 39686 37194 39738
rect 37206 39686 37258 39738
rect 41950 39686 42002 39738
rect 42014 39686 42066 39738
rect 42078 39686 42130 39738
rect 42142 39686 42194 39738
rect 42206 39686 42258 39738
rect 46950 39686 47002 39738
rect 47014 39686 47066 39738
rect 47078 39686 47130 39738
rect 47142 39686 47194 39738
rect 47206 39686 47258 39738
rect 51950 39686 52002 39738
rect 52014 39686 52066 39738
rect 52078 39686 52130 39738
rect 52142 39686 52194 39738
rect 52206 39686 52258 39738
rect 56950 39686 57002 39738
rect 57014 39686 57066 39738
rect 57078 39686 57130 39738
rect 57142 39686 57194 39738
rect 57206 39686 57258 39738
rect 58532 39423 58584 39432
rect 58532 39389 58541 39423
rect 58541 39389 58575 39423
rect 58575 39389 58584 39423
rect 58532 39380 58584 39389
rect 2610 39142 2662 39194
rect 2674 39142 2726 39194
rect 2738 39142 2790 39194
rect 2802 39142 2854 39194
rect 2866 39142 2918 39194
rect 7610 39142 7662 39194
rect 7674 39142 7726 39194
rect 7738 39142 7790 39194
rect 7802 39142 7854 39194
rect 7866 39142 7918 39194
rect 12610 39142 12662 39194
rect 12674 39142 12726 39194
rect 12738 39142 12790 39194
rect 12802 39142 12854 39194
rect 12866 39142 12918 39194
rect 17610 39142 17662 39194
rect 17674 39142 17726 39194
rect 17738 39142 17790 39194
rect 17802 39142 17854 39194
rect 17866 39142 17918 39194
rect 22610 39142 22662 39194
rect 22674 39142 22726 39194
rect 22738 39142 22790 39194
rect 22802 39142 22854 39194
rect 22866 39142 22918 39194
rect 27610 39142 27662 39194
rect 27674 39142 27726 39194
rect 27738 39142 27790 39194
rect 27802 39142 27854 39194
rect 27866 39142 27918 39194
rect 32610 39142 32662 39194
rect 32674 39142 32726 39194
rect 32738 39142 32790 39194
rect 32802 39142 32854 39194
rect 32866 39142 32918 39194
rect 37610 39142 37662 39194
rect 37674 39142 37726 39194
rect 37738 39142 37790 39194
rect 37802 39142 37854 39194
rect 37866 39142 37918 39194
rect 42610 39142 42662 39194
rect 42674 39142 42726 39194
rect 42738 39142 42790 39194
rect 42802 39142 42854 39194
rect 42866 39142 42918 39194
rect 47610 39142 47662 39194
rect 47674 39142 47726 39194
rect 47738 39142 47790 39194
rect 47802 39142 47854 39194
rect 47866 39142 47918 39194
rect 52610 39142 52662 39194
rect 52674 39142 52726 39194
rect 52738 39142 52790 39194
rect 52802 39142 52854 39194
rect 52866 39142 52918 39194
rect 57610 39142 57662 39194
rect 57674 39142 57726 39194
rect 57738 39142 57790 39194
rect 57802 39142 57854 39194
rect 57866 39142 57918 39194
rect 58532 38743 58584 38752
rect 58532 38709 58541 38743
rect 58541 38709 58575 38743
rect 58575 38709 58584 38743
rect 58532 38700 58584 38709
rect 1950 38598 2002 38650
rect 2014 38598 2066 38650
rect 2078 38598 2130 38650
rect 2142 38598 2194 38650
rect 2206 38598 2258 38650
rect 6950 38598 7002 38650
rect 7014 38598 7066 38650
rect 7078 38598 7130 38650
rect 7142 38598 7194 38650
rect 7206 38598 7258 38650
rect 11950 38598 12002 38650
rect 12014 38598 12066 38650
rect 12078 38598 12130 38650
rect 12142 38598 12194 38650
rect 12206 38598 12258 38650
rect 16950 38598 17002 38650
rect 17014 38598 17066 38650
rect 17078 38598 17130 38650
rect 17142 38598 17194 38650
rect 17206 38598 17258 38650
rect 21950 38598 22002 38650
rect 22014 38598 22066 38650
rect 22078 38598 22130 38650
rect 22142 38598 22194 38650
rect 22206 38598 22258 38650
rect 26950 38598 27002 38650
rect 27014 38598 27066 38650
rect 27078 38598 27130 38650
rect 27142 38598 27194 38650
rect 27206 38598 27258 38650
rect 31950 38598 32002 38650
rect 32014 38598 32066 38650
rect 32078 38598 32130 38650
rect 32142 38598 32194 38650
rect 32206 38598 32258 38650
rect 36950 38598 37002 38650
rect 37014 38598 37066 38650
rect 37078 38598 37130 38650
rect 37142 38598 37194 38650
rect 37206 38598 37258 38650
rect 41950 38598 42002 38650
rect 42014 38598 42066 38650
rect 42078 38598 42130 38650
rect 42142 38598 42194 38650
rect 42206 38598 42258 38650
rect 46950 38598 47002 38650
rect 47014 38598 47066 38650
rect 47078 38598 47130 38650
rect 47142 38598 47194 38650
rect 47206 38598 47258 38650
rect 51950 38598 52002 38650
rect 52014 38598 52066 38650
rect 52078 38598 52130 38650
rect 52142 38598 52194 38650
rect 52206 38598 52258 38650
rect 56950 38598 57002 38650
rect 57014 38598 57066 38650
rect 57078 38598 57130 38650
rect 57142 38598 57194 38650
rect 57206 38598 57258 38650
rect 2610 38054 2662 38106
rect 2674 38054 2726 38106
rect 2738 38054 2790 38106
rect 2802 38054 2854 38106
rect 2866 38054 2918 38106
rect 7610 38054 7662 38106
rect 7674 38054 7726 38106
rect 7738 38054 7790 38106
rect 7802 38054 7854 38106
rect 7866 38054 7918 38106
rect 12610 38054 12662 38106
rect 12674 38054 12726 38106
rect 12738 38054 12790 38106
rect 12802 38054 12854 38106
rect 12866 38054 12918 38106
rect 17610 38054 17662 38106
rect 17674 38054 17726 38106
rect 17738 38054 17790 38106
rect 17802 38054 17854 38106
rect 17866 38054 17918 38106
rect 22610 38054 22662 38106
rect 22674 38054 22726 38106
rect 22738 38054 22790 38106
rect 22802 38054 22854 38106
rect 22866 38054 22918 38106
rect 27610 38054 27662 38106
rect 27674 38054 27726 38106
rect 27738 38054 27790 38106
rect 27802 38054 27854 38106
rect 27866 38054 27918 38106
rect 32610 38054 32662 38106
rect 32674 38054 32726 38106
rect 32738 38054 32790 38106
rect 32802 38054 32854 38106
rect 32866 38054 32918 38106
rect 37610 38054 37662 38106
rect 37674 38054 37726 38106
rect 37738 38054 37790 38106
rect 37802 38054 37854 38106
rect 37866 38054 37918 38106
rect 42610 38054 42662 38106
rect 42674 38054 42726 38106
rect 42738 38054 42790 38106
rect 42802 38054 42854 38106
rect 42866 38054 42918 38106
rect 47610 38054 47662 38106
rect 47674 38054 47726 38106
rect 47738 38054 47790 38106
rect 47802 38054 47854 38106
rect 47866 38054 47918 38106
rect 52610 38054 52662 38106
rect 52674 38054 52726 38106
rect 52738 38054 52790 38106
rect 52802 38054 52854 38106
rect 52866 38054 52918 38106
rect 57610 38054 57662 38106
rect 57674 38054 57726 38106
rect 57738 38054 57790 38106
rect 57802 38054 57854 38106
rect 57866 38054 57918 38106
rect 58532 37655 58584 37664
rect 58532 37621 58541 37655
rect 58541 37621 58575 37655
rect 58575 37621 58584 37655
rect 58532 37612 58584 37621
rect 1950 37510 2002 37562
rect 2014 37510 2066 37562
rect 2078 37510 2130 37562
rect 2142 37510 2194 37562
rect 2206 37510 2258 37562
rect 6950 37510 7002 37562
rect 7014 37510 7066 37562
rect 7078 37510 7130 37562
rect 7142 37510 7194 37562
rect 7206 37510 7258 37562
rect 11950 37510 12002 37562
rect 12014 37510 12066 37562
rect 12078 37510 12130 37562
rect 12142 37510 12194 37562
rect 12206 37510 12258 37562
rect 16950 37510 17002 37562
rect 17014 37510 17066 37562
rect 17078 37510 17130 37562
rect 17142 37510 17194 37562
rect 17206 37510 17258 37562
rect 21950 37510 22002 37562
rect 22014 37510 22066 37562
rect 22078 37510 22130 37562
rect 22142 37510 22194 37562
rect 22206 37510 22258 37562
rect 26950 37510 27002 37562
rect 27014 37510 27066 37562
rect 27078 37510 27130 37562
rect 27142 37510 27194 37562
rect 27206 37510 27258 37562
rect 31950 37510 32002 37562
rect 32014 37510 32066 37562
rect 32078 37510 32130 37562
rect 32142 37510 32194 37562
rect 32206 37510 32258 37562
rect 36950 37510 37002 37562
rect 37014 37510 37066 37562
rect 37078 37510 37130 37562
rect 37142 37510 37194 37562
rect 37206 37510 37258 37562
rect 41950 37510 42002 37562
rect 42014 37510 42066 37562
rect 42078 37510 42130 37562
rect 42142 37510 42194 37562
rect 42206 37510 42258 37562
rect 46950 37510 47002 37562
rect 47014 37510 47066 37562
rect 47078 37510 47130 37562
rect 47142 37510 47194 37562
rect 47206 37510 47258 37562
rect 51950 37510 52002 37562
rect 52014 37510 52066 37562
rect 52078 37510 52130 37562
rect 52142 37510 52194 37562
rect 52206 37510 52258 37562
rect 56950 37510 57002 37562
rect 57014 37510 57066 37562
rect 57078 37510 57130 37562
rect 57142 37510 57194 37562
rect 57206 37510 57258 37562
rect 58532 37315 58584 37324
rect 58532 37281 58541 37315
rect 58541 37281 58575 37315
rect 58575 37281 58584 37315
rect 58532 37272 58584 37281
rect 2610 36966 2662 37018
rect 2674 36966 2726 37018
rect 2738 36966 2790 37018
rect 2802 36966 2854 37018
rect 2866 36966 2918 37018
rect 7610 36966 7662 37018
rect 7674 36966 7726 37018
rect 7738 36966 7790 37018
rect 7802 36966 7854 37018
rect 7866 36966 7918 37018
rect 12610 36966 12662 37018
rect 12674 36966 12726 37018
rect 12738 36966 12790 37018
rect 12802 36966 12854 37018
rect 12866 36966 12918 37018
rect 17610 36966 17662 37018
rect 17674 36966 17726 37018
rect 17738 36966 17790 37018
rect 17802 36966 17854 37018
rect 17866 36966 17918 37018
rect 22610 36966 22662 37018
rect 22674 36966 22726 37018
rect 22738 36966 22790 37018
rect 22802 36966 22854 37018
rect 22866 36966 22918 37018
rect 27610 36966 27662 37018
rect 27674 36966 27726 37018
rect 27738 36966 27790 37018
rect 27802 36966 27854 37018
rect 27866 36966 27918 37018
rect 32610 36966 32662 37018
rect 32674 36966 32726 37018
rect 32738 36966 32790 37018
rect 32802 36966 32854 37018
rect 32866 36966 32918 37018
rect 37610 36966 37662 37018
rect 37674 36966 37726 37018
rect 37738 36966 37790 37018
rect 37802 36966 37854 37018
rect 37866 36966 37918 37018
rect 42610 36966 42662 37018
rect 42674 36966 42726 37018
rect 42738 36966 42790 37018
rect 42802 36966 42854 37018
rect 42866 36966 42918 37018
rect 47610 36966 47662 37018
rect 47674 36966 47726 37018
rect 47738 36966 47790 37018
rect 47802 36966 47854 37018
rect 47866 36966 47918 37018
rect 52610 36966 52662 37018
rect 52674 36966 52726 37018
rect 52738 36966 52790 37018
rect 52802 36966 52854 37018
rect 52866 36966 52918 37018
rect 57610 36966 57662 37018
rect 57674 36966 57726 37018
rect 57738 36966 57790 37018
rect 57802 36966 57854 37018
rect 57866 36966 57918 37018
rect 1950 36422 2002 36474
rect 2014 36422 2066 36474
rect 2078 36422 2130 36474
rect 2142 36422 2194 36474
rect 2206 36422 2258 36474
rect 6950 36422 7002 36474
rect 7014 36422 7066 36474
rect 7078 36422 7130 36474
rect 7142 36422 7194 36474
rect 7206 36422 7258 36474
rect 11950 36422 12002 36474
rect 12014 36422 12066 36474
rect 12078 36422 12130 36474
rect 12142 36422 12194 36474
rect 12206 36422 12258 36474
rect 16950 36422 17002 36474
rect 17014 36422 17066 36474
rect 17078 36422 17130 36474
rect 17142 36422 17194 36474
rect 17206 36422 17258 36474
rect 21950 36422 22002 36474
rect 22014 36422 22066 36474
rect 22078 36422 22130 36474
rect 22142 36422 22194 36474
rect 22206 36422 22258 36474
rect 26950 36422 27002 36474
rect 27014 36422 27066 36474
rect 27078 36422 27130 36474
rect 27142 36422 27194 36474
rect 27206 36422 27258 36474
rect 31950 36422 32002 36474
rect 32014 36422 32066 36474
rect 32078 36422 32130 36474
rect 32142 36422 32194 36474
rect 32206 36422 32258 36474
rect 36950 36422 37002 36474
rect 37014 36422 37066 36474
rect 37078 36422 37130 36474
rect 37142 36422 37194 36474
rect 37206 36422 37258 36474
rect 41950 36422 42002 36474
rect 42014 36422 42066 36474
rect 42078 36422 42130 36474
rect 42142 36422 42194 36474
rect 42206 36422 42258 36474
rect 46950 36422 47002 36474
rect 47014 36422 47066 36474
rect 47078 36422 47130 36474
rect 47142 36422 47194 36474
rect 47206 36422 47258 36474
rect 51950 36422 52002 36474
rect 52014 36422 52066 36474
rect 52078 36422 52130 36474
rect 52142 36422 52194 36474
rect 52206 36422 52258 36474
rect 56950 36422 57002 36474
rect 57014 36422 57066 36474
rect 57078 36422 57130 36474
rect 57142 36422 57194 36474
rect 57206 36422 57258 36474
rect 58532 36159 58584 36168
rect 58532 36125 58541 36159
rect 58541 36125 58575 36159
rect 58575 36125 58584 36159
rect 58532 36116 58584 36125
rect 2610 35878 2662 35930
rect 2674 35878 2726 35930
rect 2738 35878 2790 35930
rect 2802 35878 2854 35930
rect 2866 35878 2918 35930
rect 7610 35878 7662 35930
rect 7674 35878 7726 35930
rect 7738 35878 7790 35930
rect 7802 35878 7854 35930
rect 7866 35878 7918 35930
rect 12610 35878 12662 35930
rect 12674 35878 12726 35930
rect 12738 35878 12790 35930
rect 12802 35878 12854 35930
rect 12866 35878 12918 35930
rect 17610 35878 17662 35930
rect 17674 35878 17726 35930
rect 17738 35878 17790 35930
rect 17802 35878 17854 35930
rect 17866 35878 17918 35930
rect 22610 35878 22662 35930
rect 22674 35878 22726 35930
rect 22738 35878 22790 35930
rect 22802 35878 22854 35930
rect 22866 35878 22918 35930
rect 27610 35878 27662 35930
rect 27674 35878 27726 35930
rect 27738 35878 27790 35930
rect 27802 35878 27854 35930
rect 27866 35878 27918 35930
rect 32610 35878 32662 35930
rect 32674 35878 32726 35930
rect 32738 35878 32790 35930
rect 32802 35878 32854 35930
rect 32866 35878 32918 35930
rect 37610 35878 37662 35930
rect 37674 35878 37726 35930
rect 37738 35878 37790 35930
rect 37802 35878 37854 35930
rect 37866 35878 37918 35930
rect 42610 35878 42662 35930
rect 42674 35878 42726 35930
rect 42738 35878 42790 35930
rect 42802 35878 42854 35930
rect 42866 35878 42918 35930
rect 47610 35878 47662 35930
rect 47674 35878 47726 35930
rect 47738 35878 47790 35930
rect 47802 35878 47854 35930
rect 47866 35878 47918 35930
rect 52610 35878 52662 35930
rect 52674 35878 52726 35930
rect 52738 35878 52790 35930
rect 52802 35878 52854 35930
rect 52866 35878 52918 35930
rect 57610 35878 57662 35930
rect 57674 35878 57726 35930
rect 57738 35878 57790 35930
rect 57802 35878 57854 35930
rect 57866 35878 57918 35930
rect 58532 35479 58584 35488
rect 58532 35445 58541 35479
rect 58541 35445 58575 35479
rect 58575 35445 58584 35479
rect 58532 35436 58584 35445
rect 1950 35334 2002 35386
rect 2014 35334 2066 35386
rect 2078 35334 2130 35386
rect 2142 35334 2194 35386
rect 2206 35334 2258 35386
rect 6950 35334 7002 35386
rect 7014 35334 7066 35386
rect 7078 35334 7130 35386
rect 7142 35334 7194 35386
rect 7206 35334 7258 35386
rect 11950 35334 12002 35386
rect 12014 35334 12066 35386
rect 12078 35334 12130 35386
rect 12142 35334 12194 35386
rect 12206 35334 12258 35386
rect 16950 35334 17002 35386
rect 17014 35334 17066 35386
rect 17078 35334 17130 35386
rect 17142 35334 17194 35386
rect 17206 35334 17258 35386
rect 21950 35334 22002 35386
rect 22014 35334 22066 35386
rect 22078 35334 22130 35386
rect 22142 35334 22194 35386
rect 22206 35334 22258 35386
rect 26950 35334 27002 35386
rect 27014 35334 27066 35386
rect 27078 35334 27130 35386
rect 27142 35334 27194 35386
rect 27206 35334 27258 35386
rect 31950 35334 32002 35386
rect 32014 35334 32066 35386
rect 32078 35334 32130 35386
rect 32142 35334 32194 35386
rect 32206 35334 32258 35386
rect 36950 35334 37002 35386
rect 37014 35334 37066 35386
rect 37078 35334 37130 35386
rect 37142 35334 37194 35386
rect 37206 35334 37258 35386
rect 41950 35334 42002 35386
rect 42014 35334 42066 35386
rect 42078 35334 42130 35386
rect 42142 35334 42194 35386
rect 42206 35334 42258 35386
rect 46950 35334 47002 35386
rect 47014 35334 47066 35386
rect 47078 35334 47130 35386
rect 47142 35334 47194 35386
rect 47206 35334 47258 35386
rect 51950 35334 52002 35386
rect 52014 35334 52066 35386
rect 52078 35334 52130 35386
rect 52142 35334 52194 35386
rect 52206 35334 52258 35386
rect 56950 35334 57002 35386
rect 57014 35334 57066 35386
rect 57078 35334 57130 35386
rect 57142 35334 57194 35386
rect 57206 35334 57258 35386
rect 2610 34790 2662 34842
rect 2674 34790 2726 34842
rect 2738 34790 2790 34842
rect 2802 34790 2854 34842
rect 2866 34790 2918 34842
rect 7610 34790 7662 34842
rect 7674 34790 7726 34842
rect 7738 34790 7790 34842
rect 7802 34790 7854 34842
rect 7866 34790 7918 34842
rect 12610 34790 12662 34842
rect 12674 34790 12726 34842
rect 12738 34790 12790 34842
rect 12802 34790 12854 34842
rect 12866 34790 12918 34842
rect 17610 34790 17662 34842
rect 17674 34790 17726 34842
rect 17738 34790 17790 34842
rect 17802 34790 17854 34842
rect 17866 34790 17918 34842
rect 22610 34790 22662 34842
rect 22674 34790 22726 34842
rect 22738 34790 22790 34842
rect 22802 34790 22854 34842
rect 22866 34790 22918 34842
rect 27610 34790 27662 34842
rect 27674 34790 27726 34842
rect 27738 34790 27790 34842
rect 27802 34790 27854 34842
rect 27866 34790 27918 34842
rect 32610 34790 32662 34842
rect 32674 34790 32726 34842
rect 32738 34790 32790 34842
rect 32802 34790 32854 34842
rect 32866 34790 32918 34842
rect 37610 34790 37662 34842
rect 37674 34790 37726 34842
rect 37738 34790 37790 34842
rect 37802 34790 37854 34842
rect 37866 34790 37918 34842
rect 42610 34790 42662 34842
rect 42674 34790 42726 34842
rect 42738 34790 42790 34842
rect 42802 34790 42854 34842
rect 42866 34790 42918 34842
rect 47610 34790 47662 34842
rect 47674 34790 47726 34842
rect 47738 34790 47790 34842
rect 47802 34790 47854 34842
rect 47866 34790 47918 34842
rect 52610 34790 52662 34842
rect 52674 34790 52726 34842
rect 52738 34790 52790 34842
rect 52802 34790 52854 34842
rect 52866 34790 52918 34842
rect 57610 34790 57662 34842
rect 57674 34790 57726 34842
rect 57738 34790 57790 34842
rect 57802 34790 57854 34842
rect 57866 34790 57918 34842
rect 58532 34391 58584 34400
rect 58532 34357 58541 34391
rect 58541 34357 58575 34391
rect 58575 34357 58584 34391
rect 58532 34348 58584 34357
rect 1950 34246 2002 34298
rect 2014 34246 2066 34298
rect 2078 34246 2130 34298
rect 2142 34246 2194 34298
rect 2206 34246 2258 34298
rect 6950 34246 7002 34298
rect 7014 34246 7066 34298
rect 7078 34246 7130 34298
rect 7142 34246 7194 34298
rect 7206 34246 7258 34298
rect 11950 34246 12002 34298
rect 12014 34246 12066 34298
rect 12078 34246 12130 34298
rect 12142 34246 12194 34298
rect 12206 34246 12258 34298
rect 16950 34246 17002 34298
rect 17014 34246 17066 34298
rect 17078 34246 17130 34298
rect 17142 34246 17194 34298
rect 17206 34246 17258 34298
rect 21950 34246 22002 34298
rect 22014 34246 22066 34298
rect 22078 34246 22130 34298
rect 22142 34246 22194 34298
rect 22206 34246 22258 34298
rect 26950 34246 27002 34298
rect 27014 34246 27066 34298
rect 27078 34246 27130 34298
rect 27142 34246 27194 34298
rect 27206 34246 27258 34298
rect 31950 34246 32002 34298
rect 32014 34246 32066 34298
rect 32078 34246 32130 34298
rect 32142 34246 32194 34298
rect 32206 34246 32258 34298
rect 36950 34246 37002 34298
rect 37014 34246 37066 34298
rect 37078 34246 37130 34298
rect 37142 34246 37194 34298
rect 37206 34246 37258 34298
rect 41950 34246 42002 34298
rect 42014 34246 42066 34298
rect 42078 34246 42130 34298
rect 42142 34246 42194 34298
rect 42206 34246 42258 34298
rect 46950 34246 47002 34298
rect 47014 34246 47066 34298
rect 47078 34246 47130 34298
rect 47142 34246 47194 34298
rect 47206 34246 47258 34298
rect 51950 34246 52002 34298
rect 52014 34246 52066 34298
rect 52078 34246 52130 34298
rect 52142 34246 52194 34298
rect 52206 34246 52258 34298
rect 56950 34246 57002 34298
rect 57014 34246 57066 34298
rect 57078 34246 57130 34298
rect 57142 34246 57194 34298
rect 57206 34246 57258 34298
rect 58532 33983 58584 33992
rect 58532 33949 58541 33983
rect 58541 33949 58575 33983
rect 58575 33949 58584 33983
rect 58532 33940 58584 33949
rect 2610 33702 2662 33754
rect 2674 33702 2726 33754
rect 2738 33702 2790 33754
rect 2802 33702 2854 33754
rect 2866 33702 2918 33754
rect 7610 33702 7662 33754
rect 7674 33702 7726 33754
rect 7738 33702 7790 33754
rect 7802 33702 7854 33754
rect 7866 33702 7918 33754
rect 12610 33702 12662 33754
rect 12674 33702 12726 33754
rect 12738 33702 12790 33754
rect 12802 33702 12854 33754
rect 12866 33702 12918 33754
rect 17610 33702 17662 33754
rect 17674 33702 17726 33754
rect 17738 33702 17790 33754
rect 17802 33702 17854 33754
rect 17866 33702 17918 33754
rect 22610 33702 22662 33754
rect 22674 33702 22726 33754
rect 22738 33702 22790 33754
rect 22802 33702 22854 33754
rect 22866 33702 22918 33754
rect 27610 33702 27662 33754
rect 27674 33702 27726 33754
rect 27738 33702 27790 33754
rect 27802 33702 27854 33754
rect 27866 33702 27918 33754
rect 32610 33702 32662 33754
rect 32674 33702 32726 33754
rect 32738 33702 32790 33754
rect 32802 33702 32854 33754
rect 32866 33702 32918 33754
rect 37610 33702 37662 33754
rect 37674 33702 37726 33754
rect 37738 33702 37790 33754
rect 37802 33702 37854 33754
rect 37866 33702 37918 33754
rect 42610 33702 42662 33754
rect 42674 33702 42726 33754
rect 42738 33702 42790 33754
rect 42802 33702 42854 33754
rect 42866 33702 42918 33754
rect 47610 33702 47662 33754
rect 47674 33702 47726 33754
rect 47738 33702 47790 33754
rect 47802 33702 47854 33754
rect 47866 33702 47918 33754
rect 52610 33702 52662 33754
rect 52674 33702 52726 33754
rect 52738 33702 52790 33754
rect 52802 33702 52854 33754
rect 52866 33702 52918 33754
rect 57610 33702 57662 33754
rect 57674 33702 57726 33754
rect 57738 33702 57790 33754
rect 57802 33702 57854 33754
rect 57866 33702 57918 33754
rect 1950 33158 2002 33210
rect 2014 33158 2066 33210
rect 2078 33158 2130 33210
rect 2142 33158 2194 33210
rect 2206 33158 2258 33210
rect 6950 33158 7002 33210
rect 7014 33158 7066 33210
rect 7078 33158 7130 33210
rect 7142 33158 7194 33210
rect 7206 33158 7258 33210
rect 11950 33158 12002 33210
rect 12014 33158 12066 33210
rect 12078 33158 12130 33210
rect 12142 33158 12194 33210
rect 12206 33158 12258 33210
rect 16950 33158 17002 33210
rect 17014 33158 17066 33210
rect 17078 33158 17130 33210
rect 17142 33158 17194 33210
rect 17206 33158 17258 33210
rect 21950 33158 22002 33210
rect 22014 33158 22066 33210
rect 22078 33158 22130 33210
rect 22142 33158 22194 33210
rect 22206 33158 22258 33210
rect 26950 33158 27002 33210
rect 27014 33158 27066 33210
rect 27078 33158 27130 33210
rect 27142 33158 27194 33210
rect 27206 33158 27258 33210
rect 31950 33158 32002 33210
rect 32014 33158 32066 33210
rect 32078 33158 32130 33210
rect 32142 33158 32194 33210
rect 32206 33158 32258 33210
rect 36950 33158 37002 33210
rect 37014 33158 37066 33210
rect 37078 33158 37130 33210
rect 37142 33158 37194 33210
rect 37206 33158 37258 33210
rect 41950 33158 42002 33210
rect 42014 33158 42066 33210
rect 42078 33158 42130 33210
rect 42142 33158 42194 33210
rect 42206 33158 42258 33210
rect 46950 33158 47002 33210
rect 47014 33158 47066 33210
rect 47078 33158 47130 33210
rect 47142 33158 47194 33210
rect 47206 33158 47258 33210
rect 51950 33158 52002 33210
rect 52014 33158 52066 33210
rect 52078 33158 52130 33210
rect 52142 33158 52194 33210
rect 52206 33158 52258 33210
rect 56950 33158 57002 33210
rect 57014 33158 57066 33210
rect 57078 33158 57130 33210
rect 57142 33158 57194 33210
rect 57206 33158 57258 33210
rect 58532 32895 58584 32904
rect 58532 32861 58541 32895
rect 58541 32861 58575 32895
rect 58575 32861 58584 32895
rect 58532 32852 58584 32861
rect 2610 32614 2662 32666
rect 2674 32614 2726 32666
rect 2738 32614 2790 32666
rect 2802 32614 2854 32666
rect 2866 32614 2918 32666
rect 7610 32614 7662 32666
rect 7674 32614 7726 32666
rect 7738 32614 7790 32666
rect 7802 32614 7854 32666
rect 7866 32614 7918 32666
rect 12610 32614 12662 32666
rect 12674 32614 12726 32666
rect 12738 32614 12790 32666
rect 12802 32614 12854 32666
rect 12866 32614 12918 32666
rect 17610 32614 17662 32666
rect 17674 32614 17726 32666
rect 17738 32614 17790 32666
rect 17802 32614 17854 32666
rect 17866 32614 17918 32666
rect 22610 32614 22662 32666
rect 22674 32614 22726 32666
rect 22738 32614 22790 32666
rect 22802 32614 22854 32666
rect 22866 32614 22918 32666
rect 27610 32614 27662 32666
rect 27674 32614 27726 32666
rect 27738 32614 27790 32666
rect 27802 32614 27854 32666
rect 27866 32614 27918 32666
rect 32610 32614 32662 32666
rect 32674 32614 32726 32666
rect 32738 32614 32790 32666
rect 32802 32614 32854 32666
rect 32866 32614 32918 32666
rect 37610 32614 37662 32666
rect 37674 32614 37726 32666
rect 37738 32614 37790 32666
rect 37802 32614 37854 32666
rect 37866 32614 37918 32666
rect 42610 32614 42662 32666
rect 42674 32614 42726 32666
rect 42738 32614 42790 32666
rect 42802 32614 42854 32666
rect 42866 32614 42918 32666
rect 47610 32614 47662 32666
rect 47674 32614 47726 32666
rect 47738 32614 47790 32666
rect 47802 32614 47854 32666
rect 47866 32614 47918 32666
rect 52610 32614 52662 32666
rect 52674 32614 52726 32666
rect 52738 32614 52790 32666
rect 52802 32614 52854 32666
rect 52866 32614 52918 32666
rect 57610 32614 57662 32666
rect 57674 32614 57726 32666
rect 57738 32614 57790 32666
rect 57802 32614 57854 32666
rect 57866 32614 57918 32666
rect 58532 32215 58584 32224
rect 58532 32181 58541 32215
rect 58541 32181 58575 32215
rect 58575 32181 58584 32215
rect 58532 32172 58584 32181
rect 1950 32070 2002 32122
rect 2014 32070 2066 32122
rect 2078 32070 2130 32122
rect 2142 32070 2194 32122
rect 2206 32070 2258 32122
rect 6950 32070 7002 32122
rect 7014 32070 7066 32122
rect 7078 32070 7130 32122
rect 7142 32070 7194 32122
rect 7206 32070 7258 32122
rect 11950 32070 12002 32122
rect 12014 32070 12066 32122
rect 12078 32070 12130 32122
rect 12142 32070 12194 32122
rect 12206 32070 12258 32122
rect 16950 32070 17002 32122
rect 17014 32070 17066 32122
rect 17078 32070 17130 32122
rect 17142 32070 17194 32122
rect 17206 32070 17258 32122
rect 21950 32070 22002 32122
rect 22014 32070 22066 32122
rect 22078 32070 22130 32122
rect 22142 32070 22194 32122
rect 22206 32070 22258 32122
rect 26950 32070 27002 32122
rect 27014 32070 27066 32122
rect 27078 32070 27130 32122
rect 27142 32070 27194 32122
rect 27206 32070 27258 32122
rect 31950 32070 32002 32122
rect 32014 32070 32066 32122
rect 32078 32070 32130 32122
rect 32142 32070 32194 32122
rect 32206 32070 32258 32122
rect 36950 32070 37002 32122
rect 37014 32070 37066 32122
rect 37078 32070 37130 32122
rect 37142 32070 37194 32122
rect 37206 32070 37258 32122
rect 41950 32070 42002 32122
rect 42014 32070 42066 32122
rect 42078 32070 42130 32122
rect 42142 32070 42194 32122
rect 42206 32070 42258 32122
rect 46950 32070 47002 32122
rect 47014 32070 47066 32122
rect 47078 32070 47130 32122
rect 47142 32070 47194 32122
rect 47206 32070 47258 32122
rect 51950 32070 52002 32122
rect 52014 32070 52066 32122
rect 52078 32070 52130 32122
rect 52142 32070 52194 32122
rect 52206 32070 52258 32122
rect 56950 32070 57002 32122
rect 57014 32070 57066 32122
rect 57078 32070 57130 32122
rect 57142 32070 57194 32122
rect 57206 32070 57258 32122
rect 2610 31526 2662 31578
rect 2674 31526 2726 31578
rect 2738 31526 2790 31578
rect 2802 31526 2854 31578
rect 2866 31526 2918 31578
rect 7610 31526 7662 31578
rect 7674 31526 7726 31578
rect 7738 31526 7790 31578
rect 7802 31526 7854 31578
rect 7866 31526 7918 31578
rect 12610 31526 12662 31578
rect 12674 31526 12726 31578
rect 12738 31526 12790 31578
rect 12802 31526 12854 31578
rect 12866 31526 12918 31578
rect 17610 31526 17662 31578
rect 17674 31526 17726 31578
rect 17738 31526 17790 31578
rect 17802 31526 17854 31578
rect 17866 31526 17918 31578
rect 22610 31526 22662 31578
rect 22674 31526 22726 31578
rect 22738 31526 22790 31578
rect 22802 31526 22854 31578
rect 22866 31526 22918 31578
rect 27610 31526 27662 31578
rect 27674 31526 27726 31578
rect 27738 31526 27790 31578
rect 27802 31526 27854 31578
rect 27866 31526 27918 31578
rect 32610 31526 32662 31578
rect 32674 31526 32726 31578
rect 32738 31526 32790 31578
rect 32802 31526 32854 31578
rect 32866 31526 32918 31578
rect 37610 31526 37662 31578
rect 37674 31526 37726 31578
rect 37738 31526 37790 31578
rect 37802 31526 37854 31578
rect 37866 31526 37918 31578
rect 42610 31526 42662 31578
rect 42674 31526 42726 31578
rect 42738 31526 42790 31578
rect 42802 31526 42854 31578
rect 42866 31526 42918 31578
rect 47610 31526 47662 31578
rect 47674 31526 47726 31578
rect 47738 31526 47790 31578
rect 47802 31526 47854 31578
rect 47866 31526 47918 31578
rect 52610 31526 52662 31578
rect 52674 31526 52726 31578
rect 52738 31526 52790 31578
rect 52802 31526 52854 31578
rect 52866 31526 52918 31578
rect 57610 31526 57662 31578
rect 57674 31526 57726 31578
rect 57738 31526 57790 31578
rect 57802 31526 57854 31578
rect 57866 31526 57918 31578
rect 58532 31127 58584 31136
rect 58532 31093 58541 31127
rect 58541 31093 58575 31127
rect 58575 31093 58584 31127
rect 58532 31084 58584 31093
rect 1950 30982 2002 31034
rect 2014 30982 2066 31034
rect 2078 30982 2130 31034
rect 2142 30982 2194 31034
rect 2206 30982 2258 31034
rect 6950 30982 7002 31034
rect 7014 30982 7066 31034
rect 7078 30982 7130 31034
rect 7142 30982 7194 31034
rect 7206 30982 7258 31034
rect 11950 30982 12002 31034
rect 12014 30982 12066 31034
rect 12078 30982 12130 31034
rect 12142 30982 12194 31034
rect 12206 30982 12258 31034
rect 16950 30982 17002 31034
rect 17014 30982 17066 31034
rect 17078 30982 17130 31034
rect 17142 30982 17194 31034
rect 17206 30982 17258 31034
rect 21950 30982 22002 31034
rect 22014 30982 22066 31034
rect 22078 30982 22130 31034
rect 22142 30982 22194 31034
rect 22206 30982 22258 31034
rect 26950 30982 27002 31034
rect 27014 30982 27066 31034
rect 27078 30982 27130 31034
rect 27142 30982 27194 31034
rect 27206 30982 27258 31034
rect 31950 30982 32002 31034
rect 32014 30982 32066 31034
rect 32078 30982 32130 31034
rect 32142 30982 32194 31034
rect 32206 30982 32258 31034
rect 36950 30982 37002 31034
rect 37014 30982 37066 31034
rect 37078 30982 37130 31034
rect 37142 30982 37194 31034
rect 37206 30982 37258 31034
rect 41950 30982 42002 31034
rect 42014 30982 42066 31034
rect 42078 30982 42130 31034
rect 42142 30982 42194 31034
rect 42206 30982 42258 31034
rect 46950 30982 47002 31034
rect 47014 30982 47066 31034
rect 47078 30982 47130 31034
rect 47142 30982 47194 31034
rect 47206 30982 47258 31034
rect 51950 30982 52002 31034
rect 52014 30982 52066 31034
rect 52078 30982 52130 31034
rect 52142 30982 52194 31034
rect 52206 30982 52258 31034
rect 56950 30982 57002 31034
rect 57014 30982 57066 31034
rect 57078 30982 57130 31034
rect 57142 30982 57194 31034
rect 57206 30982 57258 31034
rect 58532 30719 58584 30728
rect 58532 30685 58541 30719
rect 58541 30685 58575 30719
rect 58575 30685 58584 30719
rect 58532 30676 58584 30685
rect 2610 30438 2662 30490
rect 2674 30438 2726 30490
rect 2738 30438 2790 30490
rect 2802 30438 2854 30490
rect 2866 30438 2918 30490
rect 7610 30438 7662 30490
rect 7674 30438 7726 30490
rect 7738 30438 7790 30490
rect 7802 30438 7854 30490
rect 7866 30438 7918 30490
rect 12610 30438 12662 30490
rect 12674 30438 12726 30490
rect 12738 30438 12790 30490
rect 12802 30438 12854 30490
rect 12866 30438 12918 30490
rect 17610 30438 17662 30490
rect 17674 30438 17726 30490
rect 17738 30438 17790 30490
rect 17802 30438 17854 30490
rect 17866 30438 17918 30490
rect 22610 30438 22662 30490
rect 22674 30438 22726 30490
rect 22738 30438 22790 30490
rect 22802 30438 22854 30490
rect 22866 30438 22918 30490
rect 27610 30438 27662 30490
rect 27674 30438 27726 30490
rect 27738 30438 27790 30490
rect 27802 30438 27854 30490
rect 27866 30438 27918 30490
rect 32610 30438 32662 30490
rect 32674 30438 32726 30490
rect 32738 30438 32790 30490
rect 32802 30438 32854 30490
rect 32866 30438 32918 30490
rect 37610 30438 37662 30490
rect 37674 30438 37726 30490
rect 37738 30438 37790 30490
rect 37802 30438 37854 30490
rect 37866 30438 37918 30490
rect 42610 30438 42662 30490
rect 42674 30438 42726 30490
rect 42738 30438 42790 30490
rect 42802 30438 42854 30490
rect 42866 30438 42918 30490
rect 47610 30438 47662 30490
rect 47674 30438 47726 30490
rect 47738 30438 47790 30490
rect 47802 30438 47854 30490
rect 47866 30438 47918 30490
rect 52610 30438 52662 30490
rect 52674 30438 52726 30490
rect 52738 30438 52790 30490
rect 52802 30438 52854 30490
rect 52866 30438 52918 30490
rect 57610 30438 57662 30490
rect 57674 30438 57726 30490
rect 57738 30438 57790 30490
rect 57802 30438 57854 30490
rect 57866 30438 57918 30490
rect 1950 29894 2002 29946
rect 2014 29894 2066 29946
rect 2078 29894 2130 29946
rect 2142 29894 2194 29946
rect 2206 29894 2258 29946
rect 6950 29894 7002 29946
rect 7014 29894 7066 29946
rect 7078 29894 7130 29946
rect 7142 29894 7194 29946
rect 7206 29894 7258 29946
rect 11950 29894 12002 29946
rect 12014 29894 12066 29946
rect 12078 29894 12130 29946
rect 12142 29894 12194 29946
rect 12206 29894 12258 29946
rect 16950 29894 17002 29946
rect 17014 29894 17066 29946
rect 17078 29894 17130 29946
rect 17142 29894 17194 29946
rect 17206 29894 17258 29946
rect 21950 29894 22002 29946
rect 22014 29894 22066 29946
rect 22078 29894 22130 29946
rect 22142 29894 22194 29946
rect 22206 29894 22258 29946
rect 26950 29894 27002 29946
rect 27014 29894 27066 29946
rect 27078 29894 27130 29946
rect 27142 29894 27194 29946
rect 27206 29894 27258 29946
rect 31950 29894 32002 29946
rect 32014 29894 32066 29946
rect 32078 29894 32130 29946
rect 32142 29894 32194 29946
rect 32206 29894 32258 29946
rect 36950 29894 37002 29946
rect 37014 29894 37066 29946
rect 37078 29894 37130 29946
rect 37142 29894 37194 29946
rect 37206 29894 37258 29946
rect 41950 29894 42002 29946
rect 42014 29894 42066 29946
rect 42078 29894 42130 29946
rect 42142 29894 42194 29946
rect 42206 29894 42258 29946
rect 46950 29894 47002 29946
rect 47014 29894 47066 29946
rect 47078 29894 47130 29946
rect 47142 29894 47194 29946
rect 47206 29894 47258 29946
rect 51950 29894 52002 29946
rect 52014 29894 52066 29946
rect 52078 29894 52130 29946
rect 52142 29894 52194 29946
rect 52206 29894 52258 29946
rect 56950 29894 57002 29946
rect 57014 29894 57066 29946
rect 57078 29894 57130 29946
rect 57142 29894 57194 29946
rect 57206 29894 57258 29946
rect 58532 29631 58584 29640
rect 58532 29597 58541 29631
rect 58541 29597 58575 29631
rect 58575 29597 58584 29631
rect 58532 29588 58584 29597
rect 2610 29350 2662 29402
rect 2674 29350 2726 29402
rect 2738 29350 2790 29402
rect 2802 29350 2854 29402
rect 2866 29350 2918 29402
rect 7610 29350 7662 29402
rect 7674 29350 7726 29402
rect 7738 29350 7790 29402
rect 7802 29350 7854 29402
rect 7866 29350 7918 29402
rect 12610 29350 12662 29402
rect 12674 29350 12726 29402
rect 12738 29350 12790 29402
rect 12802 29350 12854 29402
rect 12866 29350 12918 29402
rect 17610 29350 17662 29402
rect 17674 29350 17726 29402
rect 17738 29350 17790 29402
rect 17802 29350 17854 29402
rect 17866 29350 17918 29402
rect 22610 29350 22662 29402
rect 22674 29350 22726 29402
rect 22738 29350 22790 29402
rect 22802 29350 22854 29402
rect 22866 29350 22918 29402
rect 27610 29350 27662 29402
rect 27674 29350 27726 29402
rect 27738 29350 27790 29402
rect 27802 29350 27854 29402
rect 27866 29350 27918 29402
rect 32610 29350 32662 29402
rect 32674 29350 32726 29402
rect 32738 29350 32790 29402
rect 32802 29350 32854 29402
rect 32866 29350 32918 29402
rect 37610 29350 37662 29402
rect 37674 29350 37726 29402
rect 37738 29350 37790 29402
rect 37802 29350 37854 29402
rect 37866 29350 37918 29402
rect 42610 29350 42662 29402
rect 42674 29350 42726 29402
rect 42738 29350 42790 29402
rect 42802 29350 42854 29402
rect 42866 29350 42918 29402
rect 47610 29350 47662 29402
rect 47674 29350 47726 29402
rect 47738 29350 47790 29402
rect 47802 29350 47854 29402
rect 47866 29350 47918 29402
rect 52610 29350 52662 29402
rect 52674 29350 52726 29402
rect 52738 29350 52790 29402
rect 52802 29350 52854 29402
rect 52866 29350 52918 29402
rect 57610 29350 57662 29402
rect 57674 29350 57726 29402
rect 57738 29350 57790 29402
rect 57802 29350 57854 29402
rect 57866 29350 57918 29402
rect 58532 29019 58584 29028
rect 58532 28985 58541 29019
rect 58541 28985 58575 29019
rect 58575 28985 58584 29019
rect 58532 28976 58584 28985
rect 1950 28806 2002 28858
rect 2014 28806 2066 28858
rect 2078 28806 2130 28858
rect 2142 28806 2194 28858
rect 2206 28806 2258 28858
rect 6950 28806 7002 28858
rect 7014 28806 7066 28858
rect 7078 28806 7130 28858
rect 7142 28806 7194 28858
rect 7206 28806 7258 28858
rect 11950 28806 12002 28858
rect 12014 28806 12066 28858
rect 12078 28806 12130 28858
rect 12142 28806 12194 28858
rect 12206 28806 12258 28858
rect 16950 28806 17002 28858
rect 17014 28806 17066 28858
rect 17078 28806 17130 28858
rect 17142 28806 17194 28858
rect 17206 28806 17258 28858
rect 21950 28806 22002 28858
rect 22014 28806 22066 28858
rect 22078 28806 22130 28858
rect 22142 28806 22194 28858
rect 22206 28806 22258 28858
rect 26950 28806 27002 28858
rect 27014 28806 27066 28858
rect 27078 28806 27130 28858
rect 27142 28806 27194 28858
rect 27206 28806 27258 28858
rect 31950 28806 32002 28858
rect 32014 28806 32066 28858
rect 32078 28806 32130 28858
rect 32142 28806 32194 28858
rect 32206 28806 32258 28858
rect 36950 28806 37002 28858
rect 37014 28806 37066 28858
rect 37078 28806 37130 28858
rect 37142 28806 37194 28858
rect 37206 28806 37258 28858
rect 41950 28806 42002 28858
rect 42014 28806 42066 28858
rect 42078 28806 42130 28858
rect 42142 28806 42194 28858
rect 42206 28806 42258 28858
rect 46950 28806 47002 28858
rect 47014 28806 47066 28858
rect 47078 28806 47130 28858
rect 47142 28806 47194 28858
rect 47206 28806 47258 28858
rect 51950 28806 52002 28858
rect 52014 28806 52066 28858
rect 52078 28806 52130 28858
rect 52142 28806 52194 28858
rect 52206 28806 52258 28858
rect 56950 28806 57002 28858
rect 57014 28806 57066 28858
rect 57078 28806 57130 28858
rect 57142 28806 57194 28858
rect 57206 28806 57258 28858
rect 2610 28262 2662 28314
rect 2674 28262 2726 28314
rect 2738 28262 2790 28314
rect 2802 28262 2854 28314
rect 2866 28262 2918 28314
rect 7610 28262 7662 28314
rect 7674 28262 7726 28314
rect 7738 28262 7790 28314
rect 7802 28262 7854 28314
rect 7866 28262 7918 28314
rect 12610 28262 12662 28314
rect 12674 28262 12726 28314
rect 12738 28262 12790 28314
rect 12802 28262 12854 28314
rect 12866 28262 12918 28314
rect 17610 28262 17662 28314
rect 17674 28262 17726 28314
rect 17738 28262 17790 28314
rect 17802 28262 17854 28314
rect 17866 28262 17918 28314
rect 22610 28262 22662 28314
rect 22674 28262 22726 28314
rect 22738 28262 22790 28314
rect 22802 28262 22854 28314
rect 22866 28262 22918 28314
rect 27610 28262 27662 28314
rect 27674 28262 27726 28314
rect 27738 28262 27790 28314
rect 27802 28262 27854 28314
rect 27866 28262 27918 28314
rect 32610 28262 32662 28314
rect 32674 28262 32726 28314
rect 32738 28262 32790 28314
rect 32802 28262 32854 28314
rect 32866 28262 32918 28314
rect 37610 28262 37662 28314
rect 37674 28262 37726 28314
rect 37738 28262 37790 28314
rect 37802 28262 37854 28314
rect 37866 28262 37918 28314
rect 42610 28262 42662 28314
rect 42674 28262 42726 28314
rect 42738 28262 42790 28314
rect 42802 28262 42854 28314
rect 42866 28262 42918 28314
rect 47610 28262 47662 28314
rect 47674 28262 47726 28314
rect 47738 28262 47790 28314
rect 47802 28262 47854 28314
rect 47866 28262 47918 28314
rect 52610 28262 52662 28314
rect 52674 28262 52726 28314
rect 52738 28262 52790 28314
rect 52802 28262 52854 28314
rect 52866 28262 52918 28314
rect 57610 28262 57662 28314
rect 57674 28262 57726 28314
rect 57738 28262 57790 28314
rect 57802 28262 57854 28314
rect 57866 28262 57918 28314
rect 58532 27863 58584 27872
rect 58532 27829 58541 27863
rect 58541 27829 58575 27863
rect 58575 27829 58584 27863
rect 58532 27820 58584 27829
rect 1950 27718 2002 27770
rect 2014 27718 2066 27770
rect 2078 27718 2130 27770
rect 2142 27718 2194 27770
rect 2206 27718 2258 27770
rect 6950 27718 7002 27770
rect 7014 27718 7066 27770
rect 7078 27718 7130 27770
rect 7142 27718 7194 27770
rect 7206 27718 7258 27770
rect 11950 27718 12002 27770
rect 12014 27718 12066 27770
rect 12078 27718 12130 27770
rect 12142 27718 12194 27770
rect 12206 27718 12258 27770
rect 16950 27718 17002 27770
rect 17014 27718 17066 27770
rect 17078 27718 17130 27770
rect 17142 27718 17194 27770
rect 17206 27718 17258 27770
rect 21950 27718 22002 27770
rect 22014 27718 22066 27770
rect 22078 27718 22130 27770
rect 22142 27718 22194 27770
rect 22206 27718 22258 27770
rect 26950 27718 27002 27770
rect 27014 27718 27066 27770
rect 27078 27718 27130 27770
rect 27142 27718 27194 27770
rect 27206 27718 27258 27770
rect 31950 27718 32002 27770
rect 32014 27718 32066 27770
rect 32078 27718 32130 27770
rect 32142 27718 32194 27770
rect 32206 27718 32258 27770
rect 36950 27718 37002 27770
rect 37014 27718 37066 27770
rect 37078 27718 37130 27770
rect 37142 27718 37194 27770
rect 37206 27718 37258 27770
rect 41950 27718 42002 27770
rect 42014 27718 42066 27770
rect 42078 27718 42130 27770
rect 42142 27718 42194 27770
rect 42206 27718 42258 27770
rect 46950 27718 47002 27770
rect 47014 27718 47066 27770
rect 47078 27718 47130 27770
rect 47142 27718 47194 27770
rect 47206 27718 47258 27770
rect 51950 27718 52002 27770
rect 52014 27718 52066 27770
rect 52078 27718 52130 27770
rect 52142 27718 52194 27770
rect 52206 27718 52258 27770
rect 56950 27718 57002 27770
rect 57014 27718 57066 27770
rect 57078 27718 57130 27770
rect 57142 27718 57194 27770
rect 57206 27718 57258 27770
rect 58532 27455 58584 27464
rect 58532 27421 58541 27455
rect 58541 27421 58575 27455
rect 58575 27421 58584 27455
rect 58532 27412 58584 27421
rect 2610 27174 2662 27226
rect 2674 27174 2726 27226
rect 2738 27174 2790 27226
rect 2802 27174 2854 27226
rect 2866 27174 2918 27226
rect 7610 27174 7662 27226
rect 7674 27174 7726 27226
rect 7738 27174 7790 27226
rect 7802 27174 7854 27226
rect 7866 27174 7918 27226
rect 12610 27174 12662 27226
rect 12674 27174 12726 27226
rect 12738 27174 12790 27226
rect 12802 27174 12854 27226
rect 12866 27174 12918 27226
rect 17610 27174 17662 27226
rect 17674 27174 17726 27226
rect 17738 27174 17790 27226
rect 17802 27174 17854 27226
rect 17866 27174 17918 27226
rect 22610 27174 22662 27226
rect 22674 27174 22726 27226
rect 22738 27174 22790 27226
rect 22802 27174 22854 27226
rect 22866 27174 22918 27226
rect 27610 27174 27662 27226
rect 27674 27174 27726 27226
rect 27738 27174 27790 27226
rect 27802 27174 27854 27226
rect 27866 27174 27918 27226
rect 32610 27174 32662 27226
rect 32674 27174 32726 27226
rect 32738 27174 32790 27226
rect 32802 27174 32854 27226
rect 32866 27174 32918 27226
rect 37610 27174 37662 27226
rect 37674 27174 37726 27226
rect 37738 27174 37790 27226
rect 37802 27174 37854 27226
rect 37866 27174 37918 27226
rect 42610 27174 42662 27226
rect 42674 27174 42726 27226
rect 42738 27174 42790 27226
rect 42802 27174 42854 27226
rect 42866 27174 42918 27226
rect 47610 27174 47662 27226
rect 47674 27174 47726 27226
rect 47738 27174 47790 27226
rect 47802 27174 47854 27226
rect 47866 27174 47918 27226
rect 52610 27174 52662 27226
rect 52674 27174 52726 27226
rect 52738 27174 52790 27226
rect 52802 27174 52854 27226
rect 52866 27174 52918 27226
rect 57610 27174 57662 27226
rect 57674 27174 57726 27226
rect 57738 27174 57790 27226
rect 57802 27174 57854 27226
rect 57866 27174 57918 27226
rect 1950 26630 2002 26682
rect 2014 26630 2066 26682
rect 2078 26630 2130 26682
rect 2142 26630 2194 26682
rect 2206 26630 2258 26682
rect 6950 26630 7002 26682
rect 7014 26630 7066 26682
rect 7078 26630 7130 26682
rect 7142 26630 7194 26682
rect 7206 26630 7258 26682
rect 11950 26630 12002 26682
rect 12014 26630 12066 26682
rect 12078 26630 12130 26682
rect 12142 26630 12194 26682
rect 12206 26630 12258 26682
rect 16950 26630 17002 26682
rect 17014 26630 17066 26682
rect 17078 26630 17130 26682
rect 17142 26630 17194 26682
rect 17206 26630 17258 26682
rect 21950 26630 22002 26682
rect 22014 26630 22066 26682
rect 22078 26630 22130 26682
rect 22142 26630 22194 26682
rect 22206 26630 22258 26682
rect 26950 26630 27002 26682
rect 27014 26630 27066 26682
rect 27078 26630 27130 26682
rect 27142 26630 27194 26682
rect 27206 26630 27258 26682
rect 31950 26630 32002 26682
rect 32014 26630 32066 26682
rect 32078 26630 32130 26682
rect 32142 26630 32194 26682
rect 32206 26630 32258 26682
rect 36950 26630 37002 26682
rect 37014 26630 37066 26682
rect 37078 26630 37130 26682
rect 37142 26630 37194 26682
rect 37206 26630 37258 26682
rect 41950 26630 42002 26682
rect 42014 26630 42066 26682
rect 42078 26630 42130 26682
rect 42142 26630 42194 26682
rect 42206 26630 42258 26682
rect 46950 26630 47002 26682
rect 47014 26630 47066 26682
rect 47078 26630 47130 26682
rect 47142 26630 47194 26682
rect 47206 26630 47258 26682
rect 51950 26630 52002 26682
rect 52014 26630 52066 26682
rect 52078 26630 52130 26682
rect 52142 26630 52194 26682
rect 52206 26630 52258 26682
rect 56950 26630 57002 26682
rect 57014 26630 57066 26682
rect 57078 26630 57130 26682
rect 57142 26630 57194 26682
rect 57206 26630 57258 26682
rect 58348 26324 58400 26376
rect 2610 26086 2662 26138
rect 2674 26086 2726 26138
rect 2738 26086 2790 26138
rect 2802 26086 2854 26138
rect 2866 26086 2918 26138
rect 7610 26086 7662 26138
rect 7674 26086 7726 26138
rect 7738 26086 7790 26138
rect 7802 26086 7854 26138
rect 7866 26086 7918 26138
rect 12610 26086 12662 26138
rect 12674 26086 12726 26138
rect 12738 26086 12790 26138
rect 12802 26086 12854 26138
rect 12866 26086 12918 26138
rect 17610 26086 17662 26138
rect 17674 26086 17726 26138
rect 17738 26086 17790 26138
rect 17802 26086 17854 26138
rect 17866 26086 17918 26138
rect 22610 26086 22662 26138
rect 22674 26086 22726 26138
rect 22738 26086 22790 26138
rect 22802 26086 22854 26138
rect 22866 26086 22918 26138
rect 27610 26086 27662 26138
rect 27674 26086 27726 26138
rect 27738 26086 27790 26138
rect 27802 26086 27854 26138
rect 27866 26086 27918 26138
rect 32610 26086 32662 26138
rect 32674 26086 32726 26138
rect 32738 26086 32790 26138
rect 32802 26086 32854 26138
rect 32866 26086 32918 26138
rect 37610 26086 37662 26138
rect 37674 26086 37726 26138
rect 37738 26086 37790 26138
rect 37802 26086 37854 26138
rect 37866 26086 37918 26138
rect 42610 26086 42662 26138
rect 42674 26086 42726 26138
rect 42738 26086 42790 26138
rect 42802 26086 42854 26138
rect 42866 26086 42918 26138
rect 47610 26086 47662 26138
rect 47674 26086 47726 26138
rect 47738 26086 47790 26138
rect 47802 26086 47854 26138
rect 47866 26086 47918 26138
rect 52610 26086 52662 26138
rect 52674 26086 52726 26138
rect 52738 26086 52790 26138
rect 52802 26086 52854 26138
rect 52866 26086 52918 26138
rect 57610 26086 57662 26138
rect 57674 26086 57726 26138
rect 57738 26086 57790 26138
rect 57802 26086 57854 26138
rect 57866 26086 57918 26138
rect 58532 25687 58584 25696
rect 58532 25653 58541 25687
rect 58541 25653 58575 25687
rect 58575 25653 58584 25687
rect 58532 25644 58584 25653
rect 1950 25542 2002 25594
rect 2014 25542 2066 25594
rect 2078 25542 2130 25594
rect 2142 25542 2194 25594
rect 2206 25542 2258 25594
rect 6950 25542 7002 25594
rect 7014 25542 7066 25594
rect 7078 25542 7130 25594
rect 7142 25542 7194 25594
rect 7206 25542 7258 25594
rect 11950 25542 12002 25594
rect 12014 25542 12066 25594
rect 12078 25542 12130 25594
rect 12142 25542 12194 25594
rect 12206 25542 12258 25594
rect 16950 25542 17002 25594
rect 17014 25542 17066 25594
rect 17078 25542 17130 25594
rect 17142 25542 17194 25594
rect 17206 25542 17258 25594
rect 21950 25542 22002 25594
rect 22014 25542 22066 25594
rect 22078 25542 22130 25594
rect 22142 25542 22194 25594
rect 22206 25542 22258 25594
rect 26950 25542 27002 25594
rect 27014 25542 27066 25594
rect 27078 25542 27130 25594
rect 27142 25542 27194 25594
rect 27206 25542 27258 25594
rect 31950 25542 32002 25594
rect 32014 25542 32066 25594
rect 32078 25542 32130 25594
rect 32142 25542 32194 25594
rect 32206 25542 32258 25594
rect 36950 25542 37002 25594
rect 37014 25542 37066 25594
rect 37078 25542 37130 25594
rect 37142 25542 37194 25594
rect 37206 25542 37258 25594
rect 41950 25542 42002 25594
rect 42014 25542 42066 25594
rect 42078 25542 42130 25594
rect 42142 25542 42194 25594
rect 42206 25542 42258 25594
rect 46950 25542 47002 25594
rect 47014 25542 47066 25594
rect 47078 25542 47130 25594
rect 47142 25542 47194 25594
rect 47206 25542 47258 25594
rect 51950 25542 52002 25594
rect 52014 25542 52066 25594
rect 52078 25542 52130 25594
rect 52142 25542 52194 25594
rect 52206 25542 52258 25594
rect 56950 25542 57002 25594
rect 57014 25542 57066 25594
rect 57078 25542 57130 25594
rect 57142 25542 57194 25594
rect 57206 25542 57258 25594
rect 2610 24998 2662 25050
rect 2674 24998 2726 25050
rect 2738 24998 2790 25050
rect 2802 24998 2854 25050
rect 2866 24998 2918 25050
rect 7610 24998 7662 25050
rect 7674 24998 7726 25050
rect 7738 24998 7790 25050
rect 7802 24998 7854 25050
rect 7866 24998 7918 25050
rect 12610 24998 12662 25050
rect 12674 24998 12726 25050
rect 12738 24998 12790 25050
rect 12802 24998 12854 25050
rect 12866 24998 12918 25050
rect 17610 24998 17662 25050
rect 17674 24998 17726 25050
rect 17738 24998 17790 25050
rect 17802 24998 17854 25050
rect 17866 24998 17918 25050
rect 22610 24998 22662 25050
rect 22674 24998 22726 25050
rect 22738 24998 22790 25050
rect 22802 24998 22854 25050
rect 22866 24998 22918 25050
rect 27610 24998 27662 25050
rect 27674 24998 27726 25050
rect 27738 24998 27790 25050
rect 27802 24998 27854 25050
rect 27866 24998 27918 25050
rect 32610 24998 32662 25050
rect 32674 24998 32726 25050
rect 32738 24998 32790 25050
rect 32802 24998 32854 25050
rect 32866 24998 32918 25050
rect 37610 24998 37662 25050
rect 37674 24998 37726 25050
rect 37738 24998 37790 25050
rect 37802 24998 37854 25050
rect 37866 24998 37918 25050
rect 42610 24998 42662 25050
rect 42674 24998 42726 25050
rect 42738 24998 42790 25050
rect 42802 24998 42854 25050
rect 42866 24998 42918 25050
rect 47610 24998 47662 25050
rect 47674 24998 47726 25050
rect 47738 24998 47790 25050
rect 47802 24998 47854 25050
rect 47866 24998 47918 25050
rect 52610 24998 52662 25050
rect 52674 24998 52726 25050
rect 52738 24998 52790 25050
rect 52802 24998 52854 25050
rect 52866 24998 52918 25050
rect 57610 24998 57662 25050
rect 57674 24998 57726 25050
rect 57738 24998 57790 25050
rect 57802 24998 57854 25050
rect 57866 24998 57918 25050
rect 58532 24599 58584 24608
rect 58532 24565 58541 24599
rect 58541 24565 58575 24599
rect 58575 24565 58584 24599
rect 58532 24556 58584 24565
rect 1950 24454 2002 24506
rect 2014 24454 2066 24506
rect 2078 24454 2130 24506
rect 2142 24454 2194 24506
rect 2206 24454 2258 24506
rect 6950 24454 7002 24506
rect 7014 24454 7066 24506
rect 7078 24454 7130 24506
rect 7142 24454 7194 24506
rect 7206 24454 7258 24506
rect 11950 24454 12002 24506
rect 12014 24454 12066 24506
rect 12078 24454 12130 24506
rect 12142 24454 12194 24506
rect 12206 24454 12258 24506
rect 16950 24454 17002 24506
rect 17014 24454 17066 24506
rect 17078 24454 17130 24506
rect 17142 24454 17194 24506
rect 17206 24454 17258 24506
rect 21950 24454 22002 24506
rect 22014 24454 22066 24506
rect 22078 24454 22130 24506
rect 22142 24454 22194 24506
rect 22206 24454 22258 24506
rect 26950 24454 27002 24506
rect 27014 24454 27066 24506
rect 27078 24454 27130 24506
rect 27142 24454 27194 24506
rect 27206 24454 27258 24506
rect 31950 24454 32002 24506
rect 32014 24454 32066 24506
rect 32078 24454 32130 24506
rect 32142 24454 32194 24506
rect 32206 24454 32258 24506
rect 36950 24454 37002 24506
rect 37014 24454 37066 24506
rect 37078 24454 37130 24506
rect 37142 24454 37194 24506
rect 37206 24454 37258 24506
rect 41950 24454 42002 24506
rect 42014 24454 42066 24506
rect 42078 24454 42130 24506
rect 42142 24454 42194 24506
rect 42206 24454 42258 24506
rect 46950 24454 47002 24506
rect 47014 24454 47066 24506
rect 47078 24454 47130 24506
rect 47142 24454 47194 24506
rect 47206 24454 47258 24506
rect 51950 24454 52002 24506
rect 52014 24454 52066 24506
rect 52078 24454 52130 24506
rect 52142 24454 52194 24506
rect 52206 24454 52258 24506
rect 56950 24454 57002 24506
rect 57014 24454 57066 24506
rect 57078 24454 57130 24506
rect 57142 24454 57194 24506
rect 57206 24454 57258 24506
rect 58532 24191 58584 24200
rect 58532 24157 58541 24191
rect 58541 24157 58575 24191
rect 58575 24157 58584 24191
rect 58532 24148 58584 24157
rect 2610 23910 2662 23962
rect 2674 23910 2726 23962
rect 2738 23910 2790 23962
rect 2802 23910 2854 23962
rect 2866 23910 2918 23962
rect 7610 23910 7662 23962
rect 7674 23910 7726 23962
rect 7738 23910 7790 23962
rect 7802 23910 7854 23962
rect 7866 23910 7918 23962
rect 12610 23910 12662 23962
rect 12674 23910 12726 23962
rect 12738 23910 12790 23962
rect 12802 23910 12854 23962
rect 12866 23910 12918 23962
rect 17610 23910 17662 23962
rect 17674 23910 17726 23962
rect 17738 23910 17790 23962
rect 17802 23910 17854 23962
rect 17866 23910 17918 23962
rect 22610 23910 22662 23962
rect 22674 23910 22726 23962
rect 22738 23910 22790 23962
rect 22802 23910 22854 23962
rect 22866 23910 22918 23962
rect 27610 23910 27662 23962
rect 27674 23910 27726 23962
rect 27738 23910 27790 23962
rect 27802 23910 27854 23962
rect 27866 23910 27918 23962
rect 32610 23910 32662 23962
rect 32674 23910 32726 23962
rect 32738 23910 32790 23962
rect 32802 23910 32854 23962
rect 32866 23910 32918 23962
rect 37610 23910 37662 23962
rect 37674 23910 37726 23962
rect 37738 23910 37790 23962
rect 37802 23910 37854 23962
rect 37866 23910 37918 23962
rect 42610 23910 42662 23962
rect 42674 23910 42726 23962
rect 42738 23910 42790 23962
rect 42802 23910 42854 23962
rect 42866 23910 42918 23962
rect 47610 23910 47662 23962
rect 47674 23910 47726 23962
rect 47738 23910 47790 23962
rect 47802 23910 47854 23962
rect 47866 23910 47918 23962
rect 52610 23910 52662 23962
rect 52674 23910 52726 23962
rect 52738 23910 52790 23962
rect 52802 23910 52854 23962
rect 52866 23910 52918 23962
rect 57610 23910 57662 23962
rect 57674 23910 57726 23962
rect 57738 23910 57790 23962
rect 57802 23910 57854 23962
rect 57866 23910 57918 23962
rect 1950 23366 2002 23418
rect 2014 23366 2066 23418
rect 2078 23366 2130 23418
rect 2142 23366 2194 23418
rect 2206 23366 2258 23418
rect 6950 23366 7002 23418
rect 7014 23366 7066 23418
rect 7078 23366 7130 23418
rect 7142 23366 7194 23418
rect 7206 23366 7258 23418
rect 11950 23366 12002 23418
rect 12014 23366 12066 23418
rect 12078 23366 12130 23418
rect 12142 23366 12194 23418
rect 12206 23366 12258 23418
rect 16950 23366 17002 23418
rect 17014 23366 17066 23418
rect 17078 23366 17130 23418
rect 17142 23366 17194 23418
rect 17206 23366 17258 23418
rect 21950 23366 22002 23418
rect 22014 23366 22066 23418
rect 22078 23366 22130 23418
rect 22142 23366 22194 23418
rect 22206 23366 22258 23418
rect 26950 23366 27002 23418
rect 27014 23366 27066 23418
rect 27078 23366 27130 23418
rect 27142 23366 27194 23418
rect 27206 23366 27258 23418
rect 31950 23366 32002 23418
rect 32014 23366 32066 23418
rect 32078 23366 32130 23418
rect 32142 23366 32194 23418
rect 32206 23366 32258 23418
rect 36950 23366 37002 23418
rect 37014 23366 37066 23418
rect 37078 23366 37130 23418
rect 37142 23366 37194 23418
rect 37206 23366 37258 23418
rect 41950 23366 42002 23418
rect 42014 23366 42066 23418
rect 42078 23366 42130 23418
rect 42142 23366 42194 23418
rect 42206 23366 42258 23418
rect 46950 23366 47002 23418
rect 47014 23366 47066 23418
rect 47078 23366 47130 23418
rect 47142 23366 47194 23418
rect 47206 23366 47258 23418
rect 51950 23366 52002 23418
rect 52014 23366 52066 23418
rect 52078 23366 52130 23418
rect 52142 23366 52194 23418
rect 52206 23366 52258 23418
rect 56950 23366 57002 23418
rect 57014 23366 57066 23418
rect 57078 23366 57130 23418
rect 57142 23366 57194 23418
rect 57206 23366 57258 23418
rect 58532 23103 58584 23112
rect 58532 23069 58541 23103
rect 58541 23069 58575 23103
rect 58575 23069 58584 23103
rect 58532 23060 58584 23069
rect 2610 22822 2662 22874
rect 2674 22822 2726 22874
rect 2738 22822 2790 22874
rect 2802 22822 2854 22874
rect 2866 22822 2918 22874
rect 7610 22822 7662 22874
rect 7674 22822 7726 22874
rect 7738 22822 7790 22874
rect 7802 22822 7854 22874
rect 7866 22822 7918 22874
rect 12610 22822 12662 22874
rect 12674 22822 12726 22874
rect 12738 22822 12790 22874
rect 12802 22822 12854 22874
rect 12866 22822 12918 22874
rect 17610 22822 17662 22874
rect 17674 22822 17726 22874
rect 17738 22822 17790 22874
rect 17802 22822 17854 22874
rect 17866 22822 17918 22874
rect 22610 22822 22662 22874
rect 22674 22822 22726 22874
rect 22738 22822 22790 22874
rect 22802 22822 22854 22874
rect 22866 22822 22918 22874
rect 27610 22822 27662 22874
rect 27674 22822 27726 22874
rect 27738 22822 27790 22874
rect 27802 22822 27854 22874
rect 27866 22822 27918 22874
rect 32610 22822 32662 22874
rect 32674 22822 32726 22874
rect 32738 22822 32790 22874
rect 32802 22822 32854 22874
rect 32866 22822 32918 22874
rect 37610 22822 37662 22874
rect 37674 22822 37726 22874
rect 37738 22822 37790 22874
rect 37802 22822 37854 22874
rect 37866 22822 37918 22874
rect 42610 22822 42662 22874
rect 42674 22822 42726 22874
rect 42738 22822 42790 22874
rect 42802 22822 42854 22874
rect 42866 22822 42918 22874
rect 47610 22822 47662 22874
rect 47674 22822 47726 22874
rect 47738 22822 47790 22874
rect 47802 22822 47854 22874
rect 47866 22822 47918 22874
rect 52610 22822 52662 22874
rect 52674 22822 52726 22874
rect 52738 22822 52790 22874
rect 52802 22822 52854 22874
rect 52866 22822 52918 22874
rect 57610 22822 57662 22874
rect 57674 22822 57726 22874
rect 57738 22822 57790 22874
rect 57802 22822 57854 22874
rect 57866 22822 57918 22874
rect 58532 22423 58584 22432
rect 58532 22389 58541 22423
rect 58541 22389 58575 22423
rect 58575 22389 58584 22423
rect 58532 22380 58584 22389
rect 1950 22278 2002 22330
rect 2014 22278 2066 22330
rect 2078 22278 2130 22330
rect 2142 22278 2194 22330
rect 2206 22278 2258 22330
rect 6950 22278 7002 22330
rect 7014 22278 7066 22330
rect 7078 22278 7130 22330
rect 7142 22278 7194 22330
rect 7206 22278 7258 22330
rect 11950 22278 12002 22330
rect 12014 22278 12066 22330
rect 12078 22278 12130 22330
rect 12142 22278 12194 22330
rect 12206 22278 12258 22330
rect 16950 22278 17002 22330
rect 17014 22278 17066 22330
rect 17078 22278 17130 22330
rect 17142 22278 17194 22330
rect 17206 22278 17258 22330
rect 21950 22278 22002 22330
rect 22014 22278 22066 22330
rect 22078 22278 22130 22330
rect 22142 22278 22194 22330
rect 22206 22278 22258 22330
rect 26950 22278 27002 22330
rect 27014 22278 27066 22330
rect 27078 22278 27130 22330
rect 27142 22278 27194 22330
rect 27206 22278 27258 22330
rect 31950 22278 32002 22330
rect 32014 22278 32066 22330
rect 32078 22278 32130 22330
rect 32142 22278 32194 22330
rect 32206 22278 32258 22330
rect 36950 22278 37002 22330
rect 37014 22278 37066 22330
rect 37078 22278 37130 22330
rect 37142 22278 37194 22330
rect 37206 22278 37258 22330
rect 41950 22278 42002 22330
rect 42014 22278 42066 22330
rect 42078 22278 42130 22330
rect 42142 22278 42194 22330
rect 42206 22278 42258 22330
rect 46950 22278 47002 22330
rect 47014 22278 47066 22330
rect 47078 22278 47130 22330
rect 47142 22278 47194 22330
rect 47206 22278 47258 22330
rect 51950 22278 52002 22330
rect 52014 22278 52066 22330
rect 52078 22278 52130 22330
rect 52142 22278 52194 22330
rect 52206 22278 52258 22330
rect 56950 22278 57002 22330
rect 57014 22278 57066 22330
rect 57078 22278 57130 22330
rect 57142 22278 57194 22330
rect 57206 22278 57258 22330
rect 2610 21734 2662 21786
rect 2674 21734 2726 21786
rect 2738 21734 2790 21786
rect 2802 21734 2854 21786
rect 2866 21734 2918 21786
rect 7610 21734 7662 21786
rect 7674 21734 7726 21786
rect 7738 21734 7790 21786
rect 7802 21734 7854 21786
rect 7866 21734 7918 21786
rect 12610 21734 12662 21786
rect 12674 21734 12726 21786
rect 12738 21734 12790 21786
rect 12802 21734 12854 21786
rect 12866 21734 12918 21786
rect 17610 21734 17662 21786
rect 17674 21734 17726 21786
rect 17738 21734 17790 21786
rect 17802 21734 17854 21786
rect 17866 21734 17918 21786
rect 22610 21734 22662 21786
rect 22674 21734 22726 21786
rect 22738 21734 22790 21786
rect 22802 21734 22854 21786
rect 22866 21734 22918 21786
rect 27610 21734 27662 21786
rect 27674 21734 27726 21786
rect 27738 21734 27790 21786
rect 27802 21734 27854 21786
rect 27866 21734 27918 21786
rect 32610 21734 32662 21786
rect 32674 21734 32726 21786
rect 32738 21734 32790 21786
rect 32802 21734 32854 21786
rect 32866 21734 32918 21786
rect 37610 21734 37662 21786
rect 37674 21734 37726 21786
rect 37738 21734 37790 21786
rect 37802 21734 37854 21786
rect 37866 21734 37918 21786
rect 42610 21734 42662 21786
rect 42674 21734 42726 21786
rect 42738 21734 42790 21786
rect 42802 21734 42854 21786
rect 42866 21734 42918 21786
rect 47610 21734 47662 21786
rect 47674 21734 47726 21786
rect 47738 21734 47790 21786
rect 47802 21734 47854 21786
rect 47866 21734 47918 21786
rect 52610 21734 52662 21786
rect 52674 21734 52726 21786
rect 52738 21734 52790 21786
rect 52802 21734 52854 21786
rect 52866 21734 52918 21786
rect 57610 21734 57662 21786
rect 57674 21734 57726 21786
rect 57738 21734 57790 21786
rect 57802 21734 57854 21786
rect 57866 21734 57918 21786
rect 58532 21335 58584 21344
rect 58532 21301 58541 21335
rect 58541 21301 58575 21335
rect 58575 21301 58584 21335
rect 58532 21292 58584 21301
rect 1950 21190 2002 21242
rect 2014 21190 2066 21242
rect 2078 21190 2130 21242
rect 2142 21190 2194 21242
rect 2206 21190 2258 21242
rect 6950 21190 7002 21242
rect 7014 21190 7066 21242
rect 7078 21190 7130 21242
rect 7142 21190 7194 21242
rect 7206 21190 7258 21242
rect 11950 21190 12002 21242
rect 12014 21190 12066 21242
rect 12078 21190 12130 21242
rect 12142 21190 12194 21242
rect 12206 21190 12258 21242
rect 16950 21190 17002 21242
rect 17014 21190 17066 21242
rect 17078 21190 17130 21242
rect 17142 21190 17194 21242
rect 17206 21190 17258 21242
rect 21950 21190 22002 21242
rect 22014 21190 22066 21242
rect 22078 21190 22130 21242
rect 22142 21190 22194 21242
rect 22206 21190 22258 21242
rect 26950 21190 27002 21242
rect 27014 21190 27066 21242
rect 27078 21190 27130 21242
rect 27142 21190 27194 21242
rect 27206 21190 27258 21242
rect 31950 21190 32002 21242
rect 32014 21190 32066 21242
rect 32078 21190 32130 21242
rect 32142 21190 32194 21242
rect 32206 21190 32258 21242
rect 36950 21190 37002 21242
rect 37014 21190 37066 21242
rect 37078 21190 37130 21242
rect 37142 21190 37194 21242
rect 37206 21190 37258 21242
rect 41950 21190 42002 21242
rect 42014 21190 42066 21242
rect 42078 21190 42130 21242
rect 42142 21190 42194 21242
rect 42206 21190 42258 21242
rect 46950 21190 47002 21242
rect 47014 21190 47066 21242
rect 47078 21190 47130 21242
rect 47142 21190 47194 21242
rect 47206 21190 47258 21242
rect 51950 21190 52002 21242
rect 52014 21190 52066 21242
rect 52078 21190 52130 21242
rect 52142 21190 52194 21242
rect 52206 21190 52258 21242
rect 56950 21190 57002 21242
rect 57014 21190 57066 21242
rect 57078 21190 57130 21242
rect 57142 21190 57194 21242
rect 57206 21190 57258 21242
rect 58532 20927 58584 20936
rect 58532 20893 58541 20927
rect 58541 20893 58575 20927
rect 58575 20893 58584 20927
rect 58532 20884 58584 20893
rect 2610 20646 2662 20698
rect 2674 20646 2726 20698
rect 2738 20646 2790 20698
rect 2802 20646 2854 20698
rect 2866 20646 2918 20698
rect 7610 20646 7662 20698
rect 7674 20646 7726 20698
rect 7738 20646 7790 20698
rect 7802 20646 7854 20698
rect 7866 20646 7918 20698
rect 12610 20646 12662 20698
rect 12674 20646 12726 20698
rect 12738 20646 12790 20698
rect 12802 20646 12854 20698
rect 12866 20646 12918 20698
rect 17610 20646 17662 20698
rect 17674 20646 17726 20698
rect 17738 20646 17790 20698
rect 17802 20646 17854 20698
rect 17866 20646 17918 20698
rect 22610 20646 22662 20698
rect 22674 20646 22726 20698
rect 22738 20646 22790 20698
rect 22802 20646 22854 20698
rect 22866 20646 22918 20698
rect 27610 20646 27662 20698
rect 27674 20646 27726 20698
rect 27738 20646 27790 20698
rect 27802 20646 27854 20698
rect 27866 20646 27918 20698
rect 32610 20646 32662 20698
rect 32674 20646 32726 20698
rect 32738 20646 32790 20698
rect 32802 20646 32854 20698
rect 32866 20646 32918 20698
rect 37610 20646 37662 20698
rect 37674 20646 37726 20698
rect 37738 20646 37790 20698
rect 37802 20646 37854 20698
rect 37866 20646 37918 20698
rect 42610 20646 42662 20698
rect 42674 20646 42726 20698
rect 42738 20646 42790 20698
rect 42802 20646 42854 20698
rect 42866 20646 42918 20698
rect 47610 20646 47662 20698
rect 47674 20646 47726 20698
rect 47738 20646 47790 20698
rect 47802 20646 47854 20698
rect 47866 20646 47918 20698
rect 52610 20646 52662 20698
rect 52674 20646 52726 20698
rect 52738 20646 52790 20698
rect 52802 20646 52854 20698
rect 52866 20646 52918 20698
rect 57610 20646 57662 20698
rect 57674 20646 57726 20698
rect 57738 20646 57790 20698
rect 57802 20646 57854 20698
rect 57866 20646 57918 20698
rect 1950 20102 2002 20154
rect 2014 20102 2066 20154
rect 2078 20102 2130 20154
rect 2142 20102 2194 20154
rect 2206 20102 2258 20154
rect 6950 20102 7002 20154
rect 7014 20102 7066 20154
rect 7078 20102 7130 20154
rect 7142 20102 7194 20154
rect 7206 20102 7258 20154
rect 11950 20102 12002 20154
rect 12014 20102 12066 20154
rect 12078 20102 12130 20154
rect 12142 20102 12194 20154
rect 12206 20102 12258 20154
rect 16950 20102 17002 20154
rect 17014 20102 17066 20154
rect 17078 20102 17130 20154
rect 17142 20102 17194 20154
rect 17206 20102 17258 20154
rect 21950 20102 22002 20154
rect 22014 20102 22066 20154
rect 22078 20102 22130 20154
rect 22142 20102 22194 20154
rect 22206 20102 22258 20154
rect 26950 20102 27002 20154
rect 27014 20102 27066 20154
rect 27078 20102 27130 20154
rect 27142 20102 27194 20154
rect 27206 20102 27258 20154
rect 31950 20102 32002 20154
rect 32014 20102 32066 20154
rect 32078 20102 32130 20154
rect 32142 20102 32194 20154
rect 32206 20102 32258 20154
rect 36950 20102 37002 20154
rect 37014 20102 37066 20154
rect 37078 20102 37130 20154
rect 37142 20102 37194 20154
rect 37206 20102 37258 20154
rect 41950 20102 42002 20154
rect 42014 20102 42066 20154
rect 42078 20102 42130 20154
rect 42142 20102 42194 20154
rect 42206 20102 42258 20154
rect 46950 20102 47002 20154
rect 47014 20102 47066 20154
rect 47078 20102 47130 20154
rect 47142 20102 47194 20154
rect 47206 20102 47258 20154
rect 51950 20102 52002 20154
rect 52014 20102 52066 20154
rect 52078 20102 52130 20154
rect 52142 20102 52194 20154
rect 52206 20102 52258 20154
rect 56950 20102 57002 20154
rect 57014 20102 57066 20154
rect 57078 20102 57130 20154
rect 57142 20102 57194 20154
rect 57206 20102 57258 20154
rect 58532 19839 58584 19848
rect 58532 19805 58541 19839
rect 58541 19805 58575 19839
rect 58575 19805 58584 19839
rect 58532 19796 58584 19805
rect 2610 19558 2662 19610
rect 2674 19558 2726 19610
rect 2738 19558 2790 19610
rect 2802 19558 2854 19610
rect 2866 19558 2918 19610
rect 7610 19558 7662 19610
rect 7674 19558 7726 19610
rect 7738 19558 7790 19610
rect 7802 19558 7854 19610
rect 7866 19558 7918 19610
rect 12610 19558 12662 19610
rect 12674 19558 12726 19610
rect 12738 19558 12790 19610
rect 12802 19558 12854 19610
rect 12866 19558 12918 19610
rect 17610 19558 17662 19610
rect 17674 19558 17726 19610
rect 17738 19558 17790 19610
rect 17802 19558 17854 19610
rect 17866 19558 17918 19610
rect 22610 19558 22662 19610
rect 22674 19558 22726 19610
rect 22738 19558 22790 19610
rect 22802 19558 22854 19610
rect 22866 19558 22918 19610
rect 27610 19558 27662 19610
rect 27674 19558 27726 19610
rect 27738 19558 27790 19610
rect 27802 19558 27854 19610
rect 27866 19558 27918 19610
rect 32610 19558 32662 19610
rect 32674 19558 32726 19610
rect 32738 19558 32790 19610
rect 32802 19558 32854 19610
rect 32866 19558 32918 19610
rect 37610 19558 37662 19610
rect 37674 19558 37726 19610
rect 37738 19558 37790 19610
rect 37802 19558 37854 19610
rect 37866 19558 37918 19610
rect 42610 19558 42662 19610
rect 42674 19558 42726 19610
rect 42738 19558 42790 19610
rect 42802 19558 42854 19610
rect 42866 19558 42918 19610
rect 47610 19558 47662 19610
rect 47674 19558 47726 19610
rect 47738 19558 47790 19610
rect 47802 19558 47854 19610
rect 47866 19558 47918 19610
rect 52610 19558 52662 19610
rect 52674 19558 52726 19610
rect 52738 19558 52790 19610
rect 52802 19558 52854 19610
rect 52866 19558 52918 19610
rect 57610 19558 57662 19610
rect 57674 19558 57726 19610
rect 57738 19558 57790 19610
rect 57802 19558 57854 19610
rect 57866 19558 57918 19610
rect 58532 19159 58584 19168
rect 58532 19125 58541 19159
rect 58541 19125 58575 19159
rect 58575 19125 58584 19159
rect 58532 19116 58584 19125
rect 1950 19014 2002 19066
rect 2014 19014 2066 19066
rect 2078 19014 2130 19066
rect 2142 19014 2194 19066
rect 2206 19014 2258 19066
rect 6950 19014 7002 19066
rect 7014 19014 7066 19066
rect 7078 19014 7130 19066
rect 7142 19014 7194 19066
rect 7206 19014 7258 19066
rect 11950 19014 12002 19066
rect 12014 19014 12066 19066
rect 12078 19014 12130 19066
rect 12142 19014 12194 19066
rect 12206 19014 12258 19066
rect 16950 19014 17002 19066
rect 17014 19014 17066 19066
rect 17078 19014 17130 19066
rect 17142 19014 17194 19066
rect 17206 19014 17258 19066
rect 21950 19014 22002 19066
rect 22014 19014 22066 19066
rect 22078 19014 22130 19066
rect 22142 19014 22194 19066
rect 22206 19014 22258 19066
rect 26950 19014 27002 19066
rect 27014 19014 27066 19066
rect 27078 19014 27130 19066
rect 27142 19014 27194 19066
rect 27206 19014 27258 19066
rect 31950 19014 32002 19066
rect 32014 19014 32066 19066
rect 32078 19014 32130 19066
rect 32142 19014 32194 19066
rect 32206 19014 32258 19066
rect 36950 19014 37002 19066
rect 37014 19014 37066 19066
rect 37078 19014 37130 19066
rect 37142 19014 37194 19066
rect 37206 19014 37258 19066
rect 41950 19014 42002 19066
rect 42014 19014 42066 19066
rect 42078 19014 42130 19066
rect 42142 19014 42194 19066
rect 42206 19014 42258 19066
rect 46950 19014 47002 19066
rect 47014 19014 47066 19066
rect 47078 19014 47130 19066
rect 47142 19014 47194 19066
rect 47206 19014 47258 19066
rect 51950 19014 52002 19066
rect 52014 19014 52066 19066
rect 52078 19014 52130 19066
rect 52142 19014 52194 19066
rect 52206 19014 52258 19066
rect 56950 19014 57002 19066
rect 57014 19014 57066 19066
rect 57078 19014 57130 19066
rect 57142 19014 57194 19066
rect 57206 19014 57258 19066
rect 2610 18470 2662 18522
rect 2674 18470 2726 18522
rect 2738 18470 2790 18522
rect 2802 18470 2854 18522
rect 2866 18470 2918 18522
rect 7610 18470 7662 18522
rect 7674 18470 7726 18522
rect 7738 18470 7790 18522
rect 7802 18470 7854 18522
rect 7866 18470 7918 18522
rect 12610 18470 12662 18522
rect 12674 18470 12726 18522
rect 12738 18470 12790 18522
rect 12802 18470 12854 18522
rect 12866 18470 12918 18522
rect 17610 18470 17662 18522
rect 17674 18470 17726 18522
rect 17738 18470 17790 18522
rect 17802 18470 17854 18522
rect 17866 18470 17918 18522
rect 22610 18470 22662 18522
rect 22674 18470 22726 18522
rect 22738 18470 22790 18522
rect 22802 18470 22854 18522
rect 22866 18470 22918 18522
rect 27610 18470 27662 18522
rect 27674 18470 27726 18522
rect 27738 18470 27790 18522
rect 27802 18470 27854 18522
rect 27866 18470 27918 18522
rect 32610 18470 32662 18522
rect 32674 18470 32726 18522
rect 32738 18470 32790 18522
rect 32802 18470 32854 18522
rect 32866 18470 32918 18522
rect 37610 18470 37662 18522
rect 37674 18470 37726 18522
rect 37738 18470 37790 18522
rect 37802 18470 37854 18522
rect 37866 18470 37918 18522
rect 42610 18470 42662 18522
rect 42674 18470 42726 18522
rect 42738 18470 42790 18522
rect 42802 18470 42854 18522
rect 42866 18470 42918 18522
rect 47610 18470 47662 18522
rect 47674 18470 47726 18522
rect 47738 18470 47790 18522
rect 47802 18470 47854 18522
rect 47866 18470 47918 18522
rect 52610 18470 52662 18522
rect 52674 18470 52726 18522
rect 52738 18470 52790 18522
rect 52802 18470 52854 18522
rect 52866 18470 52918 18522
rect 57610 18470 57662 18522
rect 57674 18470 57726 18522
rect 57738 18470 57790 18522
rect 57802 18470 57854 18522
rect 57866 18470 57918 18522
rect 58532 18071 58584 18080
rect 58532 18037 58541 18071
rect 58541 18037 58575 18071
rect 58575 18037 58584 18071
rect 58532 18028 58584 18037
rect 1950 17926 2002 17978
rect 2014 17926 2066 17978
rect 2078 17926 2130 17978
rect 2142 17926 2194 17978
rect 2206 17926 2258 17978
rect 6950 17926 7002 17978
rect 7014 17926 7066 17978
rect 7078 17926 7130 17978
rect 7142 17926 7194 17978
rect 7206 17926 7258 17978
rect 11950 17926 12002 17978
rect 12014 17926 12066 17978
rect 12078 17926 12130 17978
rect 12142 17926 12194 17978
rect 12206 17926 12258 17978
rect 16950 17926 17002 17978
rect 17014 17926 17066 17978
rect 17078 17926 17130 17978
rect 17142 17926 17194 17978
rect 17206 17926 17258 17978
rect 21950 17926 22002 17978
rect 22014 17926 22066 17978
rect 22078 17926 22130 17978
rect 22142 17926 22194 17978
rect 22206 17926 22258 17978
rect 26950 17926 27002 17978
rect 27014 17926 27066 17978
rect 27078 17926 27130 17978
rect 27142 17926 27194 17978
rect 27206 17926 27258 17978
rect 31950 17926 32002 17978
rect 32014 17926 32066 17978
rect 32078 17926 32130 17978
rect 32142 17926 32194 17978
rect 32206 17926 32258 17978
rect 36950 17926 37002 17978
rect 37014 17926 37066 17978
rect 37078 17926 37130 17978
rect 37142 17926 37194 17978
rect 37206 17926 37258 17978
rect 41950 17926 42002 17978
rect 42014 17926 42066 17978
rect 42078 17926 42130 17978
rect 42142 17926 42194 17978
rect 42206 17926 42258 17978
rect 46950 17926 47002 17978
rect 47014 17926 47066 17978
rect 47078 17926 47130 17978
rect 47142 17926 47194 17978
rect 47206 17926 47258 17978
rect 51950 17926 52002 17978
rect 52014 17926 52066 17978
rect 52078 17926 52130 17978
rect 52142 17926 52194 17978
rect 52206 17926 52258 17978
rect 56950 17926 57002 17978
rect 57014 17926 57066 17978
rect 57078 17926 57130 17978
rect 57142 17926 57194 17978
rect 57206 17926 57258 17978
rect 58532 17663 58584 17672
rect 58532 17629 58541 17663
rect 58541 17629 58575 17663
rect 58575 17629 58584 17663
rect 58532 17620 58584 17629
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 22610 17382 22662 17434
rect 22674 17382 22726 17434
rect 22738 17382 22790 17434
rect 22802 17382 22854 17434
rect 22866 17382 22918 17434
rect 27610 17382 27662 17434
rect 27674 17382 27726 17434
rect 27738 17382 27790 17434
rect 27802 17382 27854 17434
rect 27866 17382 27918 17434
rect 32610 17382 32662 17434
rect 32674 17382 32726 17434
rect 32738 17382 32790 17434
rect 32802 17382 32854 17434
rect 32866 17382 32918 17434
rect 37610 17382 37662 17434
rect 37674 17382 37726 17434
rect 37738 17382 37790 17434
rect 37802 17382 37854 17434
rect 37866 17382 37918 17434
rect 42610 17382 42662 17434
rect 42674 17382 42726 17434
rect 42738 17382 42790 17434
rect 42802 17382 42854 17434
rect 42866 17382 42918 17434
rect 47610 17382 47662 17434
rect 47674 17382 47726 17434
rect 47738 17382 47790 17434
rect 47802 17382 47854 17434
rect 47866 17382 47918 17434
rect 52610 17382 52662 17434
rect 52674 17382 52726 17434
rect 52738 17382 52790 17434
rect 52802 17382 52854 17434
rect 52866 17382 52918 17434
rect 57610 17382 57662 17434
rect 57674 17382 57726 17434
rect 57738 17382 57790 17434
rect 57802 17382 57854 17434
rect 57866 17382 57918 17434
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 21950 16838 22002 16890
rect 22014 16838 22066 16890
rect 22078 16838 22130 16890
rect 22142 16838 22194 16890
rect 22206 16838 22258 16890
rect 26950 16838 27002 16890
rect 27014 16838 27066 16890
rect 27078 16838 27130 16890
rect 27142 16838 27194 16890
rect 27206 16838 27258 16890
rect 31950 16838 32002 16890
rect 32014 16838 32066 16890
rect 32078 16838 32130 16890
rect 32142 16838 32194 16890
rect 32206 16838 32258 16890
rect 36950 16838 37002 16890
rect 37014 16838 37066 16890
rect 37078 16838 37130 16890
rect 37142 16838 37194 16890
rect 37206 16838 37258 16890
rect 41950 16838 42002 16890
rect 42014 16838 42066 16890
rect 42078 16838 42130 16890
rect 42142 16838 42194 16890
rect 42206 16838 42258 16890
rect 46950 16838 47002 16890
rect 47014 16838 47066 16890
rect 47078 16838 47130 16890
rect 47142 16838 47194 16890
rect 47206 16838 47258 16890
rect 51950 16838 52002 16890
rect 52014 16838 52066 16890
rect 52078 16838 52130 16890
rect 52142 16838 52194 16890
rect 52206 16838 52258 16890
rect 56950 16838 57002 16890
rect 57014 16838 57066 16890
rect 57078 16838 57130 16890
rect 57142 16838 57194 16890
rect 57206 16838 57258 16890
rect 57980 16600 58032 16652
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 22610 16294 22662 16346
rect 22674 16294 22726 16346
rect 22738 16294 22790 16346
rect 22802 16294 22854 16346
rect 22866 16294 22918 16346
rect 27610 16294 27662 16346
rect 27674 16294 27726 16346
rect 27738 16294 27790 16346
rect 27802 16294 27854 16346
rect 27866 16294 27918 16346
rect 32610 16294 32662 16346
rect 32674 16294 32726 16346
rect 32738 16294 32790 16346
rect 32802 16294 32854 16346
rect 32866 16294 32918 16346
rect 37610 16294 37662 16346
rect 37674 16294 37726 16346
rect 37738 16294 37790 16346
rect 37802 16294 37854 16346
rect 37866 16294 37918 16346
rect 42610 16294 42662 16346
rect 42674 16294 42726 16346
rect 42738 16294 42790 16346
rect 42802 16294 42854 16346
rect 42866 16294 42918 16346
rect 47610 16294 47662 16346
rect 47674 16294 47726 16346
rect 47738 16294 47790 16346
rect 47802 16294 47854 16346
rect 47866 16294 47918 16346
rect 52610 16294 52662 16346
rect 52674 16294 52726 16346
rect 52738 16294 52790 16346
rect 52802 16294 52854 16346
rect 52866 16294 52918 16346
rect 57610 16294 57662 16346
rect 57674 16294 57726 16346
rect 57738 16294 57790 16346
rect 57802 16294 57854 16346
rect 57866 16294 57918 16346
rect 58532 15895 58584 15904
rect 58532 15861 58541 15895
rect 58541 15861 58575 15895
rect 58575 15861 58584 15895
rect 58532 15852 58584 15861
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 21950 15750 22002 15802
rect 22014 15750 22066 15802
rect 22078 15750 22130 15802
rect 22142 15750 22194 15802
rect 22206 15750 22258 15802
rect 26950 15750 27002 15802
rect 27014 15750 27066 15802
rect 27078 15750 27130 15802
rect 27142 15750 27194 15802
rect 27206 15750 27258 15802
rect 31950 15750 32002 15802
rect 32014 15750 32066 15802
rect 32078 15750 32130 15802
rect 32142 15750 32194 15802
rect 32206 15750 32258 15802
rect 36950 15750 37002 15802
rect 37014 15750 37066 15802
rect 37078 15750 37130 15802
rect 37142 15750 37194 15802
rect 37206 15750 37258 15802
rect 41950 15750 42002 15802
rect 42014 15750 42066 15802
rect 42078 15750 42130 15802
rect 42142 15750 42194 15802
rect 42206 15750 42258 15802
rect 46950 15750 47002 15802
rect 47014 15750 47066 15802
rect 47078 15750 47130 15802
rect 47142 15750 47194 15802
rect 47206 15750 47258 15802
rect 51950 15750 52002 15802
rect 52014 15750 52066 15802
rect 52078 15750 52130 15802
rect 52142 15750 52194 15802
rect 52206 15750 52258 15802
rect 56950 15750 57002 15802
rect 57014 15750 57066 15802
rect 57078 15750 57130 15802
rect 57142 15750 57194 15802
rect 57206 15750 57258 15802
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 22610 15206 22662 15258
rect 22674 15206 22726 15258
rect 22738 15206 22790 15258
rect 22802 15206 22854 15258
rect 22866 15206 22918 15258
rect 27610 15206 27662 15258
rect 27674 15206 27726 15258
rect 27738 15206 27790 15258
rect 27802 15206 27854 15258
rect 27866 15206 27918 15258
rect 32610 15206 32662 15258
rect 32674 15206 32726 15258
rect 32738 15206 32790 15258
rect 32802 15206 32854 15258
rect 32866 15206 32918 15258
rect 37610 15206 37662 15258
rect 37674 15206 37726 15258
rect 37738 15206 37790 15258
rect 37802 15206 37854 15258
rect 37866 15206 37918 15258
rect 42610 15206 42662 15258
rect 42674 15206 42726 15258
rect 42738 15206 42790 15258
rect 42802 15206 42854 15258
rect 42866 15206 42918 15258
rect 47610 15206 47662 15258
rect 47674 15206 47726 15258
rect 47738 15206 47790 15258
rect 47802 15206 47854 15258
rect 47866 15206 47918 15258
rect 52610 15206 52662 15258
rect 52674 15206 52726 15258
rect 52738 15206 52790 15258
rect 52802 15206 52854 15258
rect 52866 15206 52918 15258
rect 57610 15206 57662 15258
rect 57674 15206 57726 15258
rect 57738 15206 57790 15258
rect 57802 15206 57854 15258
rect 57866 15206 57918 15258
rect 58532 14807 58584 14816
rect 58532 14773 58541 14807
rect 58541 14773 58575 14807
rect 58575 14773 58584 14807
rect 58532 14764 58584 14773
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 21950 14662 22002 14714
rect 22014 14662 22066 14714
rect 22078 14662 22130 14714
rect 22142 14662 22194 14714
rect 22206 14662 22258 14714
rect 26950 14662 27002 14714
rect 27014 14662 27066 14714
rect 27078 14662 27130 14714
rect 27142 14662 27194 14714
rect 27206 14662 27258 14714
rect 31950 14662 32002 14714
rect 32014 14662 32066 14714
rect 32078 14662 32130 14714
rect 32142 14662 32194 14714
rect 32206 14662 32258 14714
rect 36950 14662 37002 14714
rect 37014 14662 37066 14714
rect 37078 14662 37130 14714
rect 37142 14662 37194 14714
rect 37206 14662 37258 14714
rect 41950 14662 42002 14714
rect 42014 14662 42066 14714
rect 42078 14662 42130 14714
rect 42142 14662 42194 14714
rect 42206 14662 42258 14714
rect 46950 14662 47002 14714
rect 47014 14662 47066 14714
rect 47078 14662 47130 14714
rect 47142 14662 47194 14714
rect 47206 14662 47258 14714
rect 51950 14662 52002 14714
rect 52014 14662 52066 14714
rect 52078 14662 52130 14714
rect 52142 14662 52194 14714
rect 52206 14662 52258 14714
rect 56950 14662 57002 14714
rect 57014 14662 57066 14714
rect 57078 14662 57130 14714
rect 57142 14662 57194 14714
rect 57206 14662 57258 14714
rect 58532 14399 58584 14408
rect 58532 14365 58541 14399
rect 58541 14365 58575 14399
rect 58575 14365 58584 14399
rect 58532 14356 58584 14365
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 22610 14118 22662 14170
rect 22674 14118 22726 14170
rect 22738 14118 22790 14170
rect 22802 14118 22854 14170
rect 22866 14118 22918 14170
rect 27610 14118 27662 14170
rect 27674 14118 27726 14170
rect 27738 14118 27790 14170
rect 27802 14118 27854 14170
rect 27866 14118 27918 14170
rect 32610 14118 32662 14170
rect 32674 14118 32726 14170
rect 32738 14118 32790 14170
rect 32802 14118 32854 14170
rect 32866 14118 32918 14170
rect 37610 14118 37662 14170
rect 37674 14118 37726 14170
rect 37738 14118 37790 14170
rect 37802 14118 37854 14170
rect 37866 14118 37918 14170
rect 42610 14118 42662 14170
rect 42674 14118 42726 14170
rect 42738 14118 42790 14170
rect 42802 14118 42854 14170
rect 42866 14118 42918 14170
rect 47610 14118 47662 14170
rect 47674 14118 47726 14170
rect 47738 14118 47790 14170
rect 47802 14118 47854 14170
rect 47866 14118 47918 14170
rect 52610 14118 52662 14170
rect 52674 14118 52726 14170
rect 52738 14118 52790 14170
rect 52802 14118 52854 14170
rect 52866 14118 52918 14170
rect 57610 14118 57662 14170
rect 57674 14118 57726 14170
rect 57738 14118 57790 14170
rect 57802 14118 57854 14170
rect 57866 14118 57918 14170
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 21950 13574 22002 13626
rect 22014 13574 22066 13626
rect 22078 13574 22130 13626
rect 22142 13574 22194 13626
rect 22206 13574 22258 13626
rect 26950 13574 27002 13626
rect 27014 13574 27066 13626
rect 27078 13574 27130 13626
rect 27142 13574 27194 13626
rect 27206 13574 27258 13626
rect 31950 13574 32002 13626
rect 32014 13574 32066 13626
rect 32078 13574 32130 13626
rect 32142 13574 32194 13626
rect 32206 13574 32258 13626
rect 36950 13574 37002 13626
rect 37014 13574 37066 13626
rect 37078 13574 37130 13626
rect 37142 13574 37194 13626
rect 37206 13574 37258 13626
rect 41950 13574 42002 13626
rect 42014 13574 42066 13626
rect 42078 13574 42130 13626
rect 42142 13574 42194 13626
rect 42206 13574 42258 13626
rect 46950 13574 47002 13626
rect 47014 13574 47066 13626
rect 47078 13574 47130 13626
rect 47142 13574 47194 13626
rect 47206 13574 47258 13626
rect 51950 13574 52002 13626
rect 52014 13574 52066 13626
rect 52078 13574 52130 13626
rect 52142 13574 52194 13626
rect 52206 13574 52258 13626
rect 56950 13574 57002 13626
rect 57014 13574 57066 13626
rect 57078 13574 57130 13626
rect 57142 13574 57194 13626
rect 57206 13574 57258 13626
rect 58532 13311 58584 13320
rect 58532 13277 58541 13311
rect 58541 13277 58575 13311
rect 58575 13277 58584 13311
rect 58532 13268 58584 13277
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 22610 13030 22662 13082
rect 22674 13030 22726 13082
rect 22738 13030 22790 13082
rect 22802 13030 22854 13082
rect 22866 13030 22918 13082
rect 27610 13030 27662 13082
rect 27674 13030 27726 13082
rect 27738 13030 27790 13082
rect 27802 13030 27854 13082
rect 27866 13030 27918 13082
rect 32610 13030 32662 13082
rect 32674 13030 32726 13082
rect 32738 13030 32790 13082
rect 32802 13030 32854 13082
rect 32866 13030 32918 13082
rect 37610 13030 37662 13082
rect 37674 13030 37726 13082
rect 37738 13030 37790 13082
rect 37802 13030 37854 13082
rect 37866 13030 37918 13082
rect 42610 13030 42662 13082
rect 42674 13030 42726 13082
rect 42738 13030 42790 13082
rect 42802 13030 42854 13082
rect 42866 13030 42918 13082
rect 47610 13030 47662 13082
rect 47674 13030 47726 13082
rect 47738 13030 47790 13082
rect 47802 13030 47854 13082
rect 47866 13030 47918 13082
rect 52610 13030 52662 13082
rect 52674 13030 52726 13082
rect 52738 13030 52790 13082
rect 52802 13030 52854 13082
rect 52866 13030 52918 13082
rect 57610 13030 57662 13082
rect 57674 13030 57726 13082
rect 57738 13030 57790 13082
rect 57802 13030 57854 13082
rect 57866 13030 57918 13082
rect 58532 12631 58584 12640
rect 58532 12597 58541 12631
rect 58541 12597 58575 12631
rect 58575 12597 58584 12631
rect 58532 12588 58584 12597
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 21950 12486 22002 12538
rect 22014 12486 22066 12538
rect 22078 12486 22130 12538
rect 22142 12486 22194 12538
rect 22206 12486 22258 12538
rect 26950 12486 27002 12538
rect 27014 12486 27066 12538
rect 27078 12486 27130 12538
rect 27142 12486 27194 12538
rect 27206 12486 27258 12538
rect 31950 12486 32002 12538
rect 32014 12486 32066 12538
rect 32078 12486 32130 12538
rect 32142 12486 32194 12538
rect 32206 12486 32258 12538
rect 36950 12486 37002 12538
rect 37014 12486 37066 12538
rect 37078 12486 37130 12538
rect 37142 12486 37194 12538
rect 37206 12486 37258 12538
rect 41950 12486 42002 12538
rect 42014 12486 42066 12538
rect 42078 12486 42130 12538
rect 42142 12486 42194 12538
rect 42206 12486 42258 12538
rect 46950 12486 47002 12538
rect 47014 12486 47066 12538
rect 47078 12486 47130 12538
rect 47142 12486 47194 12538
rect 47206 12486 47258 12538
rect 51950 12486 52002 12538
rect 52014 12486 52066 12538
rect 52078 12486 52130 12538
rect 52142 12486 52194 12538
rect 52206 12486 52258 12538
rect 56950 12486 57002 12538
rect 57014 12486 57066 12538
rect 57078 12486 57130 12538
rect 57142 12486 57194 12538
rect 57206 12486 57258 12538
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 22610 11942 22662 11994
rect 22674 11942 22726 11994
rect 22738 11942 22790 11994
rect 22802 11942 22854 11994
rect 22866 11942 22918 11994
rect 27610 11942 27662 11994
rect 27674 11942 27726 11994
rect 27738 11942 27790 11994
rect 27802 11942 27854 11994
rect 27866 11942 27918 11994
rect 32610 11942 32662 11994
rect 32674 11942 32726 11994
rect 32738 11942 32790 11994
rect 32802 11942 32854 11994
rect 32866 11942 32918 11994
rect 37610 11942 37662 11994
rect 37674 11942 37726 11994
rect 37738 11942 37790 11994
rect 37802 11942 37854 11994
rect 37866 11942 37918 11994
rect 42610 11942 42662 11994
rect 42674 11942 42726 11994
rect 42738 11942 42790 11994
rect 42802 11942 42854 11994
rect 42866 11942 42918 11994
rect 47610 11942 47662 11994
rect 47674 11942 47726 11994
rect 47738 11942 47790 11994
rect 47802 11942 47854 11994
rect 47866 11942 47918 11994
rect 52610 11942 52662 11994
rect 52674 11942 52726 11994
rect 52738 11942 52790 11994
rect 52802 11942 52854 11994
rect 52866 11942 52918 11994
rect 57610 11942 57662 11994
rect 57674 11942 57726 11994
rect 57738 11942 57790 11994
rect 57802 11942 57854 11994
rect 57866 11942 57918 11994
rect 58532 11543 58584 11552
rect 58532 11509 58541 11543
rect 58541 11509 58575 11543
rect 58575 11509 58584 11543
rect 58532 11500 58584 11509
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 21950 11398 22002 11450
rect 22014 11398 22066 11450
rect 22078 11398 22130 11450
rect 22142 11398 22194 11450
rect 22206 11398 22258 11450
rect 26950 11398 27002 11450
rect 27014 11398 27066 11450
rect 27078 11398 27130 11450
rect 27142 11398 27194 11450
rect 27206 11398 27258 11450
rect 31950 11398 32002 11450
rect 32014 11398 32066 11450
rect 32078 11398 32130 11450
rect 32142 11398 32194 11450
rect 32206 11398 32258 11450
rect 36950 11398 37002 11450
rect 37014 11398 37066 11450
rect 37078 11398 37130 11450
rect 37142 11398 37194 11450
rect 37206 11398 37258 11450
rect 41950 11398 42002 11450
rect 42014 11398 42066 11450
rect 42078 11398 42130 11450
rect 42142 11398 42194 11450
rect 42206 11398 42258 11450
rect 46950 11398 47002 11450
rect 47014 11398 47066 11450
rect 47078 11398 47130 11450
rect 47142 11398 47194 11450
rect 47206 11398 47258 11450
rect 51950 11398 52002 11450
rect 52014 11398 52066 11450
rect 52078 11398 52130 11450
rect 52142 11398 52194 11450
rect 52206 11398 52258 11450
rect 56950 11398 57002 11450
rect 57014 11398 57066 11450
rect 57078 11398 57130 11450
rect 57142 11398 57194 11450
rect 57206 11398 57258 11450
rect 58532 11135 58584 11144
rect 58532 11101 58541 11135
rect 58541 11101 58575 11135
rect 58575 11101 58584 11135
rect 58532 11092 58584 11101
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 22610 10854 22662 10906
rect 22674 10854 22726 10906
rect 22738 10854 22790 10906
rect 22802 10854 22854 10906
rect 22866 10854 22918 10906
rect 27610 10854 27662 10906
rect 27674 10854 27726 10906
rect 27738 10854 27790 10906
rect 27802 10854 27854 10906
rect 27866 10854 27918 10906
rect 32610 10854 32662 10906
rect 32674 10854 32726 10906
rect 32738 10854 32790 10906
rect 32802 10854 32854 10906
rect 32866 10854 32918 10906
rect 37610 10854 37662 10906
rect 37674 10854 37726 10906
rect 37738 10854 37790 10906
rect 37802 10854 37854 10906
rect 37866 10854 37918 10906
rect 42610 10854 42662 10906
rect 42674 10854 42726 10906
rect 42738 10854 42790 10906
rect 42802 10854 42854 10906
rect 42866 10854 42918 10906
rect 47610 10854 47662 10906
rect 47674 10854 47726 10906
rect 47738 10854 47790 10906
rect 47802 10854 47854 10906
rect 47866 10854 47918 10906
rect 52610 10854 52662 10906
rect 52674 10854 52726 10906
rect 52738 10854 52790 10906
rect 52802 10854 52854 10906
rect 52866 10854 52918 10906
rect 57610 10854 57662 10906
rect 57674 10854 57726 10906
rect 57738 10854 57790 10906
rect 57802 10854 57854 10906
rect 57866 10854 57918 10906
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 21950 10310 22002 10362
rect 22014 10310 22066 10362
rect 22078 10310 22130 10362
rect 22142 10310 22194 10362
rect 22206 10310 22258 10362
rect 26950 10310 27002 10362
rect 27014 10310 27066 10362
rect 27078 10310 27130 10362
rect 27142 10310 27194 10362
rect 27206 10310 27258 10362
rect 31950 10310 32002 10362
rect 32014 10310 32066 10362
rect 32078 10310 32130 10362
rect 32142 10310 32194 10362
rect 32206 10310 32258 10362
rect 36950 10310 37002 10362
rect 37014 10310 37066 10362
rect 37078 10310 37130 10362
rect 37142 10310 37194 10362
rect 37206 10310 37258 10362
rect 41950 10310 42002 10362
rect 42014 10310 42066 10362
rect 42078 10310 42130 10362
rect 42142 10310 42194 10362
rect 42206 10310 42258 10362
rect 46950 10310 47002 10362
rect 47014 10310 47066 10362
rect 47078 10310 47130 10362
rect 47142 10310 47194 10362
rect 47206 10310 47258 10362
rect 51950 10310 52002 10362
rect 52014 10310 52066 10362
rect 52078 10310 52130 10362
rect 52142 10310 52194 10362
rect 52206 10310 52258 10362
rect 56950 10310 57002 10362
rect 57014 10310 57066 10362
rect 57078 10310 57130 10362
rect 57142 10310 57194 10362
rect 57206 10310 57258 10362
rect 58532 10047 58584 10056
rect 58532 10013 58541 10047
rect 58541 10013 58575 10047
rect 58575 10013 58584 10047
rect 58532 10004 58584 10013
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 22610 9766 22662 9818
rect 22674 9766 22726 9818
rect 22738 9766 22790 9818
rect 22802 9766 22854 9818
rect 22866 9766 22918 9818
rect 27610 9766 27662 9818
rect 27674 9766 27726 9818
rect 27738 9766 27790 9818
rect 27802 9766 27854 9818
rect 27866 9766 27918 9818
rect 32610 9766 32662 9818
rect 32674 9766 32726 9818
rect 32738 9766 32790 9818
rect 32802 9766 32854 9818
rect 32866 9766 32918 9818
rect 37610 9766 37662 9818
rect 37674 9766 37726 9818
rect 37738 9766 37790 9818
rect 37802 9766 37854 9818
rect 37866 9766 37918 9818
rect 42610 9766 42662 9818
rect 42674 9766 42726 9818
rect 42738 9766 42790 9818
rect 42802 9766 42854 9818
rect 42866 9766 42918 9818
rect 47610 9766 47662 9818
rect 47674 9766 47726 9818
rect 47738 9766 47790 9818
rect 47802 9766 47854 9818
rect 47866 9766 47918 9818
rect 52610 9766 52662 9818
rect 52674 9766 52726 9818
rect 52738 9766 52790 9818
rect 52802 9766 52854 9818
rect 52866 9766 52918 9818
rect 57610 9766 57662 9818
rect 57674 9766 57726 9818
rect 57738 9766 57790 9818
rect 57802 9766 57854 9818
rect 57866 9766 57918 9818
rect 58532 9367 58584 9376
rect 58532 9333 58541 9367
rect 58541 9333 58575 9367
rect 58575 9333 58584 9367
rect 58532 9324 58584 9333
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 21950 9222 22002 9274
rect 22014 9222 22066 9274
rect 22078 9222 22130 9274
rect 22142 9222 22194 9274
rect 22206 9222 22258 9274
rect 26950 9222 27002 9274
rect 27014 9222 27066 9274
rect 27078 9222 27130 9274
rect 27142 9222 27194 9274
rect 27206 9222 27258 9274
rect 31950 9222 32002 9274
rect 32014 9222 32066 9274
rect 32078 9222 32130 9274
rect 32142 9222 32194 9274
rect 32206 9222 32258 9274
rect 36950 9222 37002 9274
rect 37014 9222 37066 9274
rect 37078 9222 37130 9274
rect 37142 9222 37194 9274
rect 37206 9222 37258 9274
rect 41950 9222 42002 9274
rect 42014 9222 42066 9274
rect 42078 9222 42130 9274
rect 42142 9222 42194 9274
rect 42206 9222 42258 9274
rect 46950 9222 47002 9274
rect 47014 9222 47066 9274
rect 47078 9222 47130 9274
rect 47142 9222 47194 9274
rect 47206 9222 47258 9274
rect 51950 9222 52002 9274
rect 52014 9222 52066 9274
rect 52078 9222 52130 9274
rect 52142 9222 52194 9274
rect 52206 9222 52258 9274
rect 56950 9222 57002 9274
rect 57014 9222 57066 9274
rect 57078 9222 57130 9274
rect 57142 9222 57194 9274
rect 57206 9222 57258 9274
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 22610 8678 22662 8730
rect 22674 8678 22726 8730
rect 22738 8678 22790 8730
rect 22802 8678 22854 8730
rect 22866 8678 22918 8730
rect 27610 8678 27662 8730
rect 27674 8678 27726 8730
rect 27738 8678 27790 8730
rect 27802 8678 27854 8730
rect 27866 8678 27918 8730
rect 32610 8678 32662 8730
rect 32674 8678 32726 8730
rect 32738 8678 32790 8730
rect 32802 8678 32854 8730
rect 32866 8678 32918 8730
rect 37610 8678 37662 8730
rect 37674 8678 37726 8730
rect 37738 8678 37790 8730
rect 37802 8678 37854 8730
rect 37866 8678 37918 8730
rect 42610 8678 42662 8730
rect 42674 8678 42726 8730
rect 42738 8678 42790 8730
rect 42802 8678 42854 8730
rect 42866 8678 42918 8730
rect 47610 8678 47662 8730
rect 47674 8678 47726 8730
rect 47738 8678 47790 8730
rect 47802 8678 47854 8730
rect 47866 8678 47918 8730
rect 52610 8678 52662 8730
rect 52674 8678 52726 8730
rect 52738 8678 52790 8730
rect 52802 8678 52854 8730
rect 52866 8678 52918 8730
rect 57610 8678 57662 8730
rect 57674 8678 57726 8730
rect 57738 8678 57790 8730
rect 57802 8678 57854 8730
rect 57866 8678 57918 8730
rect 58532 8347 58584 8356
rect 58532 8313 58541 8347
rect 58541 8313 58575 8347
rect 58575 8313 58584 8347
rect 58532 8304 58584 8313
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 21950 8134 22002 8186
rect 22014 8134 22066 8186
rect 22078 8134 22130 8186
rect 22142 8134 22194 8186
rect 22206 8134 22258 8186
rect 26950 8134 27002 8186
rect 27014 8134 27066 8186
rect 27078 8134 27130 8186
rect 27142 8134 27194 8186
rect 27206 8134 27258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 36950 8134 37002 8186
rect 37014 8134 37066 8186
rect 37078 8134 37130 8186
rect 37142 8134 37194 8186
rect 37206 8134 37258 8186
rect 41950 8134 42002 8186
rect 42014 8134 42066 8186
rect 42078 8134 42130 8186
rect 42142 8134 42194 8186
rect 42206 8134 42258 8186
rect 46950 8134 47002 8186
rect 47014 8134 47066 8186
rect 47078 8134 47130 8186
rect 47142 8134 47194 8186
rect 47206 8134 47258 8186
rect 51950 8134 52002 8186
rect 52014 8134 52066 8186
rect 52078 8134 52130 8186
rect 52142 8134 52194 8186
rect 52206 8134 52258 8186
rect 56950 8134 57002 8186
rect 57014 8134 57066 8186
rect 57078 8134 57130 8186
rect 57142 8134 57194 8186
rect 57206 8134 57258 8186
rect 58532 7871 58584 7880
rect 58532 7837 58541 7871
rect 58541 7837 58575 7871
rect 58575 7837 58584 7871
rect 58532 7828 58584 7837
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 22610 7590 22662 7642
rect 22674 7590 22726 7642
rect 22738 7590 22790 7642
rect 22802 7590 22854 7642
rect 22866 7590 22918 7642
rect 27610 7590 27662 7642
rect 27674 7590 27726 7642
rect 27738 7590 27790 7642
rect 27802 7590 27854 7642
rect 27866 7590 27918 7642
rect 32610 7590 32662 7642
rect 32674 7590 32726 7642
rect 32738 7590 32790 7642
rect 32802 7590 32854 7642
rect 32866 7590 32918 7642
rect 37610 7590 37662 7642
rect 37674 7590 37726 7642
rect 37738 7590 37790 7642
rect 37802 7590 37854 7642
rect 37866 7590 37918 7642
rect 42610 7590 42662 7642
rect 42674 7590 42726 7642
rect 42738 7590 42790 7642
rect 42802 7590 42854 7642
rect 42866 7590 42918 7642
rect 47610 7590 47662 7642
rect 47674 7590 47726 7642
rect 47738 7590 47790 7642
rect 47802 7590 47854 7642
rect 47866 7590 47918 7642
rect 52610 7590 52662 7642
rect 52674 7590 52726 7642
rect 52738 7590 52790 7642
rect 52802 7590 52854 7642
rect 52866 7590 52918 7642
rect 57610 7590 57662 7642
rect 57674 7590 57726 7642
rect 57738 7590 57790 7642
rect 57802 7590 57854 7642
rect 57866 7590 57918 7642
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 21950 7046 22002 7098
rect 22014 7046 22066 7098
rect 22078 7046 22130 7098
rect 22142 7046 22194 7098
rect 22206 7046 22258 7098
rect 26950 7046 27002 7098
rect 27014 7046 27066 7098
rect 27078 7046 27130 7098
rect 27142 7046 27194 7098
rect 27206 7046 27258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 36950 7046 37002 7098
rect 37014 7046 37066 7098
rect 37078 7046 37130 7098
rect 37142 7046 37194 7098
rect 37206 7046 37258 7098
rect 41950 7046 42002 7098
rect 42014 7046 42066 7098
rect 42078 7046 42130 7098
rect 42142 7046 42194 7098
rect 42206 7046 42258 7098
rect 46950 7046 47002 7098
rect 47014 7046 47066 7098
rect 47078 7046 47130 7098
rect 47142 7046 47194 7098
rect 47206 7046 47258 7098
rect 51950 7046 52002 7098
rect 52014 7046 52066 7098
rect 52078 7046 52130 7098
rect 52142 7046 52194 7098
rect 52206 7046 52258 7098
rect 56950 7046 57002 7098
rect 57014 7046 57066 7098
rect 57078 7046 57130 7098
rect 57142 7046 57194 7098
rect 57206 7046 57258 7098
rect 58532 6783 58584 6792
rect 58532 6749 58541 6783
rect 58541 6749 58575 6783
rect 58575 6749 58584 6783
rect 58532 6740 58584 6749
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 22610 6502 22662 6554
rect 22674 6502 22726 6554
rect 22738 6502 22790 6554
rect 22802 6502 22854 6554
rect 22866 6502 22918 6554
rect 27610 6502 27662 6554
rect 27674 6502 27726 6554
rect 27738 6502 27790 6554
rect 27802 6502 27854 6554
rect 27866 6502 27918 6554
rect 32610 6502 32662 6554
rect 32674 6502 32726 6554
rect 32738 6502 32790 6554
rect 32802 6502 32854 6554
rect 32866 6502 32918 6554
rect 37610 6502 37662 6554
rect 37674 6502 37726 6554
rect 37738 6502 37790 6554
rect 37802 6502 37854 6554
rect 37866 6502 37918 6554
rect 42610 6502 42662 6554
rect 42674 6502 42726 6554
rect 42738 6502 42790 6554
rect 42802 6502 42854 6554
rect 42866 6502 42918 6554
rect 47610 6502 47662 6554
rect 47674 6502 47726 6554
rect 47738 6502 47790 6554
rect 47802 6502 47854 6554
rect 47866 6502 47918 6554
rect 52610 6502 52662 6554
rect 52674 6502 52726 6554
rect 52738 6502 52790 6554
rect 52802 6502 52854 6554
rect 52866 6502 52918 6554
rect 57610 6502 57662 6554
rect 57674 6502 57726 6554
rect 57738 6502 57790 6554
rect 57802 6502 57854 6554
rect 57866 6502 57918 6554
rect 58532 6103 58584 6112
rect 58532 6069 58541 6103
rect 58541 6069 58575 6103
rect 58575 6069 58584 6103
rect 58532 6060 58584 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 21950 5958 22002 6010
rect 22014 5958 22066 6010
rect 22078 5958 22130 6010
rect 22142 5958 22194 6010
rect 22206 5958 22258 6010
rect 26950 5958 27002 6010
rect 27014 5958 27066 6010
rect 27078 5958 27130 6010
rect 27142 5958 27194 6010
rect 27206 5958 27258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 36950 5958 37002 6010
rect 37014 5958 37066 6010
rect 37078 5958 37130 6010
rect 37142 5958 37194 6010
rect 37206 5958 37258 6010
rect 41950 5958 42002 6010
rect 42014 5958 42066 6010
rect 42078 5958 42130 6010
rect 42142 5958 42194 6010
rect 42206 5958 42258 6010
rect 46950 5958 47002 6010
rect 47014 5958 47066 6010
rect 47078 5958 47130 6010
rect 47142 5958 47194 6010
rect 47206 5958 47258 6010
rect 51950 5958 52002 6010
rect 52014 5958 52066 6010
rect 52078 5958 52130 6010
rect 52142 5958 52194 6010
rect 52206 5958 52258 6010
rect 56950 5958 57002 6010
rect 57014 5958 57066 6010
rect 57078 5958 57130 6010
rect 57142 5958 57194 6010
rect 57206 5958 57258 6010
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 22610 5414 22662 5466
rect 22674 5414 22726 5466
rect 22738 5414 22790 5466
rect 22802 5414 22854 5466
rect 22866 5414 22918 5466
rect 27610 5414 27662 5466
rect 27674 5414 27726 5466
rect 27738 5414 27790 5466
rect 27802 5414 27854 5466
rect 27866 5414 27918 5466
rect 32610 5414 32662 5466
rect 32674 5414 32726 5466
rect 32738 5414 32790 5466
rect 32802 5414 32854 5466
rect 32866 5414 32918 5466
rect 37610 5414 37662 5466
rect 37674 5414 37726 5466
rect 37738 5414 37790 5466
rect 37802 5414 37854 5466
rect 37866 5414 37918 5466
rect 42610 5414 42662 5466
rect 42674 5414 42726 5466
rect 42738 5414 42790 5466
rect 42802 5414 42854 5466
rect 42866 5414 42918 5466
rect 47610 5414 47662 5466
rect 47674 5414 47726 5466
rect 47738 5414 47790 5466
rect 47802 5414 47854 5466
rect 47866 5414 47918 5466
rect 52610 5414 52662 5466
rect 52674 5414 52726 5466
rect 52738 5414 52790 5466
rect 52802 5414 52854 5466
rect 52866 5414 52918 5466
rect 57610 5414 57662 5466
rect 57674 5414 57726 5466
rect 57738 5414 57790 5466
rect 57802 5414 57854 5466
rect 57866 5414 57918 5466
rect 58532 5015 58584 5024
rect 58532 4981 58541 5015
rect 58541 4981 58575 5015
rect 58575 4981 58584 5015
rect 58532 4972 58584 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 21950 4870 22002 4922
rect 22014 4870 22066 4922
rect 22078 4870 22130 4922
rect 22142 4870 22194 4922
rect 22206 4870 22258 4922
rect 26950 4870 27002 4922
rect 27014 4870 27066 4922
rect 27078 4870 27130 4922
rect 27142 4870 27194 4922
rect 27206 4870 27258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 36950 4870 37002 4922
rect 37014 4870 37066 4922
rect 37078 4870 37130 4922
rect 37142 4870 37194 4922
rect 37206 4870 37258 4922
rect 41950 4870 42002 4922
rect 42014 4870 42066 4922
rect 42078 4870 42130 4922
rect 42142 4870 42194 4922
rect 42206 4870 42258 4922
rect 46950 4870 47002 4922
rect 47014 4870 47066 4922
rect 47078 4870 47130 4922
rect 47142 4870 47194 4922
rect 47206 4870 47258 4922
rect 51950 4870 52002 4922
rect 52014 4870 52066 4922
rect 52078 4870 52130 4922
rect 52142 4870 52194 4922
rect 52206 4870 52258 4922
rect 56950 4870 57002 4922
rect 57014 4870 57066 4922
rect 57078 4870 57130 4922
rect 57142 4870 57194 4922
rect 57206 4870 57258 4922
rect 58532 4607 58584 4616
rect 58532 4573 58541 4607
rect 58541 4573 58575 4607
rect 58575 4573 58584 4607
rect 58532 4564 58584 4573
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 22610 4326 22662 4378
rect 22674 4326 22726 4378
rect 22738 4326 22790 4378
rect 22802 4326 22854 4378
rect 22866 4326 22918 4378
rect 27610 4326 27662 4378
rect 27674 4326 27726 4378
rect 27738 4326 27790 4378
rect 27802 4326 27854 4378
rect 27866 4326 27918 4378
rect 32610 4326 32662 4378
rect 32674 4326 32726 4378
rect 32738 4326 32790 4378
rect 32802 4326 32854 4378
rect 32866 4326 32918 4378
rect 37610 4326 37662 4378
rect 37674 4326 37726 4378
rect 37738 4326 37790 4378
rect 37802 4326 37854 4378
rect 37866 4326 37918 4378
rect 42610 4326 42662 4378
rect 42674 4326 42726 4378
rect 42738 4326 42790 4378
rect 42802 4326 42854 4378
rect 42866 4326 42918 4378
rect 47610 4326 47662 4378
rect 47674 4326 47726 4378
rect 47738 4326 47790 4378
rect 47802 4326 47854 4378
rect 47866 4326 47918 4378
rect 52610 4326 52662 4378
rect 52674 4326 52726 4378
rect 52738 4326 52790 4378
rect 52802 4326 52854 4378
rect 52866 4326 52918 4378
rect 57610 4326 57662 4378
rect 57674 4326 57726 4378
rect 57738 4326 57790 4378
rect 57802 4326 57854 4378
rect 57866 4326 57918 4378
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 21950 3782 22002 3834
rect 22014 3782 22066 3834
rect 22078 3782 22130 3834
rect 22142 3782 22194 3834
rect 22206 3782 22258 3834
rect 26950 3782 27002 3834
rect 27014 3782 27066 3834
rect 27078 3782 27130 3834
rect 27142 3782 27194 3834
rect 27206 3782 27258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 36950 3782 37002 3834
rect 37014 3782 37066 3834
rect 37078 3782 37130 3834
rect 37142 3782 37194 3834
rect 37206 3782 37258 3834
rect 41950 3782 42002 3834
rect 42014 3782 42066 3834
rect 42078 3782 42130 3834
rect 42142 3782 42194 3834
rect 42206 3782 42258 3834
rect 46950 3782 47002 3834
rect 47014 3782 47066 3834
rect 47078 3782 47130 3834
rect 47142 3782 47194 3834
rect 47206 3782 47258 3834
rect 51950 3782 52002 3834
rect 52014 3782 52066 3834
rect 52078 3782 52130 3834
rect 52142 3782 52194 3834
rect 52206 3782 52258 3834
rect 56950 3782 57002 3834
rect 57014 3782 57066 3834
rect 57078 3782 57130 3834
rect 57142 3782 57194 3834
rect 57206 3782 57258 3834
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 22610 3238 22662 3290
rect 22674 3238 22726 3290
rect 22738 3238 22790 3290
rect 22802 3238 22854 3290
rect 22866 3238 22918 3290
rect 27610 3238 27662 3290
rect 27674 3238 27726 3290
rect 27738 3238 27790 3290
rect 27802 3238 27854 3290
rect 27866 3238 27918 3290
rect 32610 3238 32662 3290
rect 32674 3238 32726 3290
rect 32738 3238 32790 3290
rect 32802 3238 32854 3290
rect 32866 3238 32918 3290
rect 37610 3238 37662 3290
rect 37674 3238 37726 3290
rect 37738 3238 37790 3290
rect 37802 3238 37854 3290
rect 37866 3238 37918 3290
rect 42610 3238 42662 3290
rect 42674 3238 42726 3290
rect 42738 3238 42790 3290
rect 42802 3238 42854 3290
rect 42866 3238 42918 3290
rect 47610 3238 47662 3290
rect 47674 3238 47726 3290
rect 47738 3238 47790 3290
rect 47802 3238 47854 3290
rect 47866 3238 47918 3290
rect 52610 3238 52662 3290
rect 52674 3238 52726 3290
rect 52738 3238 52790 3290
rect 52802 3238 52854 3290
rect 52866 3238 52918 3290
rect 57610 3238 57662 3290
rect 57674 3238 57726 3290
rect 57738 3238 57790 3290
rect 57802 3238 57854 3290
rect 57866 3238 57918 3290
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 21950 2694 22002 2746
rect 22014 2694 22066 2746
rect 22078 2694 22130 2746
rect 22142 2694 22194 2746
rect 22206 2694 22258 2746
rect 26950 2694 27002 2746
rect 27014 2694 27066 2746
rect 27078 2694 27130 2746
rect 27142 2694 27194 2746
rect 27206 2694 27258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 36950 2694 37002 2746
rect 37014 2694 37066 2746
rect 37078 2694 37130 2746
rect 37142 2694 37194 2746
rect 37206 2694 37258 2746
rect 41950 2694 42002 2746
rect 42014 2694 42066 2746
rect 42078 2694 42130 2746
rect 42142 2694 42194 2746
rect 42206 2694 42258 2746
rect 46950 2694 47002 2746
rect 47014 2694 47066 2746
rect 47078 2694 47130 2746
rect 47142 2694 47194 2746
rect 47206 2694 47258 2746
rect 51950 2694 52002 2746
rect 52014 2694 52066 2746
rect 52078 2694 52130 2746
rect 52142 2694 52194 2746
rect 52206 2694 52258 2746
rect 56950 2694 57002 2746
rect 57014 2694 57066 2746
rect 57078 2694 57130 2746
rect 57142 2694 57194 2746
rect 57206 2694 57258 2746
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
rect 22610 2150 22662 2202
rect 22674 2150 22726 2202
rect 22738 2150 22790 2202
rect 22802 2150 22854 2202
rect 22866 2150 22918 2202
rect 27610 2150 27662 2202
rect 27674 2150 27726 2202
rect 27738 2150 27790 2202
rect 27802 2150 27854 2202
rect 27866 2150 27918 2202
rect 32610 2150 32662 2202
rect 32674 2150 32726 2202
rect 32738 2150 32790 2202
rect 32802 2150 32854 2202
rect 32866 2150 32918 2202
rect 37610 2150 37662 2202
rect 37674 2150 37726 2202
rect 37738 2150 37790 2202
rect 37802 2150 37854 2202
rect 37866 2150 37918 2202
rect 42610 2150 42662 2202
rect 42674 2150 42726 2202
rect 42738 2150 42790 2202
rect 42802 2150 42854 2202
rect 42866 2150 42918 2202
rect 47610 2150 47662 2202
rect 47674 2150 47726 2202
rect 47738 2150 47790 2202
rect 47802 2150 47854 2202
rect 47866 2150 47918 2202
rect 52610 2150 52662 2202
rect 52674 2150 52726 2202
rect 52738 2150 52790 2202
rect 52802 2150 52854 2202
rect 52866 2150 52918 2202
rect 57610 2150 57662 2202
rect 57674 2150 57726 2202
rect 57738 2150 57790 2202
rect 57802 2150 57854 2202
rect 57866 2150 57918 2202
<< metal2 >>
rect 2610 57692 2918 57701
rect 2610 57690 2616 57692
rect 2672 57690 2696 57692
rect 2752 57690 2776 57692
rect 2832 57690 2856 57692
rect 2912 57690 2918 57692
rect 2672 57638 2674 57690
rect 2854 57638 2856 57690
rect 2610 57636 2616 57638
rect 2672 57636 2696 57638
rect 2752 57636 2776 57638
rect 2832 57636 2856 57638
rect 2912 57636 2918 57638
rect 2610 57627 2918 57636
rect 7610 57692 7918 57701
rect 7610 57690 7616 57692
rect 7672 57690 7696 57692
rect 7752 57690 7776 57692
rect 7832 57690 7856 57692
rect 7912 57690 7918 57692
rect 7672 57638 7674 57690
rect 7854 57638 7856 57690
rect 7610 57636 7616 57638
rect 7672 57636 7696 57638
rect 7752 57636 7776 57638
rect 7832 57636 7856 57638
rect 7912 57636 7918 57638
rect 7610 57627 7918 57636
rect 12610 57692 12918 57701
rect 12610 57690 12616 57692
rect 12672 57690 12696 57692
rect 12752 57690 12776 57692
rect 12832 57690 12856 57692
rect 12912 57690 12918 57692
rect 12672 57638 12674 57690
rect 12854 57638 12856 57690
rect 12610 57636 12616 57638
rect 12672 57636 12696 57638
rect 12752 57636 12776 57638
rect 12832 57636 12856 57638
rect 12912 57636 12918 57638
rect 12610 57627 12918 57636
rect 17610 57692 17918 57701
rect 17610 57690 17616 57692
rect 17672 57690 17696 57692
rect 17752 57690 17776 57692
rect 17832 57690 17856 57692
rect 17912 57690 17918 57692
rect 17672 57638 17674 57690
rect 17854 57638 17856 57690
rect 17610 57636 17616 57638
rect 17672 57636 17696 57638
rect 17752 57636 17776 57638
rect 17832 57636 17856 57638
rect 17912 57636 17918 57638
rect 17610 57627 17918 57636
rect 22610 57692 22918 57701
rect 22610 57690 22616 57692
rect 22672 57690 22696 57692
rect 22752 57690 22776 57692
rect 22832 57690 22856 57692
rect 22912 57690 22918 57692
rect 22672 57638 22674 57690
rect 22854 57638 22856 57690
rect 22610 57636 22616 57638
rect 22672 57636 22696 57638
rect 22752 57636 22776 57638
rect 22832 57636 22856 57638
rect 22912 57636 22918 57638
rect 22610 57627 22918 57636
rect 27610 57692 27918 57701
rect 27610 57690 27616 57692
rect 27672 57690 27696 57692
rect 27752 57690 27776 57692
rect 27832 57690 27856 57692
rect 27912 57690 27918 57692
rect 27672 57638 27674 57690
rect 27854 57638 27856 57690
rect 27610 57636 27616 57638
rect 27672 57636 27696 57638
rect 27752 57636 27776 57638
rect 27832 57636 27856 57638
rect 27912 57636 27918 57638
rect 27610 57627 27918 57636
rect 32610 57692 32918 57701
rect 32610 57690 32616 57692
rect 32672 57690 32696 57692
rect 32752 57690 32776 57692
rect 32832 57690 32856 57692
rect 32912 57690 32918 57692
rect 32672 57638 32674 57690
rect 32854 57638 32856 57690
rect 32610 57636 32616 57638
rect 32672 57636 32696 57638
rect 32752 57636 32776 57638
rect 32832 57636 32856 57638
rect 32912 57636 32918 57638
rect 32610 57627 32918 57636
rect 37610 57692 37918 57701
rect 37610 57690 37616 57692
rect 37672 57690 37696 57692
rect 37752 57690 37776 57692
rect 37832 57690 37856 57692
rect 37912 57690 37918 57692
rect 37672 57638 37674 57690
rect 37854 57638 37856 57690
rect 37610 57636 37616 57638
rect 37672 57636 37696 57638
rect 37752 57636 37776 57638
rect 37832 57636 37856 57638
rect 37912 57636 37918 57638
rect 37610 57627 37918 57636
rect 42610 57692 42918 57701
rect 42610 57690 42616 57692
rect 42672 57690 42696 57692
rect 42752 57690 42776 57692
rect 42832 57690 42856 57692
rect 42912 57690 42918 57692
rect 42672 57638 42674 57690
rect 42854 57638 42856 57690
rect 42610 57636 42616 57638
rect 42672 57636 42696 57638
rect 42752 57636 42776 57638
rect 42832 57636 42856 57638
rect 42912 57636 42918 57638
rect 42610 57627 42918 57636
rect 47610 57692 47918 57701
rect 47610 57690 47616 57692
rect 47672 57690 47696 57692
rect 47752 57690 47776 57692
rect 47832 57690 47856 57692
rect 47912 57690 47918 57692
rect 47672 57638 47674 57690
rect 47854 57638 47856 57690
rect 47610 57636 47616 57638
rect 47672 57636 47696 57638
rect 47752 57636 47776 57638
rect 47832 57636 47856 57638
rect 47912 57636 47918 57638
rect 47610 57627 47918 57636
rect 52610 57692 52918 57701
rect 52610 57690 52616 57692
rect 52672 57690 52696 57692
rect 52752 57690 52776 57692
rect 52832 57690 52856 57692
rect 52912 57690 52918 57692
rect 52672 57638 52674 57690
rect 52854 57638 52856 57690
rect 52610 57636 52616 57638
rect 52672 57636 52696 57638
rect 52752 57636 52776 57638
rect 52832 57636 52856 57638
rect 52912 57636 52918 57638
rect 52610 57627 52918 57636
rect 57610 57692 57918 57701
rect 57610 57690 57616 57692
rect 57672 57690 57696 57692
rect 57752 57690 57776 57692
rect 57832 57690 57856 57692
rect 57912 57690 57918 57692
rect 57672 57638 57674 57690
rect 57854 57638 57856 57690
rect 57610 57636 57616 57638
rect 57672 57636 57696 57638
rect 57752 57636 57776 57638
rect 57832 57636 57856 57638
rect 57912 57636 57918 57638
rect 57610 57627 57918 57636
rect 1950 57148 2258 57157
rect 1950 57146 1956 57148
rect 2012 57146 2036 57148
rect 2092 57146 2116 57148
rect 2172 57146 2196 57148
rect 2252 57146 2258 57148
rect 2012 57094 2014 57146
rect 2194 57094 2196 57146
rect 1950 57092 1956 57094
rect 2012 57092 2036 57094
rect 2092 57092 2116 57094
rect 2172 57092 2196 57094
rect 2252 57092 2258 57094
rect 1950 57083 2258 57092
rect 6950 57148 7258 57157
rect 6950 57146 6956 57148
rect 7012 57146 7036 57148
rect 7092 57146 7116 57148
rect 7172 57146 7196 57148
rect 7252 57146 7258 57148
rect 7012 57094 7014 57146
rect 7194 57094 7196 57146
rect 6950 57092 6956 57094
rect 7012 57092 7036 57094
rect 7092 57092 7116 57094
rect 7172 57092 7196 57094
rect 7252 57092 7258 57094
rect 6950 57083 7258 57092
rect 11950 57148 12258 57157
rect 11950 57146 11956 57148
rect 12012 57146 12036 57148
rect 12092 57146 12116 57148
rect 12172 57146 12196 57148
rect 12252 57146 12258 57148
rect 12012 57094 12014 57146
rect 12194 57094 12196 57146
rect 11950 57092 11956 57094
rect 12012 57092 12036 57094
rect 12092 57092 12116 57094
rect 12172 57092 12196 57094
rect 12252 57092 12258 57094
rect 11950 57083 12258 57092
rect 16950 57148 17258 57157
rect 16950 57146 16956 57148
rect 17012 57146 17036 57148
rect 17092 57146 17116 57148
rect 17172 57146 17196 57148
rect 17252 57146 17258 57148
rect 17012 57094 17014 57146
rect 17194 57094 17196 57146
rect 16950 57092 16956 57094
rect 17012 57092 17036 57094
rect 17092 57092 17116 57094
rect 17172 57092 17196 57094
rect 17252 57092 17258 57094
rect 16950 57083 17258 57092
rect 21950 57148 22258 57157
rect 21950 57146 21956 57148
rect 22012 57146 22036 57148
rect 22092 57146 22116 57148
rect 22172 57146 22196 57148
rect 22252 57146 22258 57148
rect 22012 57094 22014 57146
rect 22194 57094 22196 57146
rect 21950 57092 21956 57094
rect 22012 57092 22036 57094
rect 22092 57092 22116 57094
rect 22172 57092 22196 57094
rect 22252 57092 22258 57094
rect 21950 57083 22258 57092
rect 26950 57148 27258 57157
rect 26950 57146 26956 57148
rect 27012 57146 27036 57148
rect 27092 57146 27116 57148
rect 27172 57146 27196 57148
rect 27252 57146 27258 57148
rect 27012 57094 27014 57146
rect 27194 57094 27196 57146
rect 26950 57092 26956 57094
rect 27012 57092 27036 57094
rect 27092 57092 27116 57094
rect 27172 57092 27196 57094
rect 27252 57092 27258 57094
rect 26950 57083 27258 57092
rect 31950 57148 32258 57157
rect 31950 57146 31956 57148
rect 32012 57146 32036 57148
rect 32092 57146 32116 57148
rect 32172 57146 32196 57148
rect 32252 57146 32258 57148
rect 32012 57094 32014 57146
rect 32194 57094 32196 57146
rect 31950 57092 31956 57094
rect 32012 57092 32036 57094
rect 32092 57092 32116 57094
rect 32172 57092 32196 57094
rect 32252 57092 32258 57094
rect 31950 57083 32258 57092
rect 36950 57148 37258 57157
rect 36950 57146 36956 57148
rect 37012 57146 37036 57148
rect 37092 57146 37116 57148
rect 37172 57146 37196 57148
rect 37252 57146 37258 57148
rect 37012 57094 37014 57146
rect 37194 57094 37196 57146
rect 36950 57092 36956 57094
rect 37012 57092 37036 57094
rect 37092 57092 37116 57094
rect 37172 57092 37196 57094
rect 37252 57092 37258 57094
rect 36950 57083 37258 57092
rect 41950 57148 42258 57157
rect 41950 57146 41956 57148
rect 42012 57146 42036 57148
rect 42092 57146 42116 57148
rect 42172 57146 42196 57148
rect 42252 57146 42258 57148
rect 42012 57094 42014 57146
rect 42194 57094 42196 57146
rect 41950 57092 41956 57094
rect 42012 57092 42036 57094
rect 42092 57092 42116 57094
rect 42172 57092 42196 57094
rect 42252 57092 42258 57094
rect 41950 57083 42258 57092
rect 46950 57148 47258 57157
rect 46950 57146 46956 57148
rect 47012 57146 47036 57148
rect 47092 57146 47116 57148
rect 47172 57146 47196 57148
rect 47252 57146 47258 57148
rect 47012 57094 47014 57146
rect 47194 57094 47196 57146
rect 46950 57092 46956 57094
rect 47012 57092 47036 57094
rect 47092 57092 47116 57094
rect 47172 57092 47196 57094
rect 47252 57092 47258 57094
rect 46950 57083 47258 57092
rect 51950 57148 52258 57157
rect 51950 57146 51956 57148
rect 52012 57146 52036 57148
rect 52092 57146 52116 57148
rect 52172 57146 52196 57148
rect 52252 57146 52258 57148
rect 52012 57094 52014 57146
rect 52194 57094 52196 57146
rect 51950 57092 51956 57094
rect 52012 57092 52036 57094
rect 52092 57092 52116 57094
rect 52172 57092 52196 57094
rect 52252 57092 52258 57094
rect 51950 57083 52258 57092
rect 56950 57148 57258 57157
rect 56950 57146 56956 57148
rect 57012 57146 57036 57148
rect 57092 57146 57116 57148
rect 57172 57146 57196 57148
rect 57252 57146 57258 57148
rect 57012 57094 57014 57146
rect 57194 57094 57196 57146
rect 56950 57092 56956 57094
rect 57012 57092 57036 57094
rect 57092 57092 57116 57094
rect 57172 57092 57196 57094
rect 57252 57092 57258 57094
rect 56950 57083 57258 57092
rect 2610 56604 2918 56613
rect 2610 56602 2616 56604
rect 2672 56602 2696 56604
rect 2752 56602 2776 56604
rect 2832 56602 2856 56604
rect 2912 56602 2918 56604
rect 2672 56550 2674 56602
rect 2854 56550 2856 56602
rect 2610 56548 2616 56550
rect 2672 56548 2696 56550
rect 2752 56548 2776 56550
rect 2832 56548 2856 56550
rect 2912 56548 2918 56550
rect 2610 56539 2918 56548
rect 7610 56604 7918 56613
rect 7610 56602 7616 56604
rect 7672 56602 7696 56604
rect 7752 56602 7776 56604
rect 7832 56602 7856 56604
rect 7912 56602 7918 56604
rect 7672 56550 7674 56602
rect 7854 56550 7856 56602
rect 7610 56548 7616 56550
rect 7672 56548 7696 56550
rect 7752 56548 7776 56550
rect 7832 56548 7856 56550
rect 7912 56548 7918 56550
rect 7610 56539 7918 56548
rect 12610 56604 12918 56613
rect 12610 56602 12616 56604
rect 12672 56602 12696 56604
rect 12752 56602 12776 56604
rect 12832 56602 12856 56604
rect 12912 56602 12918 56604
rect 12672 56550 12674 56602
rect 12854 56550 12856 56602
rect 12610 56548 12616 56550
rect 12672 56548 12696 56550
rect 12752 56548 12776 56550
rect 12832 56548 12856 56550
rect 12912 56548 12918 56550
rect 12610 56539 12918 56548
rect 17610 56604 17918 56613
rect 17610 56602 17616 56604
rect 17672 56602 17696 56604
rect 17752 56602 17776 56604
rect 17832 56602 17856 56604
rect 17912 56602 17918 56604
rect 17672 56550 17674 56602
rect 17854 56550 17856 56602
rect 17610 56548 17616 56550
rect 17672 56548 17696 56550
rect 17752 56548 17776 56550
rect 17832 56548 17856 56550
rect 17912 56548 17918 56550
rect 17610 56539 17918 56548
rect 22610 56604 22918 56613
rect 22610 56602 22616 56604
rect 22672 56602 22696 56604
rect 22752 56602 22776 56604
rect 22832 56602 22856 56604
rect 22912 56602 22918 56604
rect 22672 56550 22674 56602
rect 22854 56550 22856 56602
rect 22610 56548 22616 56550
rect 22672 56548 22696 56550
rect 22752 56548 22776 56550
rect 22832 56548 22856 56550
rect 22912 56548 22918 56550
rect 22610 56539 22918 56548
rect 27610 56604 27918 56613
rect 27610 56602 27616 56604
rect 27672 56602 27696 56604
rect 27752 56602 27776 56604
rect 27832 56602 27856 56604
rect 27912 56602 27918 56604
rect 27672 56550 27674 56602
rect 27854 56550 27856 56602
rect 27610 56548 27616 56550
rect 27672 56548 27696 56550
rect 27752 56548 27776 56550
rect 27832 56548 27856 56550
rect 27912 56548 27918 56550
rect 27610 56539 27918 56548
rect 32610 56604 32918 56613
rect 32610 56602 32616 56604
rect 32672 56602 32696 56604
rect 32752 56602 32776 56604
rect 32832 56602 32856 56604
rect 32912 56602 32918 56604
rect 32672 56550 32674 56602
rect 32854 56550 32856 56602
rect 32610 56548 32616 56550
rect 32672 56548 32696 56550
rect 32752 56548 32776 56550
rect 32832 56548 32856 56550
rect 32912 56548 32918 56550
rect 32610 56539 32918 56548
rect 37610 56604 37918 56613
rect 37610 56602 37616 56604
rect 37672 56602 37696 56604
rect 37752 56602 37776 56604
rect 37832 56602 37856 56604
rect 37912 56602 37918 56604
rect 37672 56550 37674 56602
rect 37854 56550 37856 56602
rect 37610 56548 37616 56550
rect 37672 56548 37696 56550
rect 37752 56548 37776 56550
rect 37832 56548 37856 56550
rect 37912 56548 37918 56550
rect 37610 56539 37918 56548
rect 42610 56604 42918 56613
rect 42610 56602 42616 56604
rect 42672 56602 42696 56604
rect 42752 56602 42776 56604
rect 42832 56602 42856 56604
rect 42912 56602 42918 56604
rect 42672 56550 42674 56602
rect 42854 56550 42856 56602
rect 42610 56548 42616 56550
rect 42672 56548 42696 56550
rect 42752 56548 42776 56550
rect 42832 56548 42856 56550
rect 42912 56548 42918 56550
rect 42610 56539 42918 56548
rect 47610 56604 47918 56613
rect 47610 56602 47616 56604
rect 47672 56602 47696 56604
rect 47752 56602 47776 56604
rect 47832 56602 47856 56604
rect 47912 56602 47918 56604
rect 47672 56550 47674 56602
rect 47854 56550 47856 56602
rect 47610 56548 47616 56550
rect 47672 56548 47696 56550
rect 47752 56548 47776 56550
rect 47832 56548 47856 56550
rect 47912 56548 47918 56550
rect 47610 56539 47918 56548
rect 52610 56604 52918 56613
rect 52610 56602 52616 56604
rect 52672 56602 52696 56604
rect 52752 56602 52776 56604
rect 52832 56602 52856 56604
rect 52912 56602 52918 56604
rect 52672 56550 52674 56602
rect 52854 56550 52856 56602
rect 52610 56548 52616 56550
rect 52672 56548 52696 56550
rect 52752 56548 52776 56550
rect 52832 56548 52856 56550
rect 52912 56548 52918 56550
rect 52610 56539 52918 56548
rect 57610 56604 57918 56613
rect 57610 56602 57616 56604
rect 57672 56602 57696 56604
rect 57752 56602 57776 56604
rect 57832 56602 57856 56604
rect 57912 56602 57918 56604
rect 57672 56550 57674 56602
rect 57854 56550 57856 56602
rect 57610 56548 57616 56550
rect 57672 56548 57696 56550
rect 57752 56548 57776 56550
rect 57832 56548 57856 56550
rect 57912 56548 57918 56550
rect 57610 56539 57918 56548
rect 1950 56060 2258 56069
rect 1950 56058 1956 56060
rect 2012 56058 2036 56060
rect 2092 56058 2116 56060
rect 2172 56058 2196 56060
rect 2252 56058 2258 56060
rect 2012 56006 2014 56058
rect 2194 56006 2196 56058
rect 1950 56004 1956 56006
rect 2012 56004 2036 56006
rect 2092 56004 2116 56006
rect 2172 56004 2196 56006
rect 2252 56004 2258 56006
rect 1950 55995 2258 56004
rect 6950 56060 7258 56069
rect 6950 56058 6956 56060
rect 7012 56058 7036 56060
rect 7092 56058 7116 56060
rect 7172 56058 7196 56060
rect 7252 56058 7258 56060
rect 7012 56006 7014 56058
rect 7194 56006 7196 56058
rect 6950 56004 6956 56006
rect 7012 56004 7036 56006
rect 7092 56004 7116 56006
rect 7172 56004 7196 56006
rect 7252 56004 7258 56006
rect 6950 55995 7258 56004
rect 11950 56060 12258 56069
rect 11950 56058 11956 56060
rect 12012 56058 12036 56060
rect 12092 56058 12116 56060
rect 12172 56058 12196 56060
rect 12252 56058 12258 56060
rect 12012 56006 12014 56058
rect 12194 56006 12196 56058
rect 11950 56004 11956 56006
rect 12012 56004 12036 56006
rect 12092 56004 12116 56006
rect 12172 56004 12196 56006
rect 12252 56004 12258 56006
rect 11950 55995 12258 56004
rect 16950 56060 17258 56069
rect 16950 56058 16956 56060
rect 17012 56058 17036 56060
rect 17092 56058 17116 56060
rect 17172 56058 17196 56060
rect 17252 56058 17258 56060
rect 17012 56006 17014 56058
rect 17194 56006 17196 56058
rect 16950 56004 16956 56006
rect 17012 56004 17036 56006
rect 17092 56004 17116 56006
rect 17172 56004 17196 56006
rect 17252 56004 17258 56006
rect 16950 55995 17258 56004
rect 21950 56060 22258 56069
rect 21950 56058 21956 56060
rect 22012 56058 22036 56060
rect 22092 56058 22116 56060
rect 22172 56058 22196 56060
rect 22252 56058 22258 56060
rect 22012 56006 22014 56058
rect 22194 56006 22196 56058
rect 21950 56004 21956 56006
rect 22012 56004 22036 56006
rect 22092 56004 22116 56006
rect 22172 56004 22196 56006
rect 22252 56004 22258 56006
rect 21950 55995 22258 56004
rect 26950 56060 27258 56069
rect 26950 56058 26956 56060
rect 27012 56058 27036 56060
rect 27092 56058 27116 56060
rect 27172 56058 27196 56060
rect 27252 56058 27258 56060
rect 27012 56006 27014 56058
rect 27194 56006 27196 56058
rect 26950 56004 26956 56006
rect 27012 56004 27036 56006
rect 27092 56004 27116 56006
rect 27172 56004 27196 56006
rect 27252 56004 27258 56006
rect 26950 55995 27258 56004
rect 31950 56060 32258 56069
rect 31950 56058 31956 56060
rect 32012 56058 32036 56060
rect 32092 56058 32116 56060
rect 32172 56058 32196 56060
rect 32252 56058 32258 56060
rect 32012 56006 32014 56058
rect 32194 56006 32196 56058
rect 31950 56004 31956 56006
rect 32012 56004 32036 56006
rect 32092 56004 32116 56006
rect 32172 56004 32196 56006
rect 32252 56004 32258 56006
rect 31950 55995 32258 56004
rect 36950 56060 37258 56069
rect 36950 56058 36956 56060
rect 37012 56058 37036 56060
rect 37092 56058 37116 56060
rect 37172 56058 37196 56060
rect 37252 56058 37258 56060
rect 37012 56006 37014 56058
rect 37194 56006 37196 56058
rect 36950 56004 36956 56006
rect 37012 56004 37036 56006
rect 37092 56004 37116 56006
rect 37172 56004 37196 56006
rect 37252 56004 37258 56006
rect 36950 55995 37258 56004
rect 41950 56060 42258 56069
rect 41950 56058 41956 56060
rect 42012 56058 42036 56060
rect 42092 56058 42116 56060
rect 42172 56058 42196 56060
rect 42252 56058 42258 56060
rect 42012 56006 42014 56058
rect 42194 56006 42196 56058
rect 41950 56004 41956 56006
rect 42012 56004 42036 56006
rect 42092 56004 42116 56006
rect 42172 56004 42196 56006
rect 42252 56004 42258 56006
rect 41950 55995 42258 56004
rect 46950 56060 47258 56069
rect 46950 56058 46956 56060
rect 47012 56058 47036 56060
rect 47092 56058 47116 56060
rect 47172 56058 47196 56060
rect 47252 56058 47258 56060
rect 47012 56006 47014 56058
rect 47194 56006 47196 56058
rect 46950 56004 46956 56006
rect 47012 56004 47036 56006
rect 47092 56004 47116 56006
rect 47172 56004 47196 56006
rect 47252 56004 47258 56006
rect 46950 55995 47258 56004
rect 51950 56060 52258 56069
rect 51950 56058 51956 56060
rect 52012 56058 52036 56060
rect 52092 56058 52116 56060
rect 52172 56058 52196 56060
rect 52252 56058 52258 56060
rect 52012 56006 52014 56058
rect 52194 56006 52196 56058
rect 51950 56004 51956 56006
rect 52012 56004 52036 56006
rect 52092 56004 52116 56006
rect 52172 56004 52196 56006
rect 52252 56004 52258 56006
rect 51950 55995 52258 56004
rect 56950 56060 57258 56069
rect 56950 56058 56956 56060
rect 57012 56058 57036 56060
rect 57092 56058 57116 56060
rect 57172 56058 57196 56060
rect 57252 56058 57258 56060
rect 57012 56006 57014 56058
rect 57194 56006 57196 56058
rect 56950 56004 56956 56006
rect 57012 56004 57036 56006
rect 57092 56004 57116 56006
rect 57172 56004 57196 56006
rect 57252 56004 57258 56006
rect 56950 55995 57258 56004
rect 58532 55752 58584 55758
rect 58532 55694 58584 55700
rect 58544 55593 58572 55694
rect 58530 55584 58586 55593
rect 2610 55516 2918 55525
rect 2610 55514 2616 55516
rect 2672 55514 2696 55516
rect 2752 55514 2776 55516
rect 2832 55514 2856 55516
rect 2912 55514 2918 55516
rect 2672 55462 2674 55514
rect 2854 55462 2856 55514
rect 2610 55460 2616 55462
rect 2672 55460 2696 55462
rect 2752 55460 2776 55462
rect 2832 55460 2856 55462
rect 2912 55460 2918 55462
rect 2610 55451 2918 55460
rect 7610 55516 7918 55525
rect 7610 55514 7616 55516
rect 7672 55514 7696 55516
rect 7752 55514 7776 55516
rect 7832 55514 7856 55516
rect 7912 55514 7918 55516
rect 7672 55462 7674 55514
rect 7854 55462 7856 55514
rect 7610 55460 7616 55462
rect 7672 55460 7696 55462
rect 7752 55460 7776 55462
rect 7832 55460 7856 55462
rect 7912 55460 7918 55462
rect 7610 55451 7918 55460
rect 12610 55516 12918 55525
rect 12610 55514 12616 55516
rect 12672 55514 12696 55516
rect 12752 55514 12776 55516
rect 12832 55514 12856 55516
rect 12912 55514 12918 55516
rect 12672 55462 12674 55514
rect 12854 55462 12856 55514
rect 12610 55460 12616 55462
rect 12672 55460 12696 55462
rect 12752 55460 12776 55462
rect 12832 55460 12856 55462
rect 12912 55460 12918 55462
rect 12610 55451 12918 55460
rect 17610 55516 17918 55525
rect 17610 55514 17616 55516
rect 17672 55514 17696 55516
rect 17752 55514 17776 55516
rect 17832 55514 17856 55516
rect 17912 55514 17918 55516
rect 17672 55462 17674 55514
rect 17854 55462 17856 55514
rect 17610 55460 17616 55462
rect 17672 55460 17696 55462
rect 17752 55460 17776 55462
rect 17832 55460 17856 55462
rect 17912 55460 17918 55462
rect 17610 55451 17918 55460
rect 22610 55516 22918 55525
rect 22610 55514 22616 55516
rect 22672 55514 22696 55516
rect 22752 55514 22776 55516
rect 22832 55514 22856 55516
rect 22912 55514 22918 55516
rect 22672 55462 22674 55514
rect 22854 55462 22856 55514
rect 22610 55460 22616 55462
rect 22672 55460 22696 55462
rect 22752 55460 22776 55462
rect 22832 55460 22856 55462
rect 22912 55460 22918 55462
rect 22610 55451 22918 55460
rect 27610 55516 27918 55525
rect 27610 55514 27616 55516
rect 27672 55514 27696 55516
rect 27752 55514 27776 55516
rect 27832 55514 27856 55516
rect 27912 55514 27918 55516
rect 27672 55462 27674 55514
rect 27854 55462 27856 55514
rect 27610 55460 27616 55462
rect 27672 55460 27696 55462
rect 27752 55460 27776 55462
rect 27832 55460 27856 55462
rect 27912 55460 27918 55462
rect 27610 55451 27918 55460
rect 32610 55516 32918 55525
rect 32610 55514 32616 55516
rect 32672 55514 32696 55516
rect 32752 55514 32776 55516
rect 32832 55514 32856 55516
rect 32912 55514 32918 55516
rect 32672 55462 32674 55514
rect 32854 55462 32856 55514
rect 32610 55460 32616 55462
rect 32672 55460 32696 55462
rect 32752 55460 32776 55462
rect 32832 55460 32856 55462
rect 32912 55460 32918 55462
rect 32610 55451 32918 55460
rect 37610 55516 37918 55525
rect 37610 55514 37616 55516
rect 37672 55514 37696 55516
rect 37752 55514 37776 55516
rect 37832 55514 37856 55516
rect 37912 55514 37918 55516
rect 37672 55462 37674 55514
rect 37854 55462 37856 55514
rect 37610 55460 37616 55462
rect 37672 55460 37696 55462
rect 37752 55460 37776 55462
rect 37832 55460 37856 55462
rect 37912 55460 37918 55462
rect 37610 55451 37918 55460
rect 42610 55516 42918 55525
rect 42610 55514 42616 55516
rect 42672 55514 42696 55516
rect 42752 55514 42776 55516
rect 42832 55514 42856 55516
rect 42912 55514 42918 55516
rect 42672 55462 42674 55514
rect 42854 55462 42856 55514
rect 42610 55460 42616 55462
rect 42672 55460 42696 55462
rect 42752 55460 42776 55462
rect 42832 55460 42856 55462
rect 42912 55460 42918 55462
rect 42610 55451 42918 55460
rect 47610 55516 47918 55525
rect 47610 55514 47616 55516
rect 47672 55514 47696 55516
rect 47752 55514 47776 55516
rect 47832 55514 47856 55516
rect 47912 55514 47918 55516
rect 47672 55462 47674 55514
rect 47854 55462 47856 55514
rect 47610 55460 47616 55462
rect 47672 55460 47696 55462
rect 47752 55460 47776 55462
rect 47832 55460 47856 55462
rect 47912 55460 47918 55462
rect 47610 55451 47918 55460
rect 52610 55516 52918 55525
rect 52610 55514 52616 55516
rect 52672 55514 52696 55516
rect 52752 55514 52776 55516
rect 52832 55514 52856 55516
rect 52912 55514 52918 55516
rect 52672 55462 52674 55514
rect 52854 55462 52856 55514
rect 52610 55460 52616 55462
rect 52672 55460 52696 55462
rect 52752 55460 52776 55462
rect 52832 55460 52856 55462
rect 52912 55460 52918 55462
rect 52610 55451 52918 55460
rect 57610 55516 57918 55525
rect 58530 55519 58586 55528
rect 57610 55514 57616 55516
rect 57672 55514 57696 55516
rect 57752 55514 57776 55516
rect 57832 55514 57856 55516
rect 57912 55514 57918 55516
rect 57672 55462 57674 55514
rect 57854 55462 57856 55514
rect 57610 55460 57616 55462
rect 57672 55460 57696 55462
rect 57752 55460 57776 55462
rect 57832 55460 57856 55462
rect 57912 55460 57918 55462
rect 57610 55451 57918 55460
rect 58532 55072 58584 55078
rect 58532 55014 58584 55020
rect 1950 54972 2258 54981
rect 1950 54970 1956 54972
rect 2012 54970 2036 54972
rect 2092 54970 2116 54972
rect 2172 54970 2196 54972
rect 2252 54970 2258 54972
rect 2012 54918 2014 54970
rect 2194 54918 2196 54970
rect 1950 54916 1956 54918
rect 2012 54916 2036 54918
rect 2092 54916 2116 54918
rect 2172 54916 2196 54918
rect 2252 54916 2258 54918
rect 1950 54907 2258 54916
rect 6950 54972 7258 54981
rect 6950 54970 6956 54972
rect 7012 54970 7036 54972
rect 7092 54970 7116 54972
rect 7172 54970 7196 54972
rect 7252 54970 7258 54972
rect 7012 54918 7014 54970
rect 7194 54918 7196 54970
rect 6950 54916 6956 54918
rect 7012 54916 7036 54918
rect 7092 54916 7116 54918
rect 7172 54916 7196 54918
rect 7252 54916 7258 54918
rect 6950 54907 7258 54916
rect 11950 54972 12258 54981
rect 11950 54970 11956 54972
rect 12012 54970 12036 54972
rect 12092 54970 12116 54972
rect 12172 54970 12196 54972
rect 12252 54970 12258 54972
rect 12012 54918 12014 54970
rect 12194 54918 12196 54970
rect 11950 54916 11956 54918
rect 12012 54916 12036 54918
rect 12092 54916 12116 54918
rect 12172 54916 12196 54918
rect 12252 54916 12258 54918
rect 11950 54907 12258 54916
rect 16950 54972 17258 54981
rect 16950 54970 16956 54972
rect 17012 54970 17036 54972
rect 17092 54970 17116 54972
rect 17172 54970 17196 54972
rect 17252 54970 17258 54972
rect 17012 54918 17014 54970
rect 17194 54918 17196 54970
rect 16950 54916 16956 54918
rect 17012 54916 17036 54918
rect 17092 54916 17116 54918
rect 17172 54916 17196 54918
rect 17252 54916 17258 54918
rect 16950 54907 17258 54916
rect 21950 54972 22258 54981
rect 21950 54970 21956 54972
rect 22012 54970 22036 54972
rect 22092 54970 22116 54972
rect 22172 54970 22196 54972
rect 22252 54970 22258 54972
rect 22012 54918 22014 54970
rect 22194 54918 22196 54970
rect 21950 54916 21956 54918
rect 22012 54916 22036 54918
rect 22092 54916 22116 54918
rect 22172 54916 22196 54918
rect 22252 54916 22258 54918
rect 21950 54907 22258 54916
rect 26950 54972 27258 54981
rect 26950 54970 26956 54972
rect 27012 54970 27036 54972
rect 27092 54970 27116 54972
rect 27172 54970 27196 54972
rect 27252 54970 27258 54972
rect 27012 54918 27014 54970
rect 27194 54918 27196 54970
rect 26950 54916 26956 54918
rect 27012 54916 27036 54918
rect 27092 54916 27116 54918
rect 27172 54916 27196 54918
rect 27252 54916 27258 54918
rect 26950 54907 27258 54916
rect 31950 54972 32258 54981
rect 31950 54970 31956 54972
rect 32012 54970 32036 54972
rect 32092 54970 32116 54972
rect 32172 54970 32196 54972
rect 32252 54970 32258 54972
rect 32012 54918 32014 54970
rect 32194 54918 32196 54970
rect 31950 54916 31956 54918
rect 32012 54916 32036 54918
rect 32092 54916 32116 54918
rect 32172 54916 32196 54918
rect 32252 54916 32258 54918
rect 31950 54907 32258 54916
rect 36950 54972 37258 54981
rect 36950 54970 36956 54972
rect 37012 54970 37036 54972
rect 37092 54970 37116 54972
rect 37172 54970 37196 54972
rect 37252 54970 37258 54972
rect 37012 54918 37014 54970
rect 37194 54918 37196 54970
rect 36950 54916 36956 54918
rect 37012 54916 37036 54918
rect 37092 54916 37116 54918
rect 37172 54916 37196 54918
rect 37252 54916 37258 54918
rect 36950 54907 37258 54916
rect 41950 54972 42258 54981
rect 41950 54970 41956 54972
rect 42012 54970 42036 54972
rect 42092 54970 42116 54972
rect 42172 54970 42196 54972
rect 42252 54970 42258 54972
rect 42012 54918 42014 54970
rect 42194 54918 42196 54970
rect 41950 54916 41956 54918
rect 42012 54916 42036 54918
rect 42092 54916 42116 54918
rect 42172 54916 42196 54918
rect 42252 54916 42258 54918
rect 41950 54907 42258 54916
rect 46950 54972 47258 54981
rect 46950 54970 46956 54972
rect 47012 54970 47036 54972
rect 47092 54970 47116 54972
rect 47172 54970 47196 54972
rect 47252 54970 47258 54972
rect 47012 54918 47014 54970
rect 47194 54918 47196 54970
rect 46950 54916 46956 54918
rect 47012 54916 47036 54918
rect 47092 54916 47116 54918
rect 47172 54916 47196 54918
rect 47252 54916 47258 54918
rect 46950 54907 47258 54916
rect 51950 54972 52258 54981
rect 51950 54970 51956 54972
rect 52012 54970 52036 54972
rect 52092 54970 52116 54972
rect 52172 54970 52196 54972
rect 52252 54970 52258 54972
rect 52012 54918 52014 54970
rect 52194 54918 52196 54970
rect 51950 54916 51956 54918
rect 52012 54916 52036 54918
rect 52092 54916 52116 54918
rect 52172 54916 52196 54918
rect 52252 54916 52258 54918
rect 51950 54907 52258 54916
rect 56950 54972 57258 54981
rect 56950 54970 56956 54972
rect 57012 54970 57036 54972
rect 57092 54970 57116 54972
rect 57172 54970 57196 54972
rect 57252 54970 57258 54972
rect 57012 54918 57014 54970
rect 57194 54918 57196 54970
rect 56950 54916 56956 54918
rect 57012 54916 57036 54918
rect 57092 54916 57116 54918
rect 57172 54916 57196 54918
rect 57252 54916 57258 54918
rect 56950 54907 57258 54916
rect 58544 54777 58572 55014
rect 58530 54768 58586 54777
rect 58530 54703 58586 54712
rect 2610 54428 2918 54437
rect 2610 54426 2616 54428
rect 2672 54426 2696 54428
rect 2752 54426 2776 54428
rect 2832 54426 2856 54428
rect 2912 54426 2918 54428
rect 2672 54374 2674 54426
rect 2854 54374 2856 54426
rect 2610 54372 2616 54374
rect 2672 54372 2696 54374
rect 2752 54372 2776 54374
rect 2832 54372 2856 54374
rect 2912 54372 2918 54374
rect 2610 54363 2918 54372
rect 7610 54428 7918 54437
rect 7610 54426 7616 54428
rect 7672 54426 7696 54428
rect 7752 54426 7776 54428
rect 7832 54426 7856 54428
rect 7912 54426 7918 54428
rect 7672 54374 7674 54426
rect 7854 54374 7856 54426
rect 7610 54372 7616 54374
rect 7672 54372 7696 54374
rect 7752 54372 7776 54374
rect 7832 54372 7856 54374
rect 7912 54372 7918 54374
rect 7610 54363 7918 54372
rect 12610 54428 12918 54437
rect 12610 54426 12616 54428
rect 12672 54426 12696 54428
rect 12752 54426 12776 54428
rect 12832 54426 12856 54428
rect 12912 54426 12918 54428
rect 12672 54374 12674 54426
rect 12854 54374 12856 54426
rect 12610 54372 12616 54374
rect 12672 54372 12696 54374
rect 12752 54372 12776 54374
rect 12832 54372 12856 54374
rect 12912 54372 12918 54374
rect 12610 54363 12918 54372
rect 17610 54428 17918 54437
rect 17610 54426 17616 54428
rect 17672 54426 17696 54428
rect 17752 54426 17776 54428
rect 17832 54426 17856 54428
rect 17912 54426 17918 54428
rect 17672 54374 17674 54426
rect 17854 54374 17856 54426
rect 17610 54372 17616 54374
rect 17672 54372 17696 54374
rect 17752 54372 17776 54374
rect 17832 54372 17856 54374
rect 17912 54372 17918 54374
rect 17610 54363 17918 54372
rect 22610 54428 22918 54437
rect 22610 54426 22616 54428
rect 22672 54426 22696 54428
rect 22752 54426 22776 54428
rect 22832 54426 22856 54428
rect 22912 54426 22918 54428
rect 22672 54374 22674 54426
rect 22854 54374 22856 54426
rect 22610 54372 22616 54374
rect 22672 54372 22696 54374
rect 22752 54372 22776 54374
rect 22832 54372 22856 54374
rect 22912 54372 22918 54374
rect 22610 54363 22918 54372
rect 27610 54428 27918 54437
rect 27610 54426 27616 54428
rect 27672 54426 27696 54428
rect 27752 54426 27776 54428
rect 27832 54426 27856 54428
rect 27912 54426 27918 54428
rect 27672 54374 27674 54426
rect 27854 54374 27856 54426
rect 27610 54372 27616 54374
rect 27672 54372 27696 54374
rect 27752 54372 27776 54374
rect 27832 54372 27856 54374
rect 27912 54372 27918 54374
rect 27610 54363 27918 54372
rect 32610 54428 32918 54437
rect 32610 54426 32616 54428
rect 32672 54426 32696 54428
rect 32752 54426 32776 54428
rect 32832 54426 32856 54428
rect 32912 54426 32918 54428
rect 32672 54374 32674 54426
rect 32854 54374 32856 54426
rect 32610 54372 32616 54374
rect 32672 54372 32696 54374
rect 32752 54372 32776 54374
rect 32832 54372 32856 54374
rect 32912 54372 32918 54374
rect 32610 54363 32918 54372
rect 37610 54428 37918 54437
rect 37610 54426 37616 54428
rect 37672 54426 37696 54428
rect 37752 54426 37776 54428
rect 37832 54426 37856 54428
rect 37912 54426 37918 54428
rect 37672 54374 37674 54426
rect 37854 54374 37856 54426
rect 37610 54372 37616 54374
rect 37672 54372 37696 54374
rect 37752 54372 37776 54374
rect 37832 54372 37856 54374
rect 37912 54372 37918 54374
rect 37610 54363 37918 54372
rect 42610 54428 42918 54437
rect 42610 54426 42616 54428
rect 42672 54426 42696 54428
rect 42752 54426 42776 54428
rect 42832 54426 42856 54428
rect 42912 54426 42918 54428
rect 42672 54374 42674 54426
rect 42854 54374 42856 54426
rect 42610 54372 42616 54374
rect 42672 54372 42696 54374
rect 42752 54372 42776 54374
rect 42832 54372 42856 54374
rect 42912 54372 42918 54374
rect 42610 54363 42918 54372
rect 47610 54428 47918 54437
rect 47610 54426 47616 54428
rect 47672 54426 47696 54428
rect 47752 54426 47776 54428
rect 47832 54426 47856 54428
rect 47912 54426 47918 54428
rect 47672 54374 47674 54426
rect 47854 54374 47856 54426
rect 47610 54372 47616 54374
rect 47672 54372 47696 54374
rect 47752 54372 47776 54374
rect 47832 54372 47856 54374
rect 47912 54372 47918 54374
rect 47610 54363 47918 54372
rect 52610 54428 52918 54437
rect 52610 54426 52616 54428
rect 52672 54426 52696 54428
rect 52752 54426 52776 54428
rect 52832 54426 52856 54428
rect 52912 54426 52918 54428
rect 52672 54374 52674 54426
rect 52854 54374 52856 54426
rect 52610 54372 52616 54374
rect 52672 54372 52696 54374
rect 52752 54372 52776 54374
rect 52832 54372 52856 54374
rect 52912 54372 52918 54374
rect 52610 54363 52918 54372
rect 57610 54428 57918 54437
rect 57610 54426 57616 54428
rect 57672 54426 57696 54428
rect 57752 54426 57776 54428
rect 57832 54426 57856 54428
rect 57912 54426 57918 54428
rect 57672 54374 57674 54426
rect 57854 54374 57856 54426
rect 57610 54372 57616 54374
rect 57672 54372 57696 54374
rect 57752 54372 57776 54374
rect 57832 54372 57856 54374
rect 57912 54372 57918 54374
rect 57610 54363 57918 54372
rect 58532 53984 58584 53990
rect 58530 53952 58532 53961
rect 58584 53952 58586 53961
rect 1950 53884 2258 53893
rect 1950 53882 1956 53884
rect 2012 53882 2036 53884
rect 2092 53882 2116 53884
rect 2172 53882 2196 53884
rect 2252 53882 2258 53884
rect 2012 53830 2014 53882
rect 2194 53830 2196 53882
rect 1950 53828 1956 53830
rect 2012 53828 2036 53830
rect 2092 53828 2116 53830
rect 2172 53828 2196 53830
rect 2252 53828 2258 53830
rect 1950 53819 2258 53828
rect 6950 53884 7258 53893
rect 6950 53882 6956 53884
rect 7012 53882 7036 53884
rect 7092 53882 7116 53884
rect 7172 53882 7196 53884
rect 7252 53882 7258 53884
rect 7012 53830 7014 53882
rect 7194 53830 7196 53882
rect 6950 53828 6956 53830
rect 7012 53828 7036 53830
rect 7092 53828 7116 53830
rect 7172 53828 7196 53830
rect 7252 53828 7258 53830
rect 6950 53819 7258 53828
rect 11950 53884 12258 53893
rect 11950 53882 11956 53884
rect 12012 53882 12036 53884
rect 12092 53882 12116 53884
rect 12172 53882 12196 53884
rect 12252 53882 12258 53884
rect 12012 53830 12014 53882
rect 12194 53830 12196 53882
rect 11950 53828 11956 53830
rect 12012 53828 12036 53830
rect 12092 53828 12116 53830
rect 12172 53828 12196 53830
rect 12252 53828 12258 53830
rect 11950 53819 12258 53828
rect 16950 53884 17258 53893
rect 16950 53882 16956 53884
rect 17012 53882 17036 53884
rect 17092 53882 17116 53884
rect 17172 53882 17196 53884
rect 17252 53882 17258 53884
rect 17012 53830 17014 53882
rect 17194 53830 17196 53882
rect 16950 53828 16956 53830
rect 17012 53828 17036 53830
rect 17092 53828 17116 53830
rect 17172 53828 17196 53830
rect 17252 53828 17258 53830
rect 16950 53819 17258 53828
rect 21950 53884 22258 53893
rect 21950 53882 21956 53884
rect 22012 53882 22036 53884
rect 22092 53882 22116 53884
rect 22172 53882 22196 53884
rect 22252 53882 22258 53884
rect 22012 53830 22014 53882
rect 22194 53830 22196 53882
rect 21950 53828 21956 53830
rect 22012 53828 22036 53830
rect 22092 53828 22116 53830
rect 22172 53828 22196 53830
rect 22252 53828 22258 53830
rect 21950 53819 22258 53828
rect 26950 53884 27258 53893
rect 26950 53882 26956 53884
rect 27012 53882 27036 53884
rect 27092 53882 27116 53884
rect 27172 53882 27196 53884
rect 27252 53882 27258 53884
rect 27012 53830 27014 53882
rect 27194 53830 27196 53882
rect 26950 53828 26956 53830
rect 27012 53828 27036 53830
rect 27092 53828 27116 53830
rect 27172 53828 27196 53830
rect 27252 53828 27258 53830
rect 26950 53819 27258 53828
rect 31950 53884 32258 53893
rect 31950 53882 31956 53884
rect 32012 53882 32036 53884
rect 32092 53882 32116 53884
rect 32172 53882 32196 53884
rect 32252 53882 32258 53884
rect 32012 53830 32014 53882
rect 32194 53830 32196 53882
rect 31950 53828 31956 53830
rect 32012 53828 32036 53830
rect 32092 53828 32116 53830
rect 32172 53828 32196 53830
rect 32252 53828 32258 53830
rect 31950 53819 32258 53828
rect 36950 53884 37258 53893
rect 36950 53882 36956 53884
rect 37012 53882 37036 53884
rect 37092 53882 37116 53884
rect 37172 53882 37196 53884
rect 37252 53882 37258 53884
rect 37012 53830 37014 53882
rect 37194 53830 37196 53882
rect 36950 53828 36956 53830
rect 37012 53828 37036 53830
rect 37092 53828 37116 53830
rect 37172 53828 37196 53830
rect 37252 53828 37258 53830
rect 36950 53819 37258 53828
rect 41950 53884 42258 53893
rect 41950 53882 41956 53884
rect 42012 53882 42036 53884
rect 42092 53882 42116 53884
rect 42172 53882 42196 53884
rect 42252 53882 42258 53884
rect 42012 53830 42014 53882
rect 42194 53830 42196 53882
rect 41950 53828 41956 53830
rect 42012 53828 42036 53830
rect 42092 53828 42116 53830
rect 42172 53828 42196 53830
rect 42252 53828 42258 53830
rect 41950 53819 42258 53828
rect 46950 53884 47258 53893
rect 46950 53882 46956 53884
rect 47012 53882 47036 53884
rect 47092 53882 47116 53884
rect 47172 53882 47196 53884
rect 47252 53882 47258 53884
rect 47012 53830 47014 53882
rect 47194 53830 47196 53882
rect 46950 53828 46956 53830
rect 47012 53828 47036 53830
rect 47092 53828 47116 53830
rect 47172 53828 47196 53830
rect 47252 53828 47258 53830
rect 46950 53819 47258 53828
rect 51950 53884 52258 53893
rect 51950 53882 51956 53884
rect 52012 53882 52036 53884
rect 52092 53882 52116 53884
rect 52172 53882 52196 53884
rect 52252 53882 52258 53884
rect 52012 53830 52014 53882
rect 52194 53830 52196 53882
rect 51950 53828 51956 53830
rect 52012 53828 52036 53830
rect 52092 53828 52116 53830
rect 52172 53828 52196 53830
rect 52252 53828 52258 53830
rect 51950 53819 52258 53828
rect 56950 53884 57258 53893
rect 58530 53887 58586 53896
rect 56950 53882 56956 53884
rect 57012 53882 57036 53884
rect 57092 53882 57116 53884
rect 57172 53882 57196 53884
rect 57252 53882 57258 53884
rect 57012 53830 57014 53882
rect 57194 53830 57196 53882
rect 56950 53828 56956 53830
rect 57012 53828 57036 53830
rect 57092 53828 57116 53830
rect 57172 53828 57196 53830
rect 57252 53828 57258 53830
rect 56950 53819 57258 53828
rect 58532 53576 58584 53582
rect 58532 53518 58584 53524
rect 2610 53340 2918 53349
rect 2610 53338 2616 53340
rect 2672 53338 2696 53340
rect 2752 53338 2776 53340
rect 2832 53338 2856 53340
rect 2912 53338 2918 53340
rect 2672 53286 2674 53338
rect 2854 53286 2856 53338
rect 2610 53284 2616 53286
rect 2672 53284 2696 53286
rect 2752 53284 2776 53286
rect 2832 53284 2856 53286
rect 2912 53284 2918 53286
rect 2610 53275 2918 53284
rect 7610 53340 7918 53349
rect 7610 53338 7616 53340
rect 7672 53338 7696 53340
rect 7752 53338 7776 53340
rect 7832 53338 7856 53340
rect 7912 53338 7918 53340
rect 7672 53286 7674 53338
rect 7854 53286 7856 53338
rect 7610 53284 7616 53286
rect 7672 53284 7696 53286
rect 7752 53284 7776 53286
rect 7832 53284 7856 53286
rect 7912 53284 7918 53286
rect 7610 53275 7918 53284
rect 12610 53340 12918 53349
rect 12610 53338 12616 53340
rect 12672 53338 12696 53340
rect 12752 53338 12776 53340
rect 12832 53338 12856 53340
rect 12912 53338 12918 53340
rect 12672 53286 12674 53338
rect 12854 53286 12856 53338
rect 12610 53284 12616 53286
rect 12672 53284 12696 53286
rect 12752 53284 12776 53286
rect 12832 53284 12856 53286
rect 12912 53284 12918 53286
rect 12610 53275 12918 53284
rect 17610 53340 17918 53349
rect 17610 53338 17616 53340
rect 17672 53338 17696 53340
rect 17752 53338 17776 53340
rect 17832 53338 17856 53340
rect 17912 53338 17918 53340
rect 17672 53286 17674 53338
rect 17854 53286 17856 53338
rect 17610 53284 17616 53286
rect 17672 53284 17696 53286
rect 17752 53284 17776 53286
rect 17832 53284 17856 53286
rect 17912 53284 17918 53286
rect 17610 53275 17918 53284
rect 22610 53340 22918 53349
rect 22610 53338 22616 53340
rect 22672 53338 22696 53340
rect 22752 53338 22776 53340
rect 22832 53338 22856 53340
rect 22912 53338 22918 53340
rect 22672 53286 22674 53338
rect 22854 53286 22856 53338
rect 22610 53284 22616 53286
rect 22672 53284 22696 53286
rect 22752 53284 22776 53286
rect 22832 53284 22856 53286
rect 22912 53284 22918 53286
rect 22610 53275 22918 53284
rect 27610 53340 27918 53349
rect 27610 53338 27616 53340
rect 27672 53338 27696 53340
rect 27752 53338 27776 53340
rect 27832 53338 27856 53340
rect 27912 53338 27918 53340
rect 27672 53286 27674 53338
rect 27854 53286 27856 53338
rect 27610 53284 27616 53286
rect 27672 53284 27696 53286
rect 27752 53284 27776 53286
rect 27832 53284 27856 53286
rect 27912 53284 27918 53286
rect 27610 53275 27918 53284
rect 32610 53340 32918 53349
rect 32610 53338 32616 53340
rect 32672 53338 32696 53340
rect 32752 53338 32776 53340
rect 32832 53338 32856 53340
rect 32912 53338 32918 53340
rect 32672 53286 32674 53338
rect 32854 53286 32856 53338
rect 32610 53284 32616 53286
rect 32672 53284 32696 53286
rect 32752 53284 32776 53286
rect 32832 53284 32856 53286
rect 32912 53284 32918 53286
rect 32610 53275 32918 53284
rect 37610 53340 37918 53349
rect 37610 53338 37616 53340
rect 37672 53338 37696 53340
rect 37752 53338 37776 53340
rect 37832 53338 37856 53340
rect 37912 53338 37918 53340
rect 37672 53286 37674 53338
rect 37854 53286 37856 53338
rect 37610 53284 37616 53286
rect 37672 53284 37696 53286
rect 37752 53284 37776 53286
rect 37832 53284 37856 53286
rect 37912 53284 37918 53286
rect 37610 53275 37918 53284
rect 42610 53340 42918 53349
rect 42610 53338 42616 53340
rect 42672 53338 42696 53340
rect 42752 53338 42776 53340
rect 42832 53338 42856 53340
rect 42912 53338 42918 53340
rect 42672 53286 42674 53338
rect 42854 53286 42856 53338
rect 42610 53284 42616 53286
rect 42672 53284 42696 53286
rect 42752 53284 42776 53286
rect 42832 53284 42856 53286
rect 42912 53284 42918 53286
rect 42610 53275 42918 53284
rect 47610 53340 47918 53349
rect 47610 53338 47616 53340
rect 47672 53338 47696 53340
rect 47752 53338 47776 53340
rect 47832 53338 47856 53340
rect 47912 53338 47918 53340
rect 47672 53286 47674 53338
rect 47854 53286 47856 53338
rect 47610 53284 47616 53286
rect 47672 53284 47696 53286
rect 47752 53284 47776 53286
rect 47832 53284 47856 53286
rect 47912 53284 47918 53286
rect 47610 53275 47918 53284
rect 52610 53340 52918 53349
rect 52610 53338 52616 53340
rect 52672 53338 52696 53340
rect 52752 53338 52776 53340
rect 52832 53338 52856 53340
rect 52912 53338 52918 53340
rect 52672 53286 52674 53338
rect 52854 53286 52856 53338
rect 52610 53284 52616 53286
rect 52672 53284 52696 53286
rect 52752 53284 52776 53286
rect 52832 53284 52856 53286
rect 52912 53284 52918 53286
rect 52610 53275 52918 53284
rect 57610 53340 57918 53349
rect 57610 53338 57616 53340
rect 57672 53338 57696 53340
rect 57752 53338 57776 53340
rect 57832 53338 57856 53340
rect 57912 53338 57918 53340
rect 57672 53286 57674 53338
rect 57854 53286 57856 53338
rect 57610 53284 57616 53286
rect 57672 53284 57696 53286
rect 57752 53284 57776 53286
rect 57832 53284 57856 53286
rect 57912 53284 57918 53286
rect 57610 53275 57918 53284
rect 58544 53145 58572 53518
rect 58530 53136 58586 53145
rect 58530 53071 58586 53080
rect 1950 52796 2258 52805
rect 1950 52794 1956 52796
rect 2012 52794 2036 52796
rect 2092 52794 2116 52796
rect 2172 52794 2196 52796
rect 2252 52794 2258 52796
rect 2012 52742 2014 52794
rect 2194 52742 2196 52794
rect 1950 52740 1956 52742
rect 2012 52740 2036 52742
rect 2092 52740 2116 52742
rect 2172 52740 2196 52742
rect 2252 52740 2258 52742
rect 1950 52731 2258 52740
rect 6950 52796 7258 52805
rect 6950 52794 6956 52796
rect 7012 52794 7036 52796
rect 7092 52794 7116 52796
rect 7172 52794 7196 52796
rect 7252 52794 7258 52796
rect 7012 52742 7014 52794
rect 7194 52742 7196 52794
rect 6950 52740 6956 52742
rect 7012 52740 7036 52742
rect 7092 52740 7116 52742
rect 7172 52740 7196 52742
rect 7252 52740 7258 52742
rect 6950 52731 7258 52740
rect 11950 52796 12258 52805
rect 11950 52794 11956 52796
rect 12012 52794 12036 52796
rect 12092 52794 12116 52796
rect 12172 52794 12196 52796
rect 12252 52794 12258 52796
rect 12012 52742 12014 52794
rect 12194 52742 12196 52794
rect 11950 52740 11956 52742
rect 12012 52740 12036 52742
rect 12092 52740 12116 52742
rect 12172 52740 12196 52742
rect 12252 52740 12258 52742
rect 11950 52731 12258 52740
rect 16950 52796 17258 52805
rect 16950 52794 16956 52796
rect 17012 52794 17036 52796
rect 17092 52794 17116 52796
rect 17172 52794 17196 52796
rect 17252 52794 17258 52796
rect 17012 52742 17014 52794
rect 17194 52742 17196 52794
rect 16950 52740 16956 52742
rect 17012 52740 17036 52742
rect 17092 52740 17116 52742
rect 17172 52740 17196 52742
rect 17252 52740 17258 52742
rect 16950 52731 17258 52740
rect 21950 52796 22258 52805
rect 21950 52794 21956 52796
rect 22012 52794 22036 52796
rect 22092 52794 22116 52796
rect 22172 52794 22196 52796
rect 22252 52794 22258 52796
rect 22012 52742 22014 52794
rect 22194 52742 22196 52794
rect 21950 52740 21956 52742
rect 22012 52740 22036 52742
rect 22092 52740 22116 52742
rect 22172 52740 22196 52742
rect 22252 52740 22258 52742
rect 21950 52731 22258 52740
rect 26950 52796 27258 52805
rect 26950 52794 26956 52796
rect 27012 52794 27036 52796
rect 27092 52794 27116 52796
rect 27172 52794 27196 52796
rect 27252 52794 27258 52796
rect 27012 52742 27014 52794
rect 27194 52742 27196 52794
rect 26950 52740 26956 52742
rect 27012 52740 27036 52742
rect 27092 52740 27116 52742
rect 27172 52740 27196 52742
rect 27252 52740 27258 52742
rect 26950 52731 27258 52740
rect 31950 52796 32258 52805
rect 31950 52794 31956 52796
rect 32012 52794 32036 52796
rect 32092 52794 32116 52796
rect 32172 52794 32196 52796
rect 32252 52794 32258 52796
rect 32012 52742 32014 52794
rect 32194 52742 32196 52794
rect 31950 52740 31956 52742
rect 32012 52740 32036 52742
rect 32092 52740 32116 52742
rect 32172 52740 32196 52742
rect 32252 52740 32258 52742
rect 31950 52731 32258 52740
rect 36950 52796 37258 52805
rect 36950 52794 36956 52796
rect 37012 52794 37036 52796
rect 37092 52794 37116 52796
rect 37172 52794 37196 52796
rect 37252 52794 37258 52796
rect 37012 52742 37014 52794
rect 37194 52742 37196 52794
rect 36950 52740 36956 52742
rect 37012 52740 37036 52742
rect 37092 52740 37116 52742
rect 37172 52740 37196 52742
rect 37252 52740 37258 52742
rect 36950 52731 37258 52740
rect 41950 52796 42258 52805
rect 41950 52794 41956 52796
rect 42012 52794 42036 52796
rect 42092 52794 42116 52796
rect 42172 52794 42196 52796
rect 42252 52794 42258 52796
rect 42012 52742 42014 52794
rect 42194 52742 42196 52794
rect 41950 52740 41956 52742
rect 42012 52740 42036 52742
rect 42092 52740 42116 52742
rect 42172 52740 42196 52742
rect 42252 52740 42258 52742
rect 41950 52731 42258 52740
rect 46950 52796 47258 52805
rect 46950 52794 46956 52796
rect 47012 52794 47036 52796
rect 47092 52794 47116 52796
rect 47172 52794 47196 52796
rect 47252 52794 47258 52796
rect 47012 52742 47014 52794
rect 47194 52742 47196 52794
rect 46950 52740 46956 52742
rect 47012 52740 47036 52742
rect 47092 52740 47116 52742
rect 47172 52740 47196 52742
rect 47252 52740 47258 52742
rect 46950 52731 47258 52740
rect 51950 52796 52258 52805
rect 51950 52794 51956 52796
rect 52012 52794 52036 52796
rect 52092 52794 52116 52796
rect 52172 52794 52196 52796
rect 52252 52794 52258 52796
rect 52012 52742 52014 52794
rect 52194 52742 52196 52794
rect 51950 52740 51956 52742
rect 52012 52740 52036 52742
rect 52092 52740 52116 52742
rect 52172 52740 52196 52742
rect 52252 52740 52258 52742
rect 51950 52731 52258 52740
rect 56950 52796 57258 52805
rect 56950 52794 56956 52796
rect 57012 52794 57036 52796
rect 57092 52794 57116 52796
rect 57172 52794 57196 52796
rect 57252 52794 57258 52796
rect 57012 52742 57014 52794
rect 57194 52742 57196 52794
rect 56950 52740 56956 52742
rect 57012 52740 57036 52742
rect 57092 52740 57116 52742
rect 57172 52740 57196 52742
rect 57252 52740 57258 52742
rect 56950 52731 57258 52740
rect 58532 52488 58584 52494
rect 58532 52430 58584 52436
rect 58544 52329 58572 52430
rect 58530 52320 58586 52329
rect 2610 52252 2918 52261
rect 2610 52250 2616 52252
rect 2672 52250 2696 52252
rect 2752 52250 2776 52252
rect 2832 52250 2856 52252
rect 2912 52250 2918 52252
rect 2672 52198 2674 52250
rect 2854 52198 2856 52250
rect 2610 52196 2616 52198
rect 2672 52196 2696 52198
rect 2752 52196 2776 52198
rect 2832 52196 2856 52198
rect 2912 52196 2918 52198
rect 2610 52187 2918 52196
rect 7610 52252 7918 52261
rect 7610 52250 7616 52252
rect 7672 52250 7696 52252
rect 7752 52250 7776 52252
rect 7832 52250 7856 52252
rect 7912 52250 7918 52252
rect 7672 52198 7674 52250
rect 7854 52198 7856 52250
rect 7610 52196 7616 52198
rect 7672 52196 7696 52198
rect 7752 52196 7776 52198
rect 7832 52196 7856 52198
rect 7912 52196 7918 52198
rect 7610 52187 7918 52196
rect 12610 52252 12918 52261
rect 12610 52250 12616 52252
rect 12672 52250 12696 52252
rect 12752 52250 12776 52252
rect 12832 52250 12856 52252
rect 12912 52250 12918 52252
rect 12672 52198 12674 52250
rect 12854 52198 12856 52250
rect 12610 52196 12616 52198
rect 12672 52196 12696 52198
rect 12752 52196 12776 52198
rect 12832 52196 12856 52198
rect 12912 52196 12918 52198
rect 12610 52187 12918 52196
rect 17610 52252 17918 52261
rect 17610 52250 17616 52252
rect 17672 52250 17696 52252
rect 17752 52250 17776 52252
rect 17832 52250 17856 52252
rect 17912 52250 17918 52252
rect 17672 52198 17674 52250
rect 17854 52198 17856 52250
rect 17610 52196 17616 52198
rect 17672 52196 17696 52198
rect 17752 52196 17776 52198
rect 17832 52196 17856 52198
rect 17912 52196 17918 52198
rect 17610 52187 17918 52196
rect 22610 52252 22918 52261
rect 22610 52250 22616 52252
rect 22672 52250 22696 52252
rect 22752 52250 22776 52252
rect 22832 52250 22856 52252
rect 22912 52250 22918 52252
rect 22672 52198 22674 52250
rect 22854 52198 22856 52250
rect 22610 52196 22616 52198
rect 22672 52196 22696 52198
rect 22752 52196 22776 52198
rect 22832 52196 22856 52198
rect 22912 52196 22918 52198
rect 22610 52187 22918 52196
rect 27610 52252 27918 52261
rect 27610 52250 27616 52252
rect 27672 52250 27696 52252
rect 27752 52250 27776 52252
rect 27832 52250 27856 52252
rect 27912 52250 27918 52252
rect 27672 52198 27674 52250
rect 27854 52198 27856 52250
rect 27610 52196 27616 52198
rect 27672 52196 27696 52198
rect 27752 52196 27776 52198
rect 27832 52196 27856 52198
rect 27912 52196 27918 52198
rect 27610 52187 27918 52196
rect 32610 52252 32918 52261
rect 32610 52250 32616 52252
rect 32672 52250 32696 52252
rect 32752 52250 32776 52252
rect 32832 52250 32856 52252
rect 32912 52250 32918 52252
rect 32672 52198 32674 52250
rect 32854 52198 32856 52250
rect 32610 52196 32616 52198
rect 32672 52196 32696 52198
rect 32752 52196 32776 52198
rect 32832 52196 32856 52198
rect 32912 52196 32918 52198
rect 32610 52187 32918 52196
rect 37610 52252 37918 52261
rect 37610 52250 37616 52252
rect 37672 52250 37696 52252
rect 37752 52250 37776 52252
rect 37832 52250 37856 52252
rect 37912 52250 37918 52252
rect 37672 52198 37674 52250
rect 37854 52198 37856 52250
rect 37610 52196 37616 52198
rect 37672 52196 37696 52198
rect 37752 52196 37776 52198
rect 37832 52196 37856 52198
rect 37912 52196 37918 52198
rect 37610 52187 37918 52196
rect 42610 52252 42918 52261
rect 42610 52250 42616 52252
rect 42672 52250 42696 52252
rect 42752 52250 42776 52252
rect 42832 52250 42856 52252
rect 42912 52250 42918 52252
rect 42672 52198 42674 52250
rect 42854 52198 42856 52250
rect 42610 52196 42616 52198
rect 42672 52196 42696 52198
rect 42752 52196 42776 52198
rect 42832 52196 42856 52198
rect 42912 52196 42918 52198
rect 42610 52187 42918 52196
rect 47610 52252 47918 52261
rect 47610 52250 47616 52252
rect 47672 52250 47696 52252
rect 47752 52250 47776 52252
rect 47832 52250 47856 52252
rect 47912 52250 47918 52252
rect 47672 52198 47674 52250
rect 47854 52198 47856 52250
rect 47610 52196 47616 52198
rect 47672 52196 47696 52198
rect 47752 52196 47776 52198
rect 47832 52196 47856 52198
rect 47912 52196 47918 52198
rect 47610 52187 47918 52196
rect 52610 52252 52918 52261
rect 52610 52250 52616 52252
rect 52672 52250 52696 52252
rect 52752 52250 52776 52252
rect 52832 52250 52856 52252
rect 52912 52250 52918 52252
rect 52672 52198 52674 52250
rect 52854 52198 52856 52250
rect 52610 52196 52616 52198
rect 52672 52196 52696 52198
rect 52752 52196 52776 52198
rect 52832 52196 52856 52198
rect 52912 52196 52918 52198
rect 52610 52187 52918 52196
rect 57610 52252 57918 52261
rect 58530 52255 58586 52264
rect 57610 52250 57616 52252
rect 57672 52250 57696 52252
rect 57752 52250 57776 52252
rect 57832 52250 57856 52252
rect 57912 52250 57918 52252
rect 57672 52198 57674 52250
rect 57854 52198 57856 52250
rect 57610 52196 57616 52198
rect 57672 52196 57696 52198
rect 57752 52196 57776 52198
rect 57832 52196 57856 52198
rect 57912 52196 57918 52198
rect 57610 52187 57918 52196
rect 58532 51808 58584 51814
rect 58532 51750 58584 51756
rect 1950 51708 2258 51717
rect 1950 51706 1956 51708
rect 2012 51706 2036 51708
rect 2092 51706 2116 51708
rect 2172 51706 2196 51708
rect 2252 51706 2258 51708
rect 2012 51654 2014 51706
rect 2194 51654 2196 51706
rect 1950 51652 1956 51654
rect 2012 51652 2036 51654
rect 2092 51652 2116 51654
rect 2172 51652 2196 51654
rect 2252 51652 2258 51654
rect 1950 51643 2258 51652
rect 6950 51708 7258 51717
rect 6950 51706 6956 51708
rect 7012 51706 7036 51708
rect 7092 51706 7116 51708
rect 7172 51706 7196 51708
rect 7252 51706 7258 51708
rect 7012 51654 7014 51706
rect 7194 51654 7196 51706
rect 6950 51652 6956 51654
rect 7012 51652 7036 51654
rect 7092 51652 7116 51654
rect 7172 51652 7196 51654
rect 7252 51652 7258 51654
rect 6950 51643 7258 51652
rect 11950 51708 12258 51717
rect 11950 51706 11956 51708
rect 12012 51706 12036 51708
rect 12092 51706 12116 51708
rect 12172 51706 12196 51708
rect 12252 51706 12258 51708
rect 12012 51654 12014 51706
rect 12194 51654 12196 51706
rect 11950 51652 11956 51654
rect 12012 51652 12036 51654
rect 12092 51652 12116 51654
rect 12172 51652 12196 51654
rect 12252 51652 12258 51654
rect 11950 51643 12258 51652
rect 16950 51708 17258 51717
rect 16950 51706 16956 51708
rect 17012 51706 17036 51708
rect 17092 51706 17116 51708
rect 17172 51706 17196 51708
rect 17252 51706 17258 51708
rect 17012 51654 17014 51706
rect 17194 51654 17196 51706
rect 16950 51652 16956 51654
rect 17012 51652 17036 51654
rect 17092 51652 17116 51654
rect 17172 51652 17196 51654
rect 17252 51652 17258 51654
rect 16950 51643 17258 51652
rect 21950 51708 22258 51717
rect 21950 51706 21956 51708
rect 22012 51706 22036 51708
rect 22092 51706 22116 51708
rect 22172 51706 22196 51708
rect 22252 51706 22258 51708
rect 22012 51654 22014 51706
rect 22194 51654 22196 51706
rect 21950 51652 21956 51654
rect 22012 51652 22036 51654
rect 22092 51652 22116 51654
rect 22172 51652 22196 51654
rect 22252 51652 22258 51654
rect 21950 51643 22258 51652
rect 26950 51708 27258 51717
rect 26950 51706 26956 51708
rect 27012 51706 27036 51708
rect 27092 51706 27116 51708
rect 27172 51706 27196 51708
rect 27252 51706 27258 51708
rect 27012 51654 27014 51706
rect 27194 51654 27196 51706
rect 26950 51652 26956 51654
rect 27012 51652 27036 51654
rect 27092 51652 27116 51654
rect 27172 51652 27196 51654
rect 27252 51652 27258 51654
rect 26950 51643 27258 51652
rect 31950 51708 32258 51717
rect 31950 51706 31956 51708
rect 32012 51706 32036 51708
rect 32092 51706 32116 51708
rect 32172 51706 32196 51708
rect 32252 51706 32258 51708
rect 32012 51654 32014 51706
rect 32194 51654 32196 51706
rect 31950 51652 31956 51654
rect 32012 51652 32036 51654
rect 32092 51652 32116 51654
rect 32172 51652 32196 51654
rect 32252 51652 32258 51654
rect 31950 51643 32258 51652
rect 36950 51708 37258 51717
rect 36950 51706 36956 51708
rect 37012 51706 37036 51708
rect 37092 51706 37116 51708
rect 37172 51706 37196 51708
rect 37252 51706 37258 51708
rect 37012 51654 37014 51706
rect 37194 51654 37196 51706
rect 36950 51652 36956 51654
rect 37012 51652 37036 51654
rect 37092 51652 37116 51654
rect 37172 51652 37196 51654
rect 37252 51652 37258 51654
rect 36950 51643 37258 51652
rect 41950 51708 42258 51717
rect 41950 51706 41956 51708
rect 42012 51706 42036 51708
rect 42092 51706 42116 51708
rect 42172 51706 42196 51708
rect 42252 51706 42258 51708
rect 42012 51654 42014 51706
rect 42194 51654 42196 51706
rect 41950 51652 41956 51654
rect 42012 51652 42036 51654
rect 42092 51652 42116 51654
rect 42172 51652 42196 51654
rect 42252 51652 42258 51654
rect 41950 51643 42258 51652
rect 46950 51708 47258 51717
rect 46950 51706 46956 51708
rect 47012 51706 47036 51708
rect 47092 51706 47116 51708
rect 47172 51706 47196 51708
rect 47252 51706 47258 51708
rect 47012 51654 47014 51706
rect 47194 51654 47196 51706
rect 46950 51652 46956 51654
rect 47012 51652 47036 51654
rect 47092 51652 47116 51654
rect 47172 51652 47196 51654
rect 47252 51652 47258 51654
rect 46950 51643 47258 51652
rect 51950 51708 52258 51717
rect 51950 51706 51956 51708
rect 52012 51706 52036 51708
rect 52092 51706 52116 51708
rect 52172 51706 52196 51708
rect 52252 51706 52258 51708
rect 52012 51654 52014 51706
rect 52194 51654 52196 51706
rect 51950 51652 51956 51654
rect 52012 51652 52036 51654
rect 52092 51652 52116 51654
rect 52172 51652 52196 51654
rect 52252 51652 52258 51654
rect 51950 51643 52258 51652
rect 56950 51708 57258 51717
rect 56950 51706 56956 51708
rect 57012 51706 57036 51708
rect 57092 51706 57116 51708
rect 57172 51706 57196 51708
rect 57252 51706 57258 51708
rect 57012 51654 57014 51706
rect 57194 51654 57196 51706
rect 56950 51652 56956 51654
rect 57012 51652 57036 51654
rect 57092 51652 57116 51654
rect 57172 51652 57196 51654
rect 57252 51652 57258 51654
rect 56950 51643 57258 51652
rect 58544 51513 58572 51750
rect 58530 51504 58586 51513
rect 58530 51439 58586 51448
rect 2610 51164 2918 51173
rect 2610 51162 2616 51164
rect 2672 51162 2696 51164
rect 2752 51162 2776 51164
rect 2832 51162 2856 51164
rect 2912 51162 2918 51164
rect 2672 51110 2674 51162
rect 2854 51110 2856 51162
rect 2610 51108 2616 51110
rect 2672 51108 2696 51110
rect 2752 51108 2776 51110
rect 2832 51108 2856 51110
rect 2912 51108 2918 51110
rect 2610 51099 2918 51108
rect 7610 51164 7918 51173
rect 7610 51162 7616 51164
rect 7672 51162 7696 51164
rect 7752 51162 7776 51164
rect 7832 51162 7856 51164
rect 7912 51162 7918 51164
rect 7672 51110 7674 51162
rect 7854 51110 7856 51162
rect 7610 51108 7616 51110
rect 7672 51108 7696 51110
rect 7752 51108 7776 51110
rect 7832 51108 7856 51110
rect 7912 51108 7918 51110
rect 7610 51099 7918 51108
rect 12610 51164 12918 51173
rect 12610 51162 12616 51164
rect 12672 51162 12696 51164
rect 12752 51162 12776 51164
rect 12832 51162 12856 51164
rect 12912 51162 12918 51164
rect 12672 51110 12674 51162
rect 12854 51110 12856 51162
rect 12610 51108 12616 51110
rect 12672 51108 12696 51110
rect 12752 51108 12776 51110
rect 12832 51108 12856 51110
rect 12912 51108 12918 51110
rect 12610 51099 12918 51108
rect 17610 51164 17918 51173
rect 17610 51162 17616 51164
rect 17672 51162 17696 51164
rect 17752 51162 17776 51164
rect 17832 51162 17856 51164
rect 17912 51162 17918 51164
rect 17672 51110 17674 51162
rect 17854 51110 17856 51162
rect 17610 51108 17616 51110
rect 17672 51108 17696 51110
rect 17752 51108 17776 51110
rect 17832 51108 17856 51110
rect 17912 51108 17918 51110
rect 17610 51099 17918 51108
rect 22610 51164 22918 51173
rect 22610 51162 22616 51164
rect 22672 51162 22696 51164
rect 22752 51162 22776 51164
rect 22832 51162 22856 51164
rect 22912 51162 22918 51164
rect 22672 51110 22674 51162
rect 22854 51110 22856 51162
rect 22610 51108 22616 51110
rect 22672 51108 22696 51110
rect 22752 51108 22776 51110
rect 22832 51108 22856 51110
rect 22912 51108 22918 51110
rect 22610 51099 22918 51108
rect 27610 51164 27918 51173
rect 27610 51162 27616 51164
rect 27672 51162 27696 51164
rect 27752 51162 27776 51164
rect 27832 51162 27856 51164
rect 27912 51162 27918 51164
rect 27672 51110 27674 51162
rect 27854 51110 27856 51162
rect 27610 51108 27616 51110
rect 27672 51108 27696 51110
rect 27752 51108 27776 51110
rect 27832 51108 27856 51110
rect 27912 51108 27918 51110
rect 27610 51099 27918 51108
rect 32610 51164 32918 51173
rect 32610 51162 32616 51164
rect 32672 51162 32696 51164
rect 32752 51162 32776 51164
rect 32832 51162 32856 51164
rect 32912 51162 32918 51164
rect 32672 51110 32674 51162
rect 32854 51110 32856 51162
rect 32610 51108 32616 51110
rect 32672 51108 32696 51110
rect 32752 51108 32776 51110
rect 32832 51108 32856 51110
rect 32912 51108 32918 51110
rect 32610 51099 32918 51108
rect 37610 51164 37918 51173
rect 37610 51162 37616 51164
rect 37672 51162 37696 51164
rect 37752 51162 37776 51164
rect 37832 51162 37856 51164
rect 37912 51162 37918 51164
rect 37672 51110 37674 51162
rect 37854 51110 37856 51162
rect 37610 51108 37616 51110
rect 37672 51108 37696 51110
rect 37752 51108 37776 51110
rect 37832 51108 37856 51110
rect 37912 51108 37918 51110
rect 37610 51099 37918 51108
rect 42610 51164 42918 51173
rect 42610 51162 42616 51164
rect 42672 51162 42696 51164
rect 42752 51162 42776 51164
rect 42832 51162 42856 51164
rect 42912 51162 42918 51164
rect 42672 51110 42674 51162
rect 42854 51110 42856 51162
rect 42610 51108 42616 51110
rect 42672 51108 42696 51110
rect 42752 51108 42776 51110
rect 42832 51108 42856 51110
rect 42912 51108 42918 51110
rect 42610 51099 42918 51108
rect 47610 51164 47918 51173
rect 47610 51162 47616 51164
rect 47672 51162 47696 51164
rect 47752 51162 47776 51164
rect 47832 51162 47856 51164
rect 47912 51162 47918 51164
rect 47672 51110 47674 51162
rect 47854 51110 47856 51162
rect 47610 51108 47616 51110
rect 47672 51108 47696 51110
rect 47752 51108 47776 51110
rect 47832 51108 47856 51110
rect 47912 51108 47918 51110
rect 47610 51099 47918 51108
rect 52610 51164 52918 51173
rect 52610 51162 52616 51164
rect 52672 51162 52696 51164
rect 52752 51162 52776 51164
rect 52832 51162 52856 51164
rect 52912 51162 52918 51164
rect 52672 51110 52674 51162
rect 52854 51110 52856 51162
rect 52610 51108 52616 51110
rect 52672 51108 52696 51110
rect 52752 51108 52776 51110
rect 52832 51108 52856 51110
rect 52912 51108 52918 51110
rect 52610 51099 52918 51108
rect 57610 51164 57918 51173
rect 57610 51162 57616 51164
rect 57672 51162 57696 51164
rect 57752 51162 57776 51164
rect 57832 51162 57856 51164
rect 57912 51162 57918 51164
rect 57672 51110 57674 51162
rect 57854 51110 57856 51162
rect 57610 51108 57616 51110
rect 57672 51108 57696 51110
rect 57752 51108 57776 51110
rect 57832 51108 57856 51110
rect 57912 51108 57918 51110
rect 57610 51099 57918 51108
rect 58532 50720 58584 50726
rect 58530 50688 58532 50697
rect 58584 50688 58586 50697
rect 1950 50620 2258 50629
rect 1950 50618 1956 50620
rect 2012 50618 2036 50620
rect 2092 50618 2116 50620
rect 2172 50618 2196 50620
rect 2252 50618 2258 50620
rect 2012 50566 2014 50618
rect 2194 50566 2196 50618
rect 1950 50564 1956 50566
rect 2012 50564 2036 50566
rect 2092 50564 2116 50566
rect 2172 50564 2196 50566
rect 2252 50564 2258 50566
rect 1950 50555 2258 50564
rect 6950 50620 7258 50629
rect 6950 50618 6956 50620
rect 7012 50618 7036 50620
rect 7092 50618 7116 50620
rect 7172 50618 7196 50620
rect 7252 50618 7258 50620
rect 7012 50566 7014 50618
rect 7194 50566 7196 50618
rect 6950 50564 6956 50566
rect 7012 50564 7036 50566
rect 7092 50564 7116 50566
rect 7172 50564 7196 50566
rect 7252 50564 7258 50566
rect 6950 50555 7258 50564
rect 11950 50620 12258 50629
rect 11950 50618 11956 50620
rect 12012 50618 12036 50620
rect 12092 50618 12116 50620
rect 12172 50618 12196 50620
rect 12252 50618 12258 50620
rect 12012 50566 12014 50618
rect 12194 50566 12196 50618
rect 11950 50564 11956 50566
rect 12012 50564 12036 50566
rect 12092 50564 12116 50566
rect 12172 50564 12196 50566
rect 12252 50564 12258 50566
rect 11950 50555 12258 50564
rect 16950 50620 17258 50629
rect 16950 50618 16956 50620
rect 17012 50618 17036 50620
rect 17092 50618 17116 50620
rect 17172 50618 17196 50620
rect 17252 50618 17258 50620
rect 17012 50566 17014 50618
rect 17194 50566 17196 50618
rect 16950 50564 16956 50566
rect 17012 50564 17036 50566
rect 17092 50564 17116 50566
rect 17172 50564 17196 50566
rect 17252 50564 17258 50566
rect 16950 50555 17258 50564
rect 21950 50620 22258 50629
rect 21950 50618 21956 50620
rect 22012 50618 22036 50620
rect 22092 50618 22116 50620
rect 22172 50618 22196 50620
rect 22252 50618 22258 50620
rect 22012 50566 22014 50618
rect 22194 50566 22196 50618
rect 21950 50564 21956 50566
rect 22012 50564 22036 50566
rect 22092 50564 22116 50566
rect 22172 50564 22196 50566
rect 22252 50564 22258 50566
rect 21950 50555 22258 50564
rect 26950 50620 27258 50629
rect 26950 50618 26956 50620
rect 27012 50618 27036 50620
rect 27092 50618 27116 50620
rect 27172 50618 27196 50620
rect 27252 50618 27258 50620
rect 27012 50566 27014 50618
rect 27194 50566 27196 50618
rect 26950 50564 26956 50566
rect 27012 50564 27036 50566
rect 27092 50564 27116 50566
rect 27172 50564 27196 50566
rect 27252 50564 27258 50566
rect 26950 50555 27258 50564
rect 31950 50620 32258 50629
rect 31950 50618 31956 50620
rect 32012 50618 32036 50620
rect 32092 50618 32116 50620
rect 32172 50618 32196 50620
rect 32252 50618 32258 50620
rect 32012 50566 32014 50618
rect 32194 50566 32196 50618
rect 31950 50564 31956 50566
rect 32012 50564 32036 50566
rect 32092 50564 32116 50566
rect 32172 50564 32196 50566
rect 32252 50564 32258 50566
rect 31950 50555 32258 50564
rect 36950 50620 37258 50629
rect 36950 50618 36956 50620
rect 37012 50618 37036 50620
rect 37092 50618 37116 50620
rect 37172 50618 37196 50620
rect 37252 50618 37258 50620
rect 37012 50566 37014 50618
rect 37194 50566 37196 50618
rect 36950 50564 36956 50566
rect 37012 50564 37036 50566
rect 37092 50564 37116 50566
rect 37172 50564 37196 50566
rect 37252 50564 37258 50566
rect 36950 50555 37258 50564
rect 41950 50620 42258 50629
rect 41950 50618 41956 50620
rect 42012 50618 42036 50620
rect 42092 50618 42116 50620
rect 42172 50618 42196 50620
rect 42252 50618 42258 50620
rect 42012 50566 42014 50618
rect 42194 50566 42196 50618
rect 41950 50564 41956 50566
rect 42012 50564 42036 50566
rect 42092 50564 42116 50566
rect 42172 50564 42196 50566
rect 42252 50564 42258 50566
rect 41950 50555 42258 50564
rect 46950 50620 47258 50629
rect 46950 50618 46956 50620
rect 47012 50618 47036 50620
rect 47092 50618 47116 50620
rect 47172 50618 47196 50620
rect 47252 50618 47258 50620
rect 47012 50566 47014 50618
rect 47194 50566 47196 50618
rect 46950 50564 46956 50566
rect 47012 50564 47036 50566
rect 47092 50564 47116 50566
rect 47172 50564 47196 50566
rect 47252 50564 47258 50566
rect 46950 50555 47258 50564
rect 51950 50620 52258 50629
rect 51950 50618 51956 50620
rect 52012 50618 52036 50620
rect 52092 50618 52116 50620
rect 52172 50618 52196 50620
rect 52252 50618 52258 50620
rect 52012 50566 52014 50618
rect 52194 50566 52196 50618
rect 51950 50564 51956 50566
rect 52012 50564 52036 50566
rect 52092 50564 52116 50566
rect 52172 50564 52196 50566
rect 52252 50564 52258 50566
rect 51950 50555 52258 50564
rect 56950 50620 57258 50629
rect 58530 50623 58586 50632
rect 56950 50618 56956 50620
rect 57012 50618 57036 50620
rect 57092 50618 57116 50620
rect 57172 50618 57196 50620
rect 57252 50618 57258 50620
rect 57012 50566 57014 50618
rect 57194 50566 57196 50618
rect 56950 50564 56956 50566
rect 57012 50564 57036 50566
rect 57092 50564 57116 50566
rect 57172 50564 57196 50566
rect 57252 50564 57258 50566
rect 56950 50555 57258 50564
rect 58532 50312 58584 50318
rect 58532 50254 58584 50260
rect 2610 50076 2918 50085
rect 2610 50074 2616 50076
rect 2672 50074 2696 50076
rect 2752 50074 2776 50076
rect 2832 50074 2856 50076
rect 2912 50074 2918 50076
rect 2672 50022 2674 50074
rect 2854 50022 2856 50074
rect 2610 50020 2616 50022
rect 2672 50020 2696 50022
rect 2752 50020 2776 50022
rect 2832 50020 2856 50022
rect 2912 50020 2918 50022
rect 2610 50011 2918 50020
rect 7610 50076 7918 50085
rect 7610 50074 7616 50076
rect 7672 50074 7696 50076
rect 7752 50074 7776 50076
rect 7832 50074 7856 50076
rect 7912 50074 7918 50076
rect 7672 50022 7674 50074
rect 7854 50022 7856 50074
rect 7610 50020 7616 50022
rect 7672 50020 7696 50022
rect 7752 50020 7776 50022
rect 7832 50020 7856 50022
rect 7912 50020 7918 50022
rect 7610 50011 7918 50020
rect 12610 50076 12918 50085
rect 12610 50074 12616 50076
rect 12672 50074 12696 50076
rect 12752 50074 12776 50076
rect 12832 50074 12856 50076
rect 12912 50074 12918 50076
rect 12672 50022 12674 50074
rect 12854 50022 12856 50074
rect 12610 50020 12616 50022
rect 12672 50020 12696 50022
rect 12752 50020 12776 50022
rect 12832 50020 12856 50022
rect 12912 50020 12918 50022
rect 12610 50011 12918 50020
rect 17610 50076 17918 50085
rect 17610 50074 17616 50076
rect 17672 50074 17696 50076
rect 17752 50074 17776 50076
rect 17832 50074 17856 50076
rect 17912 50074 17918 50076
rect 17672 50022 17674 50074
rect 17854 50022 17856 50074
rect 17610 50020 17616 50022
rect 17672 50020 17696 50022
rect 17752 50020 17776 50022
rect 17832 50020 17856 50022
rect 17912 50020 17918 50022
rect 17610 50011 17918 50020
rect 22610 50076 22918 50085
rect 22610 50074 22616 50076
rect 22672 50074 22696 50076
rect 22752 50074 22776 50076
rect 22832 50074 22856 50076
rect 22912 50074 22918 50076
rect 22672 50022 22674 50074
rect 22854 50022 22856 50074
rect 22610 50020 22616 50022
rect 22672 50020 22696 50022
rect 22752 50020 22776 50022
rect 22832 50020 22856 50022
rect 22912 50020 22918 50022
rect 22610 50011 22918 50020
rect 27610 50076 27918 50085
rect 27610 50074 27616 50076
rect 27672 50074 27696 50076
rect 27752 50074 27776 50076
rect 27832 50074 27856 50076
rect 27912 50074 27918 50076
rect 27672 50022 27674 50074
rect 27854 50022 27856 50074
rect 27610 50020 27616 50022
rect 27672 50020 27696 50022
rect 27752 50020 27776 50022
rect 27832 50020 27856 50022
rect 27912 50020 27918 50022
rect 27610 50011 27918 50020
rect 32610 50076 32918 50085
rect 32610 50074 32616 50076
rect 32672 50074 32696 50076
rect 32752 50074 32776 50076
rect 32832 50074 32856 50076
rect 32912 50074 32918 50076
rect 32672 50022 32674 50074
rect 32854 50022 32856 50074
rect 32610 50020 32616 50022
rect 32672 50020 32696 50022
rect 32752 50020 32776 50022
rect 32832 50020 32856 50022
rect 32912 50020 32918 50022
rect 32610 50011 32918 50020
rect 37610 50076 37918 50085
rect 37610 50074 37616 50076
rect 37672 50074 37696 50076
rect 37752 50074 37776 50076
rect 37832 50074 37856 50076
rect 37912 50074 37918 50076
rect 37672 50022 37674 50074
rect 37854 50022 37856 50074
rect 37610 50020 37616 50022
rect 37672 50020 37696 50022
rect 37752 50020 37776 50022
rect 37832 50020 37856 50022
rect 37912 50020 37918 50022
rect 37610 50011 37918 50020
rect 42610 50076 42918 50085
rect 42610 50074 42616 50076
rect 42672 50074 42696 50076
rect 42752 50074 42776 50076
rect 42832 50074 42856 50076
rect 42912 50074 42918 50076
rect 42672 50022 42674 50074
rect 42854 50022 42856 50074
rect 42610 50020 42616 50022
rect 42672 50020 42696 50022
rect 42752 50020 42776 50022
rect 42832 50020 42856 50022
rect 42912 50020 42918 50022
rect 42610 50011 42918 50020
rect 47610 50076 47918 50085
rect 47610 50074 47616 50076
rect 47672 50074 47696 50076
rect 47752 50074 47776 50076
rect 47832 50074 47856 50076
rect 47912 50074 47918 50076
rect 47672 50022 47674 50074
rect 47854 50022 47856 50074
rect 47610 50020 47616 50022
rect 47672 50020 47696 50022
rect 47752 50020 47776 50022
rect 47832 50020 47856 50022
rect 47912 50020 47918 50022
rect 47610 50011 47918 50020
rect 52610 50076 52918 50085
rect 52610 50074 52616 50076
rect 52672 50074 52696 50076
rect 52752 50074 52776 50076
rect 52832 50074 52856 50076
rect 52912 50074 52918 50076
rect 52672 50022 52674 50074
rect 52854 50022 52856 50074
rect 52610 50020 52616 50022
rect 52672 50020 52696 50022
rect 52752 50020 52776 50022
rect 52832 50020 52856 50022
rect 52912 50020 52918 50022
rect 52610 50011 52918 50020
rect 57610 50076 57918 50085
rect 57610 50074 57616 50076
rect 57672 50074 57696 50076
rect 57752 50074 57776 50076
rect 57832 50074 57856 50076
rect 57912 50074 57918 50076
rect 57672 50022 57674 50074
rect 57854 50022 57856 50074
rect 57610 50020 57616 50022
rect 57672 50020 57696 50022
rect 57752 50020 57776 50022
rect 57832 50020 57856 50022
rect 57912 50020 57918 50022
rect 57610 50011 57918 50020
rect 58544 49881 58572 50254
rect 58530 49872 58586 49881
rect 58530 49807 58586 49816
rect 1950 49532 2258 49541
rect 1950 49530 1956 49532
rect 2012 49530 2036 49532
rect 2092 49530 2116 49532
rect 2172 49530 2196 49532
rect 2252 49530 2258 49532
rect 2012 49478 2014 49530
rect 2194 49478 2196 49530
rect 1950 49476 1956 49478
rect 2012 49476 2036 49478
rect 2092 49476 2116 49478
rect 2172 49476 2196 49478
rect 2252 49476 2258 49478
rect 1950 49467 2258 49476
rect 6950 49532 7258 49541
rect 6950 49530 6956 49532
rect 7012 49530 7036 49532
rect 7092 49530 7116 49532
rect 7172 49530 7196 49532
rect 7252 49530 7258 49532
rect 7012 49478 7014 49530
rect 7194 49478 7196 49530
rect 6950 49476 6956 49478
rect 7012 49476 7036 49478
rect 7092 49476 7116 49478
rect 7172 49476 7196 49478
rect 7252 49476 7258 49478
rect 6950 49467 7258 49476
rect 11950 49532 12258 49541
rect 11950 49530 11956 49532
rect 12012 49530 12036 49532
rect 12092 49530 12116 49532
rect 12172 49530 12196 49532
rect 12252 49530 12258 49532
rect 12012 49478 12014 49530
rect 12194 49478 12196 49530
rect 11950 49476 11956 49478
rect 12012 49476 12036 49478
rect 12092 49476 12116 49478
rect 12172 49476 12196 49478
rect 12252 49476 12258 49478
rect 11950 49467 12258 49476
rect 16950 49532 17258 49541
rect 16950 49530 16956 49532
rect 17012 49530 17036 49532
rect 17092 49530 17116 49532
rect 17172 49530 17196 49532
rect 17252 49530 17258 49532
rect 17012 49478 17014 49530
rect 17194 49478 17196 49530
rect 16950 49476 16956 49478
rect 17012 49476 17036 49478
rect 17092 49476 17116 49478
rect 17172 49476 17196 49478
rect 17252 49476 17258 49478
rect 16950 49467 17258 49476
rect 21950 49532 22258 49541
rect 21950 49530 21956 49532
rect 22012 49530 22036 49532
rect 22092 49530 22116 49532
rect 22172 49530 22196 49532
rect 22252 49530 22258 49532
rect 22012 49478 22014 49530
rect 22194 49478 22196 49530
rect 21950 49476 21956 49478
rect 22012 49476 22036 49478
rect 22092 49476 22116 49478
rect 22172 49476 22196 49478
rect 22252 49476 22258 49478
rect 21950 49467 22258 49476
rect 26950 49532 27258 49541
rect 26950 49530 26956 49532
rect 27012 49530 27036 49532
rect 27092 49530 27116 49532
rect 27172 49530 27196 49532
rect 27252 49530 27258 49532
rect 27012 49478 27014 49530
rect 27194 49478 27196 49530
rect 26950 49476 26956 49478
rect 27012 49476 27036 49478
rect 27092 49476 27116 49478
rect 27172 49476 27196 49478
rect 27252 49476 27258 49478
rect 26950 49467 27258 49476
rect 31950 49532 32258 49541
rect 31950 49530 31956 49532
rect 32012 49530 32036 49532
rect 32092 49530 32116 49532
rect 32172 49530 32196 49532
rect 32252 49530 32258 49532
rect 32012 49478 32014 49530
rect 32194 49478 32196 49530
rect 31950 49476 31956 49478
rect 32012 49476 32036 49478
rect 32092 49476 32116 49478
rect 32172 49476 32196 49478
rect 32252 49476 32258 49478
rect 31950 49467 32258 49476
rect 36950 49532 37258 49541
rect 36950 49530 36956 49532
rect 37012 49530 37036 49532
rect 37092 49530 37116 49532
rect 37172 49530 37196 49532
rect 37252 49530 37258 49532
rect 37012 49478 37014 49530
rect 37194 49478 37196 49530
rect 36950 49476 36956 49478
rect 37012 49476 37036 49478
rect 37092 49476 37116 49478
rect 37172 49476 37196 49478
rect 37252 49476 37258 49478
rect 36950 49467 37258 49476
rect 41950 49532 42258 49541
rect 41950 49530 41956 49532
rect 42012 49530 42036 49532
rect 42092 49530 42116 49532
rect 42172 49530 42196 49532
rect 42252 49530 42258 49532
rect 42012 49478 42014 49530
rect 42194 49478 42196 49530
rect 41950 49476 41956 49478
rect 42012 49476 42036 49478
rect 42092 49476 42116 49478
rect 42172 49476 42196 49478
rect 42252 49476 42258 49478
rect 41950 49467 42258 49476
rect 46950 49532 47258 49541
rect 46950 49530 46956 49532
rect 47012 49530 47036 49532
rect 47092 49530 47116 49532
rect 47172 49530 47196 49532
rect 47252 49530 47258 49532
rect 47012 49478 47014 49530
rect 47194 49478 47196 49530
rect 46950 49476 46956 49478
rect 47012 49476 47036 49478
rect 47092 49476 47116 49478
rect 47172 49476 47196 49478
rect 47252 49476 47258 49478
rect 46950 49467 47258 49476
rect 51950 49532 52258 49541
rect 51950 49530 51956 49532
rect 52012 49530 52036 49532
rect 52092 49530 52116 49532
rect 52172 49530 52196 49532
rect 52252 49530 52258 49532
rect 52012 49478 52014 49530
rect 52194 49478 52196 49530
rect 51950 49476 51956 49478
rect 52012 49476 52036 49478
rect 52092 49476 52116 49478
rect 52172 49476 52196 49478
rect 52252 49476 52258 49478
rect 51950 49467 52258 49476
rect 56950 49532 57258 49541
rect 56950 49530 56956 49532
rect 57012 49530 57036 49532
rect 57092 49530 57116 49532
rect 57172 49530 57196 49532
rect 57252 49530 57258 49532
rect 57012 49478 57014 49530
rect 57194 49478 57196 49530
rect 56950 49476 56956 49478
rect 57012 49476 57036 49478
rect 57092 49476 57116 49478
rect 57172 49476 57196 49478
rect 57252 49476 57258 49478
rect 56950 49467 57258 49476
rect 58532 49224 58584 49230
rect 58532 49166 58584 49172
rect 58544 49065 58572 49166
rect 58530 49056 58586 49065
rect 2610 48988 2918 48997
rect 2610 48986 2616 48988
rect 2672 48986 2696 48988
rect 2752 48986 2776 48988
rect 2832 48986 2856 48988
rect 2912 48986 2918 48988
rect 2672 48934 2674 48986
rect 2854 48934 2856 48986
rect 2610 48932 2616 48934
rect 2672 48932 2696 48934
rect 2752 48932 2776 48934
rect 2832 48932 2856 48934
rect 2912 48932 2918 48934
rect 2610 48923 2918 48932
rect 7610 48988 7918 48997
rect 7610 48986 7616 48988
rect 7672 48986 7696 48988
rect 7752 48986 7776 48988
rect 7832 48986 7856 48988
rect 7912 48986 7918 48988
rect 7672 48934 7674 48986
rect 7854 48934 7856 48986
rect 7610 48932 7616 48934
rect 7672 48932 7696 48934
rect 7752 48932 7776 48934
rect 7832 48932 7856 48934
rect 7912 48932 7918 48934
rect 7610 48923 7918 48932
rect 12610 48988 12918 48997
rect 12610 48986 12616 48988
rect 12672 48986 12696 48988
rect 12752 48986 12776 48988
rect 12832 48986 12856 48988
rect 12912 48986 12918 48988
rect 12672 48934 12674 48986
rect 12854 48934 12856 48986
rect 12610 48932 12616 48934
rect 12672 48932 12696 48934
rect 12752 48932 12776 48934
rect 12832 48932 12856 48934
rect 12912 48932 12918 48934
rect 12610 48923 12918 48932
rect 17610 48988 17918 48997
rect 17610 48986 17616 48988
rect 17672 48986 17696 48988
rect 17752 48986 17776 48988
rect 17832 48986 17856 48988
rect 17912 48986 17918 48988
rect 17672 48934 17674 48986
rect 17854 48934 17856 48986
rect 17610 48932 17616 48934
rect 17672 48932 17696 48934
rect 17752 48932 17776 48934
rect 17832 48932 17856 48934
rect 17912 48932 17918 48934
rect 17610 48923 17918 48932
rect 22610 48988 22918 48997
rect 22610 48986 22616 48988
rect 22672 48986 22696 48988
rect 22752 48986 22776 48988
rect 22832 48986 22856 48988
rect 22912 48986 22918 48988
rect 22672 48934 22674 48986
rect 22854 48934 22856 48986
rect 22610 48932 22616 48934
rect 22672 48932 22696 48934
rect 22752 48932 22776 48934
rect 22832 48932 22856 48934
rect 22912 48932 22918 48934
rect 22610 48923 22918 48932
rect 27610 48988 27918 48997
rect 27610 48986 27616 48988
rect 27672 48986 27696 48988
rect 27752 48986 27776 48988
rect 27832 48986 27856 48988
rect 27912 48986 27918 48988
rect 27672 48934 27674 48986
rect 27854 48934 27856 48986
rect 27610 48932 27616 48934
rect 27672 48932 27696 48934
rect 27752 48932 27776 48934
rect 27832 48932 27856 48934
rect 27912 48932 27918 48934
rect 27610 48923 27918 48932
rect 32610 48988 32918 48997
rect 32610 48986 32616 48988
rect 32672 48986 32696 48988
rect 32752 48986 32776 48988
rect 32832 48986 32856 48988
rect 32912 48986 32918 48988
rect 32672 48934 32674 48986
rect 32854 48934 32856 48986
rect 32610 48932 32616 48934
rect 32672 48932 32696 48934
rect 32752 48932 32776 48934
rect 32832 48932 32856 48934
rect 32912 48932 32918 48934
rect 32610 48923 32918 48932
rect 37610 48988 37918 48997
rect 37610 48986 37616 48988
rect 37672 48986 37696 48988
rect 37752 48986 37776 48988
rect 37832 48986 37856 48988
rect 37912 48986 37918 48988
rect 37672 48934 37674 48986
rect 37854 48934 37856 48986
rect 37610 48932 37616 48934
rect 37672 48932 37696 48934
rect 37752 48932 37776 48934
rect 37832 48932 37856 48934
rect 37912 48932 37918 48934
rect 37610 48923 37918 48932
rect 42610 48988 42918 48997
rect 42610 48986 42616 48988
rect 42672 48986 42696 48988
rect 42752 48986 42776 48988
rect 42832 48986 42856 48988
rect 42912 48986 42918 48988
rect 42672 48934 42674 48986
rect 42854 48934 42856 48986
rect 42610 48932 42616 48934
rect 42672 48932 42696 48934
rect 42752 48932 42776 48934
rect 42832 48932 42856 48934
rect 42912 48932 42918 48934
rect 42610 48923 42918 48932
rect 47610 48988 47918 48997
rect 47610 48986 47616 48988
rect 47672 48986 47696 48988
rect 47752 48986 47776 48988
rect 47832 48986 47856 48988
rect 47912 48986 47918 48988
rect 47672 48934 47674 48986
rect 47854 48934 47856 48986
rect 47610 48932 47616 48934
rect 47672 48932 47696 48934
rect 47752 48932 47776 48934
rect 47832 48932 47856 48934
rect 47912 48932 47918 48934
rect 47610 48923 47918 48932
rect 52610 48988 52918 48997
rect 52610 48986 52616 48988
rect 52672 48986 52696 48988
rect 52752 48986 52776 48988
rect 52832 48986 52856 48988
rect 52912 48986 52918 48988
rect 52672 48934 52674 48986
rect 52854 48934 52856 48986
rect 52610 48932 52616 48934
rect 52672 48932 52696 48934
rect 52752 48932 52776 48934
rect 52832 48932 52856 48934
rect 52912 48932 52918 48934
rect 52610 48923 52918 48932
rect 57610 48988 57918 48997
rect 58530 48991 58586 49000
rect 57610 48986 57616 48988
rect 57672 48986 57696 48988
rect 57752 48986 57776 48988
rect 57832 48986 57856 48988
rect 57912 48986 57918 48988
rect 57672 48934 57674 48986
rect 57854 48934 57856 48986
rect 57610 48932 57616 48934
rect 57672 48932 57696 48934
rect 57752 48932 57776 48934
rect 57832 48932 57856 48934
rect 57912 48932 57918 48934
rect 57610 48923 57918 48932
rect 58532 48544 58584 48550
rect 58532 48486 58584 48492
rect 1950 48444 2258 48453
rect 1950 48442 1956 48444
rect 2012 48442 2036 48444
rect 2092 48442 2116 48444
rect 2172 48442 2196 48444
rect 2252 48442 2258 48444
rect 2012 48390 2014 48442
rect 2194 48390 2196 48442
rect 1950 48388 1956 48390
rect 2012 48388 2036 48390
rect 2092 48388 2116 48390
rect 2172 48388 2196 48390
rect 2252 48388 2258 48390
rect 1950 48379 2258 48388
rect 6950 48444 7258 48453
rect 6950 48442 6956 48444
rect 7012 48442 7036 48444
rect 7092 48442 7116 48444
rect 7172 48442 7196 48444
rect 7252 48442 7258 48444
rect 7012 48390 7014 48442
rect 7194 48390 7196 48442
rect 6950 48388 6956 48390
rect 7012 48388 7036 48390
rect 7092 48388 7116 48390
rect 7172 48388 7196 48390
rect 7252 48388 7258 48390
rect 6950 48379 7258 48388
rect 11950 48444 12258 48453
rect 11950 48442 11956 48444
rect 12012 48442 12036 48444
rect 12092 48442 12116 48444
rect 12172 48442 12196 48444
rect 12252 48442 12258 48444
rect 12012 48390 12014 48442
rect 12194 48390 12196 48442
rect 11950 48388 11956 48390
rect 12012 48388 12036 48390
rect 12092 48388 12116 48390
rect 12172 48388 12196 48390
rect 12252 48388 12258 48390
rect 11950 48379 12258 48388
rect 16950 48444 17258 48453
rect 16950 48442 16956 48444
rect 17012 48442 17036 48444
rect 17092 48442 17116 48444
rect 17172 48442 17196 48444
rect 17252 48442 17258 48444
rect 17012 48390 17014 48442
rect 17194 48390 17196 48442
rect 16950 48388 16956 48390
rect 17012 48388 17036 48390
rect 17092 48388 17116 48390
rect 17172 48388 17196 48390
rect 17252 48388 17258 48390
rect 16950 48379 17258 48388
rect 21950 48444 22258 48453
rect 21950 48442 21956 48444
rect 22012 48442 22036 48444
rect 22092 48442 22116 48444
rect 22172 48442 22196 48444
rect 22252 48442 22258 48444
rect 22012 48390 22014 48442
rect 22194 48390 22196 48442
rect 21950 48388 21956 48390
rect 22012 48388 22036 48390
rect 22092 48388 22116 48390
rect 22172 48388 22196 48390
rect 22252 48388 22258 48390
rect 21950 48379 22258 48388
rect 26950 48444 27258 48453
rect 26950 48442 26956 48444
rect 27012 48442 27036 48444
rect 27092 48442 27116 48444
rect 27172 48442 27196 48444
rect 27252 48442 27258 48444
rect 27012 48390 27014 48442
rect 27194 48390 27196 48442
rect 26950 48388 26956 48390
rect 27012 48388 27036 48390
rect 27092 48388 27116 48390
rect 27172 48388 27196 48390
rect 27252 48388 27258 48390
rect 26950 48379 27258 48388
rect 31950 48444 32258 48453
rect 31950 48442 31956 48444
rect 32012 48442 32036 48444
rect 32092 48442 32116 48444
rect 32172 48442 32196 48444
rect 32252 48442 32258 48444
rect 32012 48390 32014 48442
rect 32194 48390 32196 48442
rect 31950 48388 31956 48390
rect 32012 48388 32036 48390
rect 32092 48388 32116 48390
rect 32172 48388 32196 48390
rect 32252 48388 32258 48390
rect 31950 48379 32258 48388
rect 36950 48444 37258 48453
rect 36950 48442 36956 48444
rect 37012 48442 37036 48444
rect 37092 48442 37116 48444
rect 37172 48442 37196 48444
rect 37252 48442 37258 48444
rect 37012 48390 37014 48442
rect 37194 48390 37196 48442
rect 36950 48388 36956 48390
rect 37012 48388 37036 48390
rect 37092 48388 37116 48390
rect 37172 48388 37196 48390
rect 37252 48388 37258 48390
rect 36950 48379 37258 48388
rect 41950 48444 42258 48453
rect 41950 48442 41956 48444
rect 42012 48442 42036 48444
rect 42092 48442 42116 48444
rect 42172 48442 42196 48444
rect 42252 48442 42258 48444
rect 42012 48390 42014 48442
rect 42194 48390 42196 48442
rect 41950 48388 41956 48390
rect 42012 48388 42036 48390
rect 42092 48388 42116 48390
rect 42172 48388 42196 48390
rect 42252 48388 42258 48390
rect 41950 48379 42258 48388
rect 46950 48444 47258 48453
rect 46950 48442 46956 48444
rect 47012 48442 47036 48444
rect 47092 48442 47116 48444
rect 47172 48442 47196 48444
rect 47252 48442 47258 48444
rect 47012 48390 47014 48442
rect 47194 48390 47196 48442
rect 46950 48388 46956 48390
rect 47012 48388 47036 48390
rect 47092 48388 47116 48390
rect 47172 48388 47196 48390
rect 47252 48388 47258 48390
rect 46950 48379 47258 48388
rect 51950 48444 52258 48453
rect 51950 48442 51956 48444
rect 52012 48442 52036 48444
rect 52092 48442 52116 48444
rect 52172 48442 52196 48444
rect 52252 48442 52258 48444
rect 52012 48390 52014 48442
rect 52194 48390 52196 48442
rect 51950 48388 51956 48390
rect 52012 48388 52036 48390
rect 52092 48388 52116 48390
rect 52172 48388 52196 48390
rect 52252 48388 52258 48390
rect 51950 48379 52258 48388
rect 56950 48444 57258 48453
rect 56950 48442 56956 48444
rect 57012 48442 57036 48444
rect 57092 48442 57116 48444
rect 57172 48442 57196 48444
rect 57252 48442 57258 48444
rect 57012 48390 57014 48442
rect 57194 48390 57196 48442
rect 56950 48388 56956 48390
rect 57012 48388 57036 48390
rect 57092 48388 57116 48390
rect 57172 48388 57196 48390
rect 57252 48388 57258 48390
rect 56950 48379 57258 48388
rect 58544 48249 58572 48486
rect 58530 48240 58586 48249
rect 58530 48175 58586 48184
rect 2610 47900 2918 47909
rect 2610 47898 2616 47900
rect 2672 47898 2696 47900
rect 2752 47898 2776 47900
rect 2832 47898 2856 47900
rect 2912 47898 2918 47900
rect 2672 47846 2674 47898
rect 2854 47846 2856 47898
rect 2610 47844 2616 47846
rect 2672 47844 2696 47846
rect 2752 47844 2776 47846
rect 2832 47844 2856 47846
rect 2912 47844 2918 47846
rect 2610 47835 2918 47844
rect 7610 47900 7918 47909
rect 7610 47898 7616 47900
rect 7672 47898 7696 47900
rect 7752 47898 7776 47900
rect 7832 47898 7856 47900
rect 7912 47898 7918 47900
rect 7672 47846 7674 47898
rect 7854 47846 7856 47898
rect 7610 47844 7616 47846
rect 7672 47844 7696 47846
rect 7752 47844 7776 47846
rect 7832 47844 7856 47846
rect 7912 47844 7918 47846
rect 7610 47835 7918 47844
rect 12610 47900 12918 47909
rect 12610 47898 12616 47900
rect 12672 47898 12696 47900
rect 12752 47898 12776 47900
rect 12832 47898 12856 47900
rect 12912 47898 12918 47900
rect 12672 47846 12674 47898
rect 12854 47846 12856 47898
rect 12610 47844 12616 47846
rect 12672 47844 12696 47846
rect 12752 47844 12776 47846
rect 12832 47844 12856 47846
rect 12912 47844 12918 47846
rect 12610 47835 12918 47844
rect 17610 47900 17918 47909
rect 17610 47898 17616 47900
rect 17672 47898 17696 47900
rect 17752 47898 17776 47900
rect 17832 47898 17856 47900
rect 17912 47898 17918 47900
rect 17672 47846 17674 47898
rect 17854 47846 17856 47898
rect 17610 47844 17616 47846
rect 17672 47844 17696 47846
rect 17752 47844 17776 47846
rect 17832 47844 17856 47846
rect 17912 47844 17918 47846
rect 17610 47835 17918 47844
rect 22610 47900 22918 47909
rect 22610 47898 22616 47900
rect 22672 47898 22696 47900
rect 22752 47898 22776 47900
rect 22832 47898 22856 47900
rect 22912 47898 22918 47900
rect 22672 47846 22674 47898
rect 22854 47846 22856 47898
rect 22610 47844 22616 47846
rect 22672 47844 22696 47846
rect 22752 47844 22776 47846
rect 22832 47844 22856 47846
rect 22912 47844 22918 47846
rect 22610 47835 22918 47844
rect 27610 47900 27918 47909
rect 27610 47898 27616 47900
rect 27672 47898 27696 47900
rect 27752 47898 27776 47900
rect 27832 47898 27856 47900
rect 27912 47898 27918 47900
rect 27672 47846 27674 47898
rect 27854 47846 27856 47898
rect 27610 47844 27616 47846
rect 27672 47844 27696 47846
rect 27752 47844 27776 47846
rect 27832 47844 27856 47846
rect 27912 47844 27918 47846
rect 27610 47835 27918 47844
rect 32610 47900 32918 47909
rect 32610 47898 32616 47900
rect 32672 47898 32696 47900
rect 32752 47898 32776 47900
rect 32832 47898 32856 47900
rect 32912 47898 32918 47900
rect 32672 47846 32674 47898
rect 32854 47846 32856 47898
rect 32610 47844 32616 47846
rect 32672 47844 32696 47846
rect 32752 47844 32776 47846
rect 32832 47844 32856 47846
rect 32912 47844 32918 47846
rect 32610 47835 32918 47844
rect 37610 47900 37918 47909
rect 37610 47898 37616 47900
rect 37672 47898 37696 47900
rect 37752 47898 37776 47900
rect 37832 47898 37856 47900
rect 37912 47898 37918 47900
rect 37672 47846 37674 47898
rect 37854 47846 37856 47898
rect 37610 47844 37616 47846
rect 37672 47844 37696 47846
rect 37752 47844 37776 47846
rect 37832 47844 37856 47846
rect 37912 47844 37918 47846
rect 37610 47835 37918 47844
rect 42610 47900 42918 47909
rect 42610 47898 42616 47900
rect 42672 47898 42696 47900
rect 42752 47898 42776 47900
rect 42832 47898 42856 47900
rect 42912 47898 42918 47900
rect 42672 47846 42674 47898
rect 42854 47846 42856 47898
rect 42610 47844 42616 47846
rect 42672 47844 42696 47846
rect 42752 47844 42776 47846
rect 42832 47844 42856 47846
rect 42912 47844 42918 47846
rect 42610 47835 42918 47844
rect 47610 47900 47918 47909
rect 47610 47898 47616 47900
rect 47672 47898 47696 47900
rect 47752 47898 47776 47900
rect 47832 47898 47856 47900
rect 47912 47898 47918 47900
rect 47672 47846 47674 47898
rect 47854 47846 47856 47898
rect 47610 47844 47616 47846
rect 47672 47844 47696 47846
rect 47752 47844 47776 47846
rect 47832 47844 47856 47846
rect 47912 47844 47918 47846
rect 47610 47835 47918 47844
rect 52610 47900 52918 47909
rect 52610 47898 52616 47900
rect 52672 47898 52696 47900
rect 52752 47898 52776 47900
rect 52832 47898 52856 47900
rect 52912 47898 52918 47900
rect 52672 47846 52674 47898
rect 52854 47846 52856 47898
rect 52610 47844 52616 47846
rect 52672 47844 52696 47846
rect 52752 47844 52776 47846
rect 52832 47844 52856 47846
rect 52912 47844 52918 47846
rect 52610 47835 52918 47844
rect 57610 47900 57918 47909
rect 57610 47898 57616 47900
rect 57672 47898 57696 47900
rect 57752 47898 57776 47900
rect 57832 47898 57856 47900
rect 57912 47898 57918 47900
rect 57672 47846 57674 47898
rect 57854 47846 57856 47898
rect 57610 47844 57616 47846
rect 57672 47844 57696 47846
rect 57752 47844 57776 47846
rect 57832 47844 57856 47846
rect 57912 47844 57918 47846
rect 57610 47835 57918 47844
rect 58532 47456 58584 47462
rect 58530 47424 58532 47433
rect 58584 47424 58586 47433
rect 1950 47356 2258 47365
rect 1950 47354 1956 47356
rect 2012 47354 2036 47356
rect 2092 47354 2116 47356
rect 2172 47354 2196 47356
rect 2252 47354 2258 47356
rect 2012 47302 2014 47354
rect 2194 47302 2196 47354
rect 1950 47300 1956 47302
rect 2012 47300 2036 47302
rect 2092 47300 2116 47302
rect 2172 47300 2196 47302
rect 2252 47300 2258 47302
rect 1950 47291 2258 47300
rect 6950 47356 7258 47365
rect 6950 47354 6956 47356
rect 7012 47354 7036 47356
rect 7092 47354 7116 47356
rect 7172 47354 7196 47356
rect 7252 47354 7258 47356
rect 7012 47302 7014 47354
rect 7194 47302 7196 47354
rect 6950 47300 6956 47302
rect 7012 47300 7036 47302
rect 7092 47300 7116 47302
rect 7172 47300 7196 47302
rect 7252 47300 7258 47302
rect 6950 47291 7258 47300
rect 11950 47356 12258 47365
rect 11950 47354 11956 47356
rect 12012 47354 12036 47356
rect 12092 47354 12116 47356
rect 12172 47354 12196 47356
rect 12252 47354 12258 47356
rect 12012 47302 12014 47354
rect 12194 47302 12196 47354
rect 11950 47300 11956 47302
rect 12012 47300 12036 47302
rect 12092 47300 12116 47302
rect 12172 47300 12196 47302
rect 12252 47300 12258 47302
rect 11950 47291 12258 47300
rect 16950 47356 17258 47365
rect 16950 47354 16956 47356
rect 17012 47354 17036 47356
rect 17092 47354 17116 47356
rect 17172 47354 17196 47356
rect 17252 47354 17258 47356
rect 17012 47302 17014 47354
rect 17194 47302 17196 47354
rect 16950 47300 16956 47302
rect 17012 47300 17036 47302
rect 17092 47300 17116 47302
rect 17172 47300 17196 47302
rect 17252 47300 17258 47302
rect 16950 47291 17258 47300
rect 21950 47356 22258 47365
rect 21950 47354 21956 47356
rect 22012 47354 22036 47356
rect 22092 47354 22116 47356
rect 22172 47354 22196 47356
rect 22252 47354 22258 47356
rect 22012 47302 22014 47354
rect 22194 47302 22196 47354
rect 21950 47300 21956 47302
rect 22012 47300 22036 47302
rect 22092 47300 22116 47302
rect 22172 47300 22196 47302
rect 22252 47300 22258 47302
rect 21950 47291 22258 47300
rect 26950 47356 27258 47365
rect 26950 47354 26956 47356
rect 27012 47354 27036 47356
rect 27092 47354 27116 47356
rect 27172 47354 27196 47356
rect 27252 47354 27258 47356
rect 27012 47302 27014 47354
rect 27194 47302 27196 47354
rect 26950 47300 26956 47302
rect 27012 47300 27036 47302
rect 27092 47300 27116 47302
rect 27172 47300 27196 47302
rect 27252 47300 27258 47302
rect 26950 47291 27258 47300
rect 31950 47356 32258 47365
rect 31950 47354 31956 47356
rect 32012 47354 32036 47356
rect 32092 47354 32116 47356
rect 32172 47354 32196 47356
rect 32252 47354 32258 47356
rect 32012 47302 32014 47354
rect 32194 47302 32196 47354
rect 31950 47300 31956 47302
rect 32012 47300 32036 47302
rect 32092 47300 32116 47302
rect 32172 47300 32196 47302
rect 32252 47300 32258 47302
rect 31950 47291 32258 47300
rect 36950 47356 37258 47365
rect 36950 47354 36956 47356
rect 37012 47354 37036 47356
rect 37092 47354 37116 47356
rect 37172 47354 37196 47356
rect 37252 47354 37258 47356
rect 37012 47302 37014 47354
rect 37194 47302 37196 47354
rect 36950 47300 36956 47302
rect 37012 47300 37036 47302
rect 37092 47300 37116 47302
rect 37172 47300 37196 47302
rect 37252 47300 37258 47302
rect 36950 47291 37258 47300
rect 41950 47356 42258 47365
rect 41950 47354 41956 47356
rect 42012 47354 42036 47356
rect 42092 47354 42116 47356
rect 42172 47354 42196 47356
rect 42252 47354 42258 47356
rect 42012 47302 42014 47354
rect 42194 47302 42196 47354
rect 41950 47300 41956 47302
rect 42012 47300 42036 47302
rect 42092 47300 42116 47302
rect 42172 47300 42196 47302
rect 42252 47300 42258 47302
rect 41950 47291 42258 47300
rect 46950 47356 47258 47365
rect 46950 47354 46956 47356
rect 47012 47354 47036 47356
rect 47092 47354 47116 47356
rect 47172 47354 47196 47356
rect 47252 47354 47258 47356
rect 47012 47302 47014 47354
rect 47194 47302 47196 47354
rect 46950 47300 46956 47302
rect 47012 47300 47036 47302
rect 47092 47300 47116 47302
rect 47172 47300 47196 47302
rect 47252 47300 47258 47302
rect 46950 47291 47258 47300
rect 51950 47356 52258 47365
rect 51950 47354 51956 47356
rect 52012 47354 52036 47356
rect 52092 47354 52116 47356
rect 52172 47354 52196 47356
rect 52252 47354 52258 47356
rect 52012 47302 52014 47354
rect 52194 47302 52196 47354
rect 51950 47300 51956 47302
rect 52012 47300 52036 47302
rect 52092 47300 52116 47302
rect 52172 47300 52196 47302
rect 52252 47300 52258 47302
rect 51950 47291 52258 47300
rect 56950 47356 57258 47365
rect 58530 47359 58586 47368
rect 56950 47354 56956 47356
rect 57012 47354 57036 47356
rect 57092 47354 57116 47356
rect 57172 47354 57196 47356
rect 57252 47354 57258 47356
rect 57012 47302 57014 47354
rect 57194 47302 57196 47354
rect 56950 47300 56956 47302
rect 57012 47300 57036 47302
rect 57092 47300 57116 47302
rect 57172 47300 57196 47302
rect 57252 47300 57258 47302
rect 56950 47291 57258 47300
rect 58532 47048 58584 47054
rect 58532 46990 58584 46996
rect 2610 46812 2918 46821
rect 2610 46810 2616 46812
rect 2672 46810 2696 46812
rect 2752 46810 2776 46812
rect 2832 46810 2856 46812
rect 2912 46810 2918 46812
rect 2672 46758 2674 46810
rect 2854 46758 2856 46810
rect 2610 46756 2616 46758
rect 2672 46756 2696 46758
rect 2752 46756 2776 46758
rect 2832 46756 2856 46758
rect 2912 46756 2918 46758
rect 2610 46747 2918 46756
rect 7610 46812 7918 46821
rect 7610 46810 7616 46812
rect 7672 46810 7696 46812
rect 7752 46810 7776 46812
rect 7832 46810 7856 46812
rect 7912 46810 7918 46812
rect 7672 46758 7674 46810
rect 7854 46758 7856 46810
rect 7610 46756 7616 46758
rect 7672 46756 7696 46758
rect 7752 46756 7776 46758
rect 7832 46756 7856 46758
rect 7912 46756 7918 46758
rect 7610 46747 7918 46756
rect 12610 46812 12918 46821
rect 12610 46810 12616 46812
rect 12672 46810 12696 46812
rect 12752 46810 12776 46812
rect 12832 46810 12856 46812
rect 12912 46810 12918 46812
rect 12672 46758 12674 46810
rect 12854 46758 12856 46810
rect 12610 46756 12616 46758
rect 12672 46756 12696 46758
rect 12752 46756 12776 46758
rect 12832 46756 12856 46758
rect 12912 46756 12918 46758
rect 12610 46747 12918 46756
rect 17610 46812 17918 46821
rect 17610 46810 17616 46812
rect 17672 46810 17696 46812
rect 17752 46810 17776 46812
rect 17832 46810 17856 46812
rect 17912 46810 17918 46812
rect 17672 46758 17674 46810
rect 17854 46758 17856 46810
rect 17610 46756 17616 46758
rect 17672 46756 17696 46758
rect 17752 46756 17776 46758
rect 17832 46756 17856 46758
rect 17912 46756 17918 46758
rect 17610 46747 17918 46756
rect 22610 46812 22918 46821
rect 22610 46810 22616 46812
rect 22672 46810 22696 46812
rect 22752 46810 22776 46812
rect 22832 46810 22856 46812
rect 22912 46810 22918 46812
rect 22672 46758 22674 46810
rect 22854 46758 22856 46810
rect 22610 46756 22616 46758
rect 22672 46756 22696 46758
rect 22752 46756 22776 46758
rect 22832 46756 22856 46758
rect 22912 46756 22918 46758
rect 22610 46747 22918 46756
rect 27610 46812 27918 46821
rect 27610 46810 27616 46812
rect 27672 46810 27696 46812
rect 27752 46810 27776 46812
rect 27832 46810 27856 46812
rect 27912 46810 27918 46812
rect 27672 46758 27674 46810
rect 27854 46758 27856 46810
rect 27610 46756 27616 46758
rect 27672 46756 27696 46758
rect 27752 46756 27776 46758
rect 27832 46756 27856 46758
rect 27912 46756 27918 46758
rect 27610 46747 27918 46756
rect 32610 46812 32918 46821
rect 32610 46810 32616 46812
rect 32672 46810 32696 46812
rect 32752 46810 32776 46812
rect 32832 46810 32856 46812
rect 32912 46810 32918 46812
rect 32672 46758 32674 46810
rect 32854 46758 32856 46810
rect 32610 46756 32616 46758
rect 32672 46756 32696 46758
rect 32752 46756 32776 46758
rect 32832 46756 32856 46758
rect 32912 46756 32918 46758
rect 32610 46747 32918 46756
rect 37610 46812 37918 46821
rect 37610 46810 37616 46812
rect 37672 46810 37696 46812
rect 37752 46810 37776 46812
rect 37832 46810 37856 46812
rect 37912 46810 37918 46812
rect 37672 46758 37674 46810
rect 37854 46758 37856 46810
rect 37610 46756 37616 46758
rect 37672 46756 37696 46758
rect 37752 46756 37776 46758
rect 37832 46756 37856 46758
rect 37912 46756 37918 46758
rect 37610 46747 37918 46756
rect 42610 46812 42918 46821
rect 42610 46810 42616 46812
rect 42672 46810 42696 46812
rect 42752 46810 42776 46812
rect 42832 46810 42856 46812
rect 42912 46810 42918 46812
rect 42672 46758 42674 46810
rect 42854 46758 42856 46810
rect 42610 46756 42616 46758
rect 42672 46756 42696 46758
rect 42752 46756 42776 46758
rect 42832 46756 42856 46758
rect 42912 46756 42918 46758
rect 42610 46747 42918 46756
rect 47610 46812 47918 46821
rect 47610 46810 47616 46812
rect 47672 46810 47696 46812
rect 47752 46810 47776 46812
rect 47832 46810 47856 46812
rect 47912 46810 47918 46812
rect 47672 46758 47674 46810
rect 47854 46758 47856 46810
rect 47610 46756 47616 46758
rect 47672 46756 47696 46758
rect 47752 46756 47776 46758
rect 47832 46756 47856 46758
rect 47912 46756 47918 46758
rect 47610 46747 47918 46756
rect 52610 46812 52918 46821
rect 52610 46810 52616 46812
rect 52672 46810 52696 46812
rect 52752 46810 52776 46812
rect 52832 46810 52856 46812
rect 52912 46810 52918 46812
rect 52672 46758 52674 46810
rect 52854 46758 52856 46810
rect 52610 46756 52616 46758
rect 52672 46756 52696 46758
rect 52752 46756 52776 46758
rect 52832 46756 52856 46758
rect 52912 46756 52918 46758
rect 52610 46747 52918 46756
rect 57610 46812 57918 46821
rect 57610 46810 57616 46812
rect 57672 46810 57696 46812
rect 57752 46810 57776 46812
rect 57832 46810 57856 46812
rect 57912 46810 57918 46812
rect 57672 46758 57674 46810
rect 57854 46758 57856 46810
rect 57610 46756 57616 46758
rect 57672 46756 57696 46758
rect 57752 46756 57776 46758
rect 57832 46756 57856 46758
rect 57912 46756 57918 46758
rect 57610 46747 57918 46756
rect 58544 46617 58572 46990
rect 58530 46608 58586 46617
rect 58530 46543 58586 46552
rect 1950 46268 2258 46277
rect 1950 46266 1956 46268
rect 2012 46266 2036 46268
rect 2092 46266 2116 46268
rect 2172 46266 2196 46268
rect 2252 46266 2258 46268
rect 2012 46214 2014 46266
rect 2194 46214 2196 46266
rect 1950 46212 1956 46214
rect 2012 46212 2036 46214
rect 2092 46212 2116 46214
rect 2172 46212 2196 46214
rect 2252 46212 2258 46214
rect 1950 46203 2258 46212
rect 6950 46268 7258 46277
rect 6950 46266 6956 46268
rect 7012 46266 7036 46268
rect 7092 46266 7116 46268
rect 7172 46266 7196 46268
rect 7252 46266 7258 46268
rect 7012 46214 7014 46266
rect 7194 46214 7196 46266
rect 6950 46212 6956 46214
rect 7012 46212 7036 46214
rect 7092 46212 7116 46214
rect 7172 46212 7196 46214
rect 7252 46212 7258 46214
rect 6950 46203 7258 46212
rect 11950 46268 12258 46277
rect 11950 46266 11956 46268
rect 12012 46266 12036 46268
rect 12092 46266 12116 46268
rect 12172 46266 12196 46268
rect 12252 46266 12258 46268
rect 12012 46214 12014 46266
rect 12194 46214 12196 46266
rect 11950 46212 11956 46214
rect 12012 46212 12036 46214
rect 12092 46212 12116 46214
rect 12172 46212 12196 46214
rect 12252 46212 12258 46214
rect 11950 46203 12258 46212
rect 16950 46268 17258 46277
rect 16950 46266 16956 46268
rect 17012 46266 17036 46268
rect 17092 46266 17116 46268
rect 17172 46266 17196 46268
rect 17252 46266 17258 46268
rect 17012 46214 17014 46266
rect 17194 46214 17196 46266
rect 16950 46212 16956 46214
rect 17012 46212 17036 46214
rect 17092 46212 17116 46214
rect 17172 46212 17196 46214
rect 17252 46212 17258 46214
rect 16950 46203 17258 46212
rect 21950 46268 22258 46277
rect 21950 46266 21956 46268
rect 22012 46266 22036 46268
rect 22092 46266 22116 46268
rect 22172 46266 22196 46268
rect 22252 46266 22258 46268
rect 22012 46214 22014 46266
rect 22194 46214 22196 46266
rect 21950 46212 21956 46214
rect 22012 46212 22036 46214
rect 22092 46212 22116 46214
rect 22172 46212 22196 46214
rect 22252 46212 22258 46214
rect 21950 46203 22258 46212
rect 26950 46268 27258 46277
rect 26950 46266 26956 46268
rect 27012 46266 27036 46268
rect 27092 46266 27116 46268
rect 27172 46266 27196 46268
rect 27252 46266 27258 46268
rect 27012 46214 27014 46266
rect 27194 46214 27196 46266
rect 26950 46212 26956 46214
rect 27012 46212 27036 46214
rect 27092 46212 27116 46214
rect 27172 46212 27196 46214
rect 27252 46212 27258 46214
rect 26950 46203 27258 46212
rect 31950 46268 32258 46277
rect 31950 46266 31956 46268
rect 32012 46266 32036 46268
rect 32092 46266 32116 46268
rect 32172 46266 32196 46268
rect 32252 46266 32258 46268
rect 32012 46214 32014 46266
rect 32194 46214 32196 46266
rect 31950 46212 31956 46214
rect 32012 46212 32036 46214
rect 32092 46212 32116 46214
rect 32172 46212 32196 46214
rect 32252 46212 32258 46214
rect 31950 46203 32258 46212
rect 36950 46268 37258 46277
rect 36950 46266 36956 46268
rect 37012 46266 37036 46268
rect 37092 46266 37116 46268
rect 37172 46266 37196 46268
rect 37252 46266 37258 46268
rect 37012 46214 37014 46266
rect 37194 46214 37196 46266
rect 36950 46212 36956 46214
rect 37012 46212 37036 46214
rect 37092 46212 37116 46214
rect 37172 46212 37196 46214
rect 37252 46212 37258 46214
rect 36950 46203 37258 46212
rect 41950 46268 42258 46277
rect 41950 46266 41956 46268
rect 42012 46266 42036 46268
rect 42092 46266 42116 46268
rect 42172 46266 42196 46268
rect 42252 46266 42258 46268
rect 42012 46214 42014 46266
rect 42194 46214 42196 46266
rect 41950 46212 41956 46214
rect 42012 46212 42036 46214
rect 42092 46212 42116 46214
rect 42172 46212 42196 46214
rect 42252 46212 42258 46214
rect 41950 46203 42258 46212
rect 46950 46268 47258 46277
rect 46950 46266 46956 46268
rect 47012 46266 47036 46268
rect 47092 46266 47116 46268
rect 47172 46266 47196 46268
rect 47252 46266 47258 46268
rect 47012 46214 47014 46266
rect 47194 46214 47196 46266
rect 46950 46212 46956 46214
rect 47012 46212 47036 46214
rect 47092 46212 47116 46214
rect 47172 46212 47196 46214
rect 47252 46212 47258 46214
rect 46950 46203 47258 46212
rect 51950 46268 52258 46277
rect 51950 46266 51956 46268
rect 52012 46266 52036 46268
rect 52092 46266 52116 46268
rect 52172 46266 52196 46268
rect 52252 46266 52258 46268
rect 52012 46214 52014 46266
rect 52194 46214 52196 46266
rect 51950 46212 51956 46214
rect 52012 46212 52036 46214
rect 52092 46212 52116 46214
rect 52172 46212 52196 46214
rect 52252 46212 52258 46214
rect 51950 46203 52258 46212
rect 56950 46268 57258 46277
rect 56950 46266 56956 46268
rect 57012 46266 57036 46268
rect 57092 46266 57116 46268
rect 57172 46266 57196 46268
rect 57252 46266 57258 46268
rect 57012 46214 57014 46266
rect 57194 46214 57196 46266
rect 56950 46212 56956 46214
rect 57012 46212 57036 46214
rect 57092 46212 57116 46214
rect 57172 46212 57196 46214
rect 57252 46212 57258 46214
rect 56950 46203 57258 46212
rect 58532 45960 58584 45966
rect 58532 45902 58584 45908
rect 58544 45801 58572 45902
rect 58530 45792 58586 45801
rect 2610 45724 2918 45733
rect 2610 45722 2616 45724
rect 2672 45722 2696 45724
rect 2752 45722 2776 45724
rect 2832 45722 2856 45724
rect 2912 45722 2918 45724
rect 2672 45670 2674 45722
rect 2854 45670 2856 45722
rect 2610 45668 2616 45670
rect 2672 45668 2696 45670
rect 2752 45668 2776 45670
rect 2832 45668 2856 45670
rect 2912 45668 2918 45670
rect 2610 45659 2918 45668
rect 7610 45724 7918 45733
rect 7610 45722 7616 45724
rect 7672 45722 7696 45724
rect 7752 45722 7776 45724
rect 7832 45722 7856 45724
rect 7912 45722 7918 45724
rect 7672 45670 7674 45722
rect 7854 45670 7856 45722
rect 7610 45668 7616 45670
rect 7672 45668 7696 45670
rect 7752 45668 7776 45670
rect 7832 45668 7856 45670
rect 7912 45668 7918 45670
rect 7610 45659 7918 45668
rect 12610 45724 12918 45733
rect 12610 45722 12616 45724
rect 12672 45722 12696 45724
rect 12752 45722 12776 45724
rect 12832 45722 12856 45724
rect 12912 45722 12918 45724
rect 12672 45670 12674 45722
rect 12854 45670 12856 45722
rect 12610 45668 12616 45670
rect 12672 45668 12696 45670
rect 12752 45668 12776 45670
rect 12832 45668 12856 45670
rect 12912 45668 12918 45670
rect 12610 45659 12918 45668
rect 17610 45724 17918 45733
rect 17610 45722 17616 45724
rect 17672 45722 17696 45724
rect 17752 45722 17776 45724
rect 17832 45722 17856 45724
rect 17912 45722 17918 45724
rect 17672 45670 17674 45722
rect 17854 45670 17856 45722
rect 17610 45668 17616 45670
rect 17672 45668 17696 45670
rect 17752 45668 17776 45670
rect 17832 45668 17856 45670
rect 17912 45668 17918 45670
rect 17610 45659 17918 45668
rect 22610 45724 22918 45733
rect 22610 45722 22616 45724
rect 22672 45722 22696 45724
rect 22752 45722 22776 45724
rect 22832 45722 22856 45724
rect 22912 45722 22918 45724
rect 22672 45670 22674 45722
rect 22854 45670 22856 45722
rect 22610 45668 22616 45670
rect 22672 45668 22696 45670
rect 22752 45668 22776 45670
rect 22832 45668 22856 45670
rect 22912 45668 22918 45670
rect 22610 45659 22918 45668
rect 27610 45724 27918 45733
rect 27610 45722 27616 45724
rect 27672 45722 27696 45724
rect 27752 45722 27776 45724
rect 27832 45722 27856 45724
rect 27912 45722 27918 45724
rect 27672 45670 27674 45722
rect 27854 45670 27856 45722
rect 27610 45668 27616 45670
rect 27672 45668 27696 45670
rect 27752 45668 27776 45670
rect 27832 45668 27856 45670
rect 27912 45668 27918 45670
rect 27610 45659 27918 45668
rect 32610 45724 32918 45733
rect 32610 45722 32616 45724
rect 32672 45722 32696 45724
rect 32752 45722 32776 45724
rect 32832 45722 32856 45724
rect 32912 45722 32918 45724
rect 32672 45670 32674 45722
rect 32854 45670 32856 45722
rect 32610 45668 32616 45670
rect 32672 45668 32696 45670
rect 32752 45668 32776 45670
rect 32832 45668 32856 45670
rect 32912 45668 32918 45670
rect 32610 45659 32918 45668
rect 37610 45724 37918 45733
rect 37610 45722 37616 45724
rect 37672 45722 37696 45724
rect 37752 45722 37776 45724
rect 37832 45722 37856 45724
rect 37912 45722 37918 45724
rect 37672 45670 37674 45722
rect 37854 45670 37856 45722
rect 37610 45668 37616 45670
rect 37672 45668 37696 45670
rect 37752 45668 37776 45670
rect 37832 45668 37856 45670
rect 37912 45668 37918 45670
rect 37610 45659 37918 45668
rect 42610 45724 42918 45733
rect 42610 45722 42616 45724
rect 42672 45722 42696 45724
rect 42752 45722 42776 45724
rect 42832 45722 42856 45724
rect 42912 45722 42918 45724
rect 42672 45670 42674 45722
rect 42854 45670 42856 45722
rect 42610 45668 42616 45670
rect 42672 45668 42696 45670
rect 42752 45668 42776 45670
rect 42832 45668 42856 45670
rect 42912 45668 42918 45670
rect 42610 45659 42918 45668
rect 47610 45724 47918 45733
rect 47610 45722 47616 45724
rect 47672 45722 47696 45724
rect 47752 45722 47776 45724
rect 47832 45722 47856 45724
rect 47912 45722 47918 45724
rect 47672 45670 47674 45722
rect 47854 45670 47856 45722
rect 47610 45668 47616 45670
rect 47672 45668 47696 45670
rect 47752 45668 47776 45670
rect 47832 45668 47856 45670
rect 47912 45668 47918 45670
rect 47610 45659 47918 45668
rect 52610 45724 52918 45733
rect 52610 45722 52616 45724
rect 52672 45722 52696 45724
rect 52752 45722 52776 45724
rect 52832 45722 52856 45724
rect 52912 45722 52918 45724
rect 52672 45670 52674 45722
rect 52854 45670 52856 45722
rect 52610 45668 52616 45670
rect 52672 45668 52696 45670
rect 52752 45668 52776 45670
rect 52832 45668 52856 45670
rect 52912 45668 52918 45670
rect 52610 45659 52918 45668
rect 57610 45724 57918 45733
rect 58530 45727 58586 45736
rect 57610 45722 57616 45724
rect 57672 45722 57696 45724
rect 57752 45722 57776 45724
rect 57832 45722 57856 45724
rect 57912 45722 57918 45724
rect 57672 45670 57674 45722
rect 57854 45670 57856 45722
rect 57610 45668 57616 45670
rect 57672 45668 57696 45670
rect 57752 45668 57776 45670
rect 57832 45668 57856 45670
rect 57912 45668 57918 45670
rect 57610 45659 57918 45668
rect 58532 45280 58584 45286
rect 58532 45222 58584 45228
rect 1950 45180 2258 45189
rect 1950 45178 1956 45180
rect 2012 45178 2036 45180
rect 2092 45178 2116 45180
rect 2172 45178 2196 45180
rect 2252 45178 2258 45180
rect 2012 45126 2014 45178
rect 2194 45126 2196 45178
rect 1950 45124 1956 45126
rect 2012 45124 2036 45126
rect 2092 45124 2116 45126
rect 2172 45124 2196 45126
rect 2252 45124 2258 45126
rect 1950 45115 2258 45124
rect 6950 45180 7258 45189
rect 6950 45178 6956 45180
rect 7012 45178 7036 45180
rect 7092 45178 7116 45180
rect 7172 45178 7196 45180
rect 7252 45178 7258 45180
rect 7012 45126 7014 45178
rect 7194 45126 7196 45178
rect 6950 45124 6956 45126
rect 7012 45124 7036 45126
rect 7092 45124 7116 45126
rect 7172 45124 7196 45126
rect 7252 45124 7258 45126
rect 6950 45115 7258 45124
rect 11950 45180 12258 45189
rect 11950 45178 11956 45180
rect 12012 45178 12036 45180
rect 12092 45178 12116 45180
rect 12172 45178 12196 45180
rect 12252 45178 12258 45180
rect 12012 45126 12014 45178
rect 12194 45126 12196 45178
rect 11950 45124 11956 45126
rect 12012 45124 12036 45126
rect 12092 45124 12116 45126
rect 12172 45124 12196 45126
rect 12252 45124 12258 45126
rect 11950 45115 12258 45124
rect 16950 45180 17258 45189
rect 16950 45178 16956 45180
rect 17012 45178 17036 45180
rect 17092 45178 17116 45180
rect 17172 45178 17196 45180
rect 17252 45178 17258 45180
rect 17012 45126 17014 45178
rect 17194 45126 17196 45178
rect 16950 45124 16956 45126
rect 17012 45124 17036 45126
rect 17092 45124 17116 45126
rect 17172 45124 17196 45126
rect 17252 45124 17258 45126
rect 16950 45115 17258 45124
rect 21950 45180 22258 45189
rect 21950 45178 21956 45180
rect 22012 45178 22036 45180
rect 22092 45178 22116 45180
rect 22172 45178 22196 45180
rect 22252 45178 22258 45180
rect 22012 45126 22014 45178
rect 22194 45126 22196 45178
rect 21950 45124 21956 45126
rect 22012 45124 22036 45126
rect 22092 45124 22116 45126
rect 22172 45124 22196 45126
rect 22252 45124 22258 45126
rect 21950 45115 22258 45124
rect 26950 45180 27258 45189
rect 26950 45178 26956 45180
rect 27012 45178 27036 45180
rect 27092 45178 27116 45180
rect 27172 45178 27196 45180
rect 27252 45178 27258 45180
rect 27012 45126 27014 45178
rect 27194 45126 27196 45178
rect 26950 45124 26956 45126
rect 27012 45124 27036 45126
rect 27092 45124 27116 45126
rect 27172 45124 27196 45126
rect 27252 45124 27258 45126
rect 26950 45115 27258 45124
rect 31950 45180 32258 45189
rect 31950 45178 31956 45180
rect 32012 45178 32036 45180
rect 32092 45178 32116 45180
rect 32172 45178 32196 45180
rect 32252 45178 32258 45180
rect 32012 45126 32014 45178
rect 32194 45126 32196 45178
rect 31950 45124 31956 45126
rect 32012 45124 32036 45126
rect 32092 45124 32116 45126
rect 32172 45124 32196 45126
rect 32252 45124 32258 45126
rect 31950 45115 32258 45124
rect 36950 45180 37258 45189
rect 36950 45178 36956 45180
rect 37012 45178 37036 45180
rect 37092 45178 37116 45180
rect 37172 45178 37196 45180
rect 37252 45178 37258 45180
rect 37012 45126 37014 45178
rect 37194 45126 37196 45178
rect 36950 45124 36956 45126
rect 37012 45124 37036 45126
rect 37092 45124 37116 45126
rect 37172 45124 37196 45126
rect 37252 45124 37258 45126
rect 36950 45115 37258 45124
rect 41950 45180 42258 45189
rect 41950 45178 41956 45180
rect 42012 45178 42036 45180
rect 42092 45178 42116 45180
rect 42172 45178 42196 45180
rect 42252 45178 42258 45180
rect 42012 45126 42014 45178
rect 42194 45126 42196 45178
rect 41950 45124 41956 45126
rect 42012 45124 42036 45126
rect 42092 45124 42116 45126
rect 42172 45124 42196 45126
rect 42252 45124 42258 45126
rect 41950 45115 42258 45124
rect 46950 45180 47258 45189
rect 46950 45178 46956 45180
rect 47012 45178 47036 45180
rect 47092 45178 47116 45180
rect 47172 45178 47196 45180
rect 47252 45178 47258 45180
rect 47012 45126 47014 45178
rect 47194 45126 47196 45178
rect 46950 45124 46956 45126
rect 47012 45124 47036 45126
rect 47092 45124 47116 45126
rect 47172 45124 47196 45126
rect 47252 45124 47258 45126
rect 46950 45115 47258 45124
rect 51950 45180 52258 45189
rect 51950 45178 51956 45180
rect 52012 45178 52036 45180
rect 52092 45178 52116 45180
rect 52172 45178 52196 45180
rect 52252 45178 52258 45180
rect 52012 45126 52014 45178
rect 52194 45126 52196 45178
rect 51950 45124 51956 45126
rect 52012 45124 52036 45126
rect 52092 45124 52116 45126
rect 52172 45124 52196 45126
rect 52252 45124 52258 45126
rect 51950 45115 52258 45124
rect 56950 45180 57258 45189
rect 56950 45178 56956 45180
rect 57012 45178 57036 45180
rect 57092 45178 57116 45180
rect 57172 45178 57196 45180
rect 57252 45178 57258 45180
rect 57012 45126 57014 45178
rect 57194 45126 57196 45178
rect 56950 45124 56956 45126
rect 57012 45124 57036 45126
rect 57092 45124 57116 45126
rect 57172 45124 57196 45126
rect 57252 45124 57258 45126
rect 56950 45115 57258 45124
rect 58544 44985 58572 45222
rect 58530 44976 58586 44985
rect 58530 44911 58586 44920
rect 2610 44636 2918 44645
rect 2610 44634 2616 44636
rect 2672 44634 2696 44636
rect 2752 44634 2776 44636
rect 2832 44634 2856 44636
rect 2912 44634 2918 44636
rect 2672 44582 2674 44634
rect 2854 44582 2856 44634
rect 2610 44580 2616 44582
rect 2672 44580 2696 44582
rect 2752 44580 2776 44582
rect 2832 44580 2856 44582
rect 2912 44580 2918 44582
rect 2610 44571 2918 44580
rect 7610 44636 7918 44645
rect 7610 44634 7616 44636
rect 7672 44634 7696 44636
rect 7752 44634 7776 44636
rect 7832 44634 7856 44636
rect 7912 44634 7918 44636
rect 7672 44582 7674 44634
rect 7854 44582 7856 44634
rect 7610 44580 7616 44582
rect 7672 44580 7696 44582
rect 7752 44580 7776 44582
rect 7832 44580 7856 44582
rect 7912 44580 7918 44582
rect 7610 44571 7918 44580
rect 12610 44636 12918 44645
rect 12610 44634 12616 44636
rect 12672 44634 12696 44636
rect 12752 44634 12776 44636
rect 12832 44634 12856 44636
rect 12912 44634 12918 44636
rect 12672 44582 12674 44634
rect 12854 44582 12856 44634
rect 12610 44580 12616 44582
rect 12672 44580 12696 44582
rect 12752 44580 12776 44582
rect 12832 44580 12856 44582
rect 12912 44580 12918 44582
rect 12610 44571 12918 44580
rect 17610 44636 17918 44645
rect 17610 44634 17616 44636
rect 17672 44634 17696 44636
rect 17752 44634 17776 44636
rect 17832 44634 17856 44636
rect 17912 44634 17918 44636
rect 17672 44582 17674 44634
rect 17854 44582 17856 44634
rect 17610 44580 17616 44582
rect 17672 44580 17696 44582
rect 17752 44580 17776 44582
rect 17832 44580 17856 44582
rect 17912 44580 17918 44582
rect 17610 44571 17918 44580
rect 22610 44636 22918 44645
rect 22610 44634 22616 44636
rect 22672 44634 22696 44636
rect 22752 44634 22776 44636
rect 22832 44634 22856 44636
rect 22912 44634 22918 44636
rect 22672 44582 22674 44634
rect 22854 44582 22856 44634
rect 22610 44580 22616 44582
rect 22672 44580 22696 44582
rect 22752 44580 22776 44582
rect 22832 44580 22856 44582
rect 22912 44580 22918 44582
rect 22610 44571 22918 44580
rect 27610 44636 27918 44645
rect 27610 44634 27616 44636
rect 27672 44634 27696 44636
rect 27752 44634 27776 44636
rect 27832 44634 27856 44636
rect 27912 44634 27918 44636
rect 27672 44582 27674 44634
rect 27854 44582 27856 44634
rect 27610 44580 27616 44582
rect 27672 44580 27696 44582
rect 27752 44580 27776 44582
rect 27832 44580 27856 44582
rect 27912 44580 27918 44582
rect 27610 44571 27918 44580
rect 32610 44636 32918 44645
rect 32610 44634 32616 44636
rect 32672 44634 32696 44636
rect 32752 44634 32776 44636
rect 32832 44634 32856 44636
rect 32912 44634 32918 44636
rect 32672 44582 32674 44634
rect 32854 44582 32856 44634
rect 32610 44580 32616 44582
rect 32672 44580 32696 44582
rect 32752 44580 32776 44582
rect 32832 44580 32856 44582
rect 32912 44580 32918 44582
rect 32610 44571 32918 44580
rect 37610 44636 37918 44645
rect 37610 44634 37616 44636
rect 37672 44634 37696 44636
rect 37752 44634 37776 44636
rect 37832 44634 37856 44636
rect 37912 44634 37918 44636
rect 37672 44582 37674 44634
rect 37854 44582 37856 44634
rect 37610 44580 37616 44582
rect 37672 44580 37696 44582
rect 37752 44580 37776 44582
rect 37832 44580 37856 44582
rect 37912 44580 37918 44582
rect 37610 44571 37918 44580
rect 42610 44636 42918 44645
rect 42610 44634 42616 44636
rect 42672 44634 42696 44636
rect 42752 44634 42776 44636
rect 42832 44634 42856 44636
rect 42912 44634 42918 44636
rect 42672 44582 42674 44634
rect 42854 44582 42856 44634
rect 42610 44580 42616 44582
rect 42672 44580 42696 44582
rect 42752 44580 42776 44582
rect 42832 44580 42856 44582
rect 42912 44580 42918 44582
rect 42610 44571 42918 44580
rect 47610 44636 47918 44645
rect 47610 44634 47616 44636
rect 47672 44634 47696 44636
rect 47752 44634 47776 44636
rect 47832 44634 47856 44636
rect 47912 44634 47918 44636
rect 47672 44582 47674 44634
rect 47854 44582 47856 44634
rect 47610 44580 47616 44582
rect 47672 44580 47696 44582
rect 47752 44580 47776 44582
rect 47832 44580 47856 44582
rect 47912 44580 47918 44582
rect 47610 44571 47918 44580
rect 52610 44636 52918 44645
rect 52610 44634 52616 44636
rect 52672 44634 52696 44636
rect 52752 44634 52776 44636
rect 52832 44634 52856 44636
rect 52912 44634 52918 44636
rect 52672 44582 52674 44634
rect 52854 44582 52856 44634
rect 52610 44580 52616 44582
rect 52672 44580 52696 44582
rect 52752 44580 52776 44582
rect 52832 44580 52856 44582
rect 52912 44580 52918 44582
rect 52610 44571 52918 44580
rect 57610 44636 57918 44645
rect 57610 44634 57616 44636
rect 57672 44634 57696 44636
rect 57752 44634 57776 44636
rect 57832 44634 57856 44636
rect 57912 44634 57918 44636
rect 57672 44582 57674 44634
rect 57854 44582 57856 44634
rect 57610 44580 57616 44582
rect 57672 44580 57696 44582
rect 57752 44580 57776 44582
rect 57832 44580 57856 44582
rect 57912 44580 57918 44582
rect 57610 44571 57918 44580
rect 58532 44192 58584 44198
rect 58530 44160 58532 44169
rect 58584 44160 58586 44169
rect 1950 44092 2258 44101
rect 1950 44090 1956 44092
rect 2012 44090 2036 44092
rect 2092 44090 2116 44092
rect 2172 44090 2196 44092
rect 2252 44090 2258 44092
rect 2012 44038 2014 44090
rect 2194 44038 2196 44090
rect 1950 44036 1956 44038
rect 2012 44036 2036 44038
rect 2092 44036 2116 44038
rect 2172 44036 2196 44038
rect 2252 44036 2258 44038
rect 1950 44027 2258 44036
rect 6950 44092 7258 44101
rect 6950 44090 6956 44092
rect 7012 44090 7036 44092
rect 7092 44090 7116 44092
rect 7172 44090 7196 44092
rect 7252 44090 7258 44092
rect 7012 44038 7014 44090
rect 7194 44038 7196 44090
rect 6950 44036 6956 44038
rect 7012 44036 7036 44038
rect 7092 44036 7116 44038
rect 7172 44036 7196 44038
rect 7252 44036 7258 44038
rect 6950 44027 7258 44036
rect 11950 44092 12258 44101
rect 11950 44090 11956 44092
rect 12012 44090 12036 44092
rect 12092 44090 12116 44092
rect 12172 44090 12196 44092
rect 12252 44090 12258 44092
rect 12012 44038 12014 44090
rect 12194 44038 12196 44090
rect 11950 44036 11956 44038
rect 12012 44036 12036 44038
rect 12092 44036 12116 44038
rect 12172 44036 12196 44038
rect 12252 44036 12258 44038
rect 11950 44027 12258 44036
rect 16950 44092 17258 44101
rect 16950 44090 16956 44092
rect 17012 44090 17036 44092
rect 17092 44090 17116 44092
rect 17172 44090 17196 44092
rect 17252 44090 17258 44092
rect 17012 44038 17014 44090
rect 17194 44038 17196 44090
rect 16950 44036 16956 44038
rect 17012 44036 17036 44038
rect 17092 44036 17116 44038
rect 17172 44036 17196 44038
rect 17252 44036 17258 44038
rect 16950 44027 17258 44036
rect 21950 44092 22258 44101
rect 21950 44090 21956 44092
rect 22012 44090 22036 44092
rect 22092 44090 22116 44092
rect 22172 44090 22196 44092
rect 22252 44090 22258 44092
rect 22012 44038 22014 44090
rect 22194 44038 22196 44090
rect 21950 44036 21956 44038
rect 22012 44036 22036 44038
rect 22092 44036 22116 44038
rect 22172 44036 22196 44038
rect 22252 44036 22258 44038
rect 21950 44027 22258 44036
rect 26950 44092 27258 44101
rect 26950 44090 26956 44092
rect 27012 44090 27036 44092
rect 27092 44090 27116 44092
rect 27172 44090 27196 44092
rect 27252 44090 27258 44092
rect 27012 44038 27014 44090
rect 27194 44038 27196 44090
rect 26950 44036 26956 44038
rect 27012 44036 27036 44038
rect 27092 44036 27116 44038
rect 27172 44036 27196 44038
rect 27252 44036 27258 44038
rect 26950 44027 27258 44036
rect 31950 44092 32258 44101
rect 31950 44090 31956 44092
rect 32012 44090 32036 44092
rect 32092 44090 32116 44092
rect 32172 44090 32196 44092
rect 32252 44090 32258 44092
rect 32012 44038 32014 44090
rect 32194 44038 32196 44090
rect 31950 44036 31956 44038
rect 32012 44036 32036 44038
rect 32092 44036 32116 44038
rect 32172 44036 32196 44038
rect 32252 44036 32258 44038
rect 31950 44027 32258 44036
rect 36950 44092 37258 44101
rect 36950 44090 36956 44092
rect 37012 44090 37036 44092
rect 37092 44090 37116 44092
rect 37172 44090 37196 44092
rect 37252 44090 37258 44092
rect 37012 44038 37014 44090
rect 37194 44038 37196 44090
rect 36950 44036 36956 44038
rect 37012 44036 37036 44038
rect 37092 44036 37116 44038
rect 37172 44036 37196 44038
rect 37252 44036 37258 44038
rect 36950 44027 37258 44036
rect 41950 44092 42258 44101
rect 41950 44090 41956 44092
rect 42012 44090 42036 44092
rect 42092 44090 42116 44092
rect 42172 44090 42196 44092
rect 42252 44090 42258 44092
rect 42012 44038 42014 44090
rect 42194 44038 42196 44090
rect 41950 44036 41956 44038
rect 42012 44036 42036 44038
rect 42092 44036 42116 44038
rect 42172 44036 42196 44038
rect 42252 44036 42258 44038
rect 41950 44027 42258 44036
rect 46950 44092 47258 44101
rect 46950 44090 46956 44092
rect 47012 44090 47036 44092
rect 47092 44090 47116 44092
rect 47172 44090 47196 44092
rect 47252 44090 47258 44092
rect 47012 44038 47014 44090
rect 47194 44038 47196 44090
rect 46950 44036 46956 44038
rect 47012 44036 47036 44038
rect 47092 44036 47116 44038
rect 47172 44036 47196 44038
rect 47252 44036 47258 44038
rect 46950 44027 47258 44036
rect 51950 44092 52258 44101
rect 51950 44090 51956 44092
rect 52012 44090 52036 44092
rect 52092 44090 52116 44092
rect 52172 44090 52196 44092
rect 52252 44090 52258 44092
rect 52012 44038 52014 44090
rect 52194 44038 52196 44090
rect 51950 44036 51956 44038
rect 52012 44036 52036 44038
rect 52092 44036 52116 44038
rect 52172 44036 52196 44038
rect 52252 44036 52258 44038
rect 51950 44027 52258 44036
rect 56950 44092 57258 44101
rect 58530 44095 58586 44104
rect 56950 44090 56956 44092
rect 57012 44090 57036 44092
rect 57092 44090 57116 44092
rect 57172 44090 57196 44092
rect 57252 44090 57258 44092
rect 57012 44038 57014 44090
rect 57194 44038 57196 44090
rect 56950 44036 56956 44038
rect 57012 44036 57036 44038
rect 57092 44036 57116 44038
rect 57172 44036 57196 44038
rect 57252 44036 57258 44038
rect 56950 44027 57258 44036
rect 58532 43784 58584 43790
rect 58532 43726 58584 43732
rect 2610 43548 2918 43557
rect 2610 43546 2616 43548
rect 2672 43546 2696 43548
rect 2752 43546 2776 43548
rect 2832 43546 2856 43548
rect 2912 43546 2918 43548
rect 2672 43494 2674 43546
rect 2854 43494 2856 43546
rect 2610 43492 2616 43494
rect 2672 43492 2696 43494
rect 2752 43492 2776 43494
rect 2832 43492 2856 43494
rect 2912 43492 2918 43494
rect 2610 43483 2918 43492
rect 7610 43548 7918 43557
rect 7610 43546 7616 43548
rect 7672 43546 7696 43548
rect 7752 43546 7776 43548
rect 7832 43546 7856 43548
rect 7912 43546 7918 43548
rect 7672 43494 7674 43546
rect 7854 43494 7856 43546
rect 7610 43492 7616 43494
rect 7672 43492 7696 43494
rect 7752 43492 7776 43494
rect 7832 43492 7856 43494
rect 7912 43492 7918 43494
rect 7610 43483 7918 43492
rect 12610 43548 12918 43557
rect 12610 43546 12616 43548
rect 12672 43546 12696 43548
rect 12752 43546 12776 43548
rect 12832 43546 12856 43548
rect 12912 43546 12918 43548
rect 12672 43494 12674 43546
rect 12854 43494 12856 43546
rect 12610 43492 12616 43494
rect 12672 43492 12696 43494
rect 12752 43492 12776 43494
rect 12832 43492 12856 43494
rect 12912 43492 12918 43494
rect 12610 43483 12918 43492
rect 17610 43548 17918 43557
rect 17610 43546 17616 43548
rect 17672 43546 17696 43548
rect 17752 43546 17776 43548
rect 17832 43546 17856 43548
rect 17912 43546 17918 43548
rect 17672 43494 17674 43546
rect 17854 43494 17856 43546
rect 17610 43492 17616 43494
rect 17672 43492 17696 43494
rect 17752 43492 17776 43494
rect 17832 43492 17856 43494
rect 17912 43492 17918 43494
rect 17610 43483 17918 43492
rect 22610 43548 22918 43557
rect 22610 43546 22616 43548
rect 22672 43546 22696 43548
rect 22752 43546 22776 43548
rect 22832 43546 22856 43548
rect 22912 43546 22918 43548
rect 22672 43494 22674 43546
rect 22854 43494 22856 43546
rect 22610 43492 22616 43494
rect 22672 43492 22696 43494
rect 22752 43492 22776 43494
rect 22832 43492 22856 43494
rect 22912 43492 22918 43494
rect 22610 43483 22918 43492
rect 27610 43548 27918 43557
rect 27610 43546 27616 43548
rect 27672 43546 27696 43548
rect 27752 43546 27776 43548
rect 27832 43546 27856 43548
rect 27912 43546 27918 43548
rect 27672 43494 27674 43546
rect 27854 43494 27856 43546
rect 27610 43492 27616 43494
rect 27672 43492 27696 43494
rect 27752 43492 27776 43494
rect 27832 43492 27856 43494
rect 27912 43492 27918 43494
rect 27610 43483 27918 43492
rect 32610 43548 32918 43557
rect 32610 43546 32616 43548
rect 32672 43546 32696 43548
rect 32752 43546 32776 43548
rect 32832 43546 32856 43548
rect 32912 43546 32918 43548
rect 32672 43494 32674 43546
rect 32854 43494 32856 43546
rect 32610 43492 32616 43494
rect 32672 43492 32696 43494
rect 32752 43492 32776 43494
rect 32832 43492 32856 43494
rect 32912 43492 32918 43494
rect 32610 43483 32918 43492
rect 37610 43548 37918 43557
rect 37610 43546 37616 43548
rect 37672 43546 37696 43548
rect 37752 43546 37776 43548
rect 37832 43546 37856 43548
rect 37912 43546 37918 43548
rect 37672 43494 37674 43546
rect 37854 43494 37856 43546
rect 37610 43492 37616 43494
rect 37672 43492 37696 43494
rect 37752 43492 37776 43494
rect 37832 43492 37856 43494
rect 37912 43492 37918 43494
rect 37610 43483 37918 43492
rect 42610 43548 42918 43557
rect 42610 43546 42616 43548
rect 42672 43546 42696 43548
rect 42752 43546 42776 43548
rect 42832 43546 42856 43548
rect 42912 43546 42918 43548
rect 42672 43494 42674 43546
rect 42854 43494 42856 43546
rect 42610 43492 42616 43494
rect 42672 43492 42696 43494
rect 42752 43492 42776 43494
rect 42832 43492 42856 43494
rect 42912 43492 42918 43494
rect 42610 43483 42918 43492
rect 47610 43548 47918 43557
rect 47610 43546 47616 43548
rect 47672 43546 47696 43548
rect 47752 43546 47776 43548
rect 47832 43546 47856 43548
rect 47912 43546 47918 43548
rect 47672 43494 47674 43546
rect 47854 43494 47856 43546
rect 47610 43492 47616 43494
rect 47672 43492 47696 43494
rect 47752 43492 47776 43494
rect 47832 43492 47856 43494
rect 47912 43492 47918 43494
rect 47610 43483 47918 43492
rect 52610 43548 52918 43557
rect 52610 43546 52616 43548
rect 52672 43546 52696 43548
rect 52752 43546 52776 43548
rect 52832 43546 52856 43548
rect 52912 43546 52918 43548
rect 52672 43494 52674 43546
rect 52854 43494 52856 43546
rect 52610 43492 52616 43494
rect 52672 43492 52696 43494
rect 52752 43492 52776 43494
rect 52832 43492 52856 43494
rect 52912 43492 52918 43494
rect 52610 43483 52918 43492
rect 57610 43548 57918 43557
rect 57610 43546 57616 43548
rect 57672 43546 57696 43548
rect 57752 43546 57776 43548
rect 57832 43546 57856 43548
rect 57912 43546 57918 43548
rect 57672 43494 57674 43546
rect 57854 43494 57856 43546
rect 57610 43492 57616 43494
rect 57672 43492 57696 43494
rect 57752 43492 57776 43494
rect 57832 43492 57856 43494
rect 57912 43492 57918 43494
rect 57610 43483 57918 43492
rect 58544 43353 58572 43726
rect 58530 43344 58586 43353
rect 58530 43279 58586 43288
rect 1950 43004 2258 43013
rect 1950 43002 1956 43004
rect 2012 43002 2036 43004
rect 2092 43002 2116 43004
rect 2172 43002 2196 43004
rect 2252 43002 2258 43004
rect 2012 42950 2014 43002
rect 2194 42950 2196 43002
rect 1950 42948 1956 42950
rect 2012 42948 2036 42950
rect 2092 42948 2116 42950
rect 2172 42948 2196 42950
rect 2252 42948 2258 42950
rect 1950 42939 2258 42948
rect 6950 43004 7258 43013
rect 6950 43002 6956 43004
rect 7012 43002 7036 43004
rect 7092 43002 7116 43004
rect 7172 43002 7196 43004
rect 7252 43002 7258 43004
rect 7012 42950 7014 43002
rect 7194 42950 7196 43002
rect 6950 42948 6956 42950
rect 7012 42948 7036 42950
rect 7092 42948 7116 42950
rect 7172 42948 7196 42950
rect 7252 42948 7258 42950
rect 6950 42939 7258 42948
rect 11950 43004 12258 43013
rect 11950 43002 11956 43004
rect 12012 43002 12036 43004
rect 12092 43002 12116 43004
rect 12172 43002 12196 43004
rect 12252 43002 12258 43004
rect 12012 42950 12014 43002
rect 12194 42950 12196 43002
rect 11950 42948 11956 42950
rect 12012 42948 12036 42950
rect 12092 42948 12116 42950
rect 12172 42948 12196 42950
rect 12252 42948 12258 42950
rect 11950 42939 12258 42948
rect 16950 43004 17258 43013
rect 16950 43002 16956 43004
rect 17012 43002 17036 43004
rect 17092 43002 17116 43004
rect 17172 43002 17196 43004
rect 17252 43002 17258 43004
rect 17012 42950 17014 43002
rect 17194 42950 17196 43002
rect 16950 42948 16956 42950
rect 17012 42948 17036 42950
rect 17092 42948 17116 42950
rect 17172 42948 17196 42950
rect 17252 42948 17258 42950
rect 16950 42939 17258 42948
rect 21950 43004 22258 43013
rect 21950 43002 21956 43004
rect 22012 43002 22036 43004
rect 22092 43002 22116 43004
rect 22172 43002 22196 43004
rect 22252 43002 22258 43004
rect 22012 42950 22014 43002
rect 22194 42950 22196 43002
rect 21950 42948 21956 42950
rect 22012 42948 22036 42950
rect 22092 42948 22116 42950
rect 22172 42948 22196 42950
rect 22252 42948 22258 42950
rect 21950 42939 22258 42948
rect 26950 43004 27258 43013
rect 26950 43002 26956 43004
rect 27012 43002 27036 43004
rect 27092 43002 27116 43004
rect 27172 43002 27196 43004
rect 27252 43002 27258 43004
rect 27012 42950 27014 43002
rect 27194 42950 27196 43002
rect 26950 42948 26956 42950
rect 27012 42948 27036 42950
rect 27092 42948 27116 42950
rect 27172 42948 27196 42950
rect 27252 42948 27258 42950
rect 26950 42939 27258 42948
rect 31950 43004 32258 43013
rect 31950 43002 31956 43004
rect 32012 43002 32036 43004
rect 32092 43002 32116 43004
rect 32172 43002 32196 43004
rect 32252 43002 32258 43004
rect 32012 42950 32014 43002
rect 32194 42950 32196 43002
rect 31950 42948 31956 42950
rect 32012 42948 32036 42950
rect 32092 42948 32116 42950
rect 32172 42948 32196 42950
rect 32252 42948 32258 42950
rect 31950 42939 32258 42948
rect 36950 43004 37258 43013
rect 36950 43002 36956 43004
rect 37012 43002 37036 43004
rect 37092 43002 37116 43004
rect 37172 43002 37196 43004
rect 37252 43002 37258 43004
rect 37012 42950 37014 43002
rect 37194 42950 37196 43002
rect 36950 42948 36956 42950
rect 37012 42948 37036 42950
rect 37092 42948 37116 42950
rect 37172 42948 37196 42950
rect 37252 42948 37258 42950
rect 36950 42939 37258 42948
rect 41950 43004 42258 43013
rect 41950 43002 41956 43004
rect 42012 43002 42036 43004
rect 42092 43002 42116 43004
rect 42172 43002 42196 43004
rect 42252 43002 42258 43004
rect 42012 42950 42014 43002
rect 42194 42950 42196 43002
rect 41950 42948 41956 42950
rect 42012 42948 42036 42950
rect 42092 42948 42116 42950
rect 42172 42948 42196 42950
rect 42252 42948 42258 42950
rect 41950 42939 42258 42948
rect 46950 43004 47258 43013
rect 46950 43002 46956 43004
rect 47012 43002 47036 43004
rect 47092 43002 47116 43004
rect 47172 43002 47196 43004
rect 47252 43002 47258 43004
rect 47012 42950 47014 43002
rect 47194 42950 47196 43002
rect 46950 42948 46956 42950
rect 47012 42948 47036 42950
rect 47092 42948 47116 42950
rect 47172 42948 47196 42950
rect 47252 42948 47258 42950
rect 46950 42939 47258 42948
rect 51950 43004 52258 43013
rect 51950 43002 51956 43004
rect 52012 43002 52036 43004
rect 52092 43002 52116 43004
rect 52172 43002 52196 43004
rect 52252 43002 52258 43004
rect 52012 42950 52014 43002
rect 52194 42950 52196 43002
rect 51950 42948 51956 42950
rect 52012 42948 52036 42950
rect 52092 42948 52116 42950
rect 52172 42948 52196 42950
rect 52252 42948 52258 42950
rect 51950 42939 52258 42948
rect 56950 43004 57258 43013
rect 56950 43002 56956 43004
rect 57012 43002 57036 43004
rect 57092 43002 57116 43004
rect 57172 43002 57196 43004
rect 57252 43002 57258 43004
rect 57012 42950 57014 43002
rect 57194 42950 57196 43002
rect 56950 42948 56956 42950
rect 57012 42948 57036 42950
rect 57092 42948 57116 42950
rect 57172 42948 57196 42950
rect 57252 42948 57258 42950
rect 56950 42939 57258 42948
rect 58532 42696 58584 42702
rect 58532 42638 58584 42644
rect 58544 42537 58572 42638
rect 58530 42528 58586 42537
rect 2610 42460 2918 42469
rect 2610 42458 2616 42460
rect 2672 42458 2696 42460
rect 2752 42458 2776 42460
rect 2832 42458 2856 42460
rect 2912 42458 2918 42460
rect 2672 42406 2674 42458
rect 2854 42406 2856 42458
rect 2610 42404 2616 42406
rect 2672 42404 2696 42406
rect 2752 42404 2776 42406
rect 2832 42404 2856 42406
rect 2912 42404 2918 42406
rect 2610 42395 2918 42404
rect 7610 42460 7918 42469
rect 7610 42458 7616 42460
rect 7672 42458 7696 42460
rect 7752 42458 7776 42460
rect 7832 42458 7856 42460
rect 7912 42458 7918 42460
rect 7672 42406 7674 42458
rect 7854 42406 7856 42458
rect 7610 42404 7616 42406
rect 7672 42404 7696 42406
rect 7752 42404 7776 42406
rect 7832 42404 7856 42406
rect 7912 42404 7918 42406
rect 7610 42395 7918 42404
rect 12610 42460 12918 42469
rect 12610 42458 12616 42460
rect 12672 42458 12696 42460
rect 12752 42458 12776 42460
rect 12832 42458 12856 42460
rect 12912 42458 12918 42460
rect 12672 42406 12674 42458
rect 12854 42406 12856 42458
rect 12610 42404 12616 42406
rect 12672 42404 12696 42406
rect 12752 42404 12776 42406
rect 12832 42404 12856 42406
rect 12912 42404 12918 42406
rect 12610 42395 12918 42404
rect 17610 42460 17918 42469
rect 17610 42458 17616 42460
rect 17672 42458 17696 42460
rect 17752 42458 17776 42460
rect 17832 42458 17856 42460
rect 17912 42458 17918 42460
rect 17672 42406 17674 42458
rect 17854 42406 17856 42458
rect 17610 42404 17616 42406
rect 17672 42404 17696 42406
rect 17752 42404 17776 42406
rect 17832 42404 17856 42406
rect 17912 42404 17918 42406
rect 17610 42395 17918 42404
rect 22610 42460 22918 42469
rect 22610 42458 22616 42460
rect 22672 42458 22696 42460
rect 22752 42458 22776 42460
rect 22832 42458 22856 42460
rect 22912 42458 22918 42460
rect 22672 42406 22674 42458
rect 22854 42406 22856 42458
rect 22610 42404 22616 42406
rect 22672 42404 22696 42406
rect 22752 42404 22776 42406
rect 22832 42404 22856 42406
rect 22912 42404 22918 42406
rect 22610 42395 22918 42404
rect 27610 42460 27918 42469
rect 27610 42458 27616 42460
rect 27672 42458 27696 42460
rect 27752 42458 27776 42460
rect 27832 42458 27856 42460
rect 27912 42458 27918 42460
rect 27672 42406 27674 42458
rect 27854 42406 27856 42458
rect 27610 42404 27616 42406
rect 27672 42404 27696 42406
rect 27752 42404 27776 42406
rect 27832 42404 27856 42406
rect 27912 42404 27918 42406
rect 27610 42395 27918 42404
rect 32610 42460 32918 42469
rect 32610 42458 32616 42460
rect 32672 42458 32696 42460
rect 32752 42458 32776 42460
rect 32832 42458 32856 42460
rect 32912 42458 32918 42460
rect 32672 42406 32674 42458
rect 32854 42406 32856 42458
rect 32610 42404 32616 42406
rect 32672 42404 32696 42406
rect 32752 42404 32776 42406
rect 32832 42404 32856 42406
rect 32912 42404 32918 42406
rect 32610 42395 32918 42404
rect 37610 42460 37918 42469
rect 37610 42458 37616 42460
rect 37672 42458 37696 42460
rect 37752 42458 37776 42460
rect 37832 42458 37856 42460
rect 37912 42458 37918 42460
rect 37672 42406 37674 42458
rect 37854 42406 37856 42458
rect 37610 42404 37616 42406
rect 37672 42404 37696 42406
rect 37752 42404 37776 42406
rect 37832 42404 37856 42406
rect 37912 42404 37918 42406
rect 37610 42395 37918 42404
rect 42610 42460 42918 42469
rect 42610 42458 42616 42460
rect 42672 42458 42696 42460
rect 42752 42458 42776 42460
rect 42832 42458 42856 42460
rect 42912 42458 42918 42460
rect 42672 42406 42674 42458
rect 42854 42406 42856 42458
rect 42610 42404 42616 42406
rect 42672 42404 42696 42406
rect 42752 42404 42776 42406
rect 42832 42404 42856 42406
rect 42912 42404 42918 42406
rect 42610 42395 42918 42404
rect 47610 42460 47918 42469
rect 47610 42458 47616 42460
rect 47672 42458 47696 42460
rect 47752 42458 47776 42460
rect 47832 42458 47856 42460
rect 47912 42458 47918 42460
rect 47672 42406 47674 42458
rect 47854 42406 47856 42458
rect 47610 42404 47616 42406
rect 47672 42404 47696 42406
rect 47752 42404 47776 42406
rect 47832 42404 47856 42406
rect 47912 42404 47918 42406
rect 47610 42395 47918 42404
rect 52610 42460 52918 42469
rect 52610 42458 52616 42460
rect 52672 42458 52696 42460
rect 52752 42458 52776 42460
rect 52832 42458 52856 42460
rect 52912 42458 52918 42460
rect 52672 42406 52674 42458
rect 52854 42406 52856 42458
rect 52610 42404 52616 42406
rect 52672 42404 52696 42406
rect 52752 42404 52776 42406
rect 52832 42404 52856 42406
rect 52912 42404 52918 42406
rect 52610 42395 52918 42404
rect 57610 42460 57918 42469
rect 58530 42463 58586 42472
rect 57610 42458 57616 42460
rect 57672 42458 57696 42460
rect 57752 42458 57776 42460
rect 57832 42458 57856 42460
rect 57912 42458 57918 42460
rect 57672 42406 57674 42458
rect 57854 42406 57856 42458
rect 57610 42404 57616 42406
rect 57672 42404 57696 42406
rect 57752 42404 57776 42406
rect 57832 42404 57856 42406
rect 57912 42404 57918 42406
rect 57610 42395 57918 42404
rect 58532 42016 58584 42022
rect 58532 41958 58584 41964
rect 1950 41916 2258 41925
rect 1950 41914 1956 41916
rect 2012 41914 2036 41916
rect 2092 41914 2116 41916
rect 2172 41914 2196 41916
rect 2252 41914 2258 41916
rect 2012 41862 2014 41914
rect 2194 41862 2196 41914
rect 1950 41860 1956 41862
rect 2012 41860 2036 41862
rect 2092 41860 2116 41862
rect 2172 41860 2196 41862
rect 2252 41860 2258 41862
rect 1950 41851 2258 41860
rect 6950 41916 7258 41925
rect 6950 41914 6956 41916
rect 7012 41914 7036 41916
rect 7092 41914 7116 41916
rect 7172 41914 7196 41916
rect 7252 41914 7258 41916
rect 7012 41862 7014 41914
rect 7194 41862 7196 41914
rect 6950 41860 6956 41862
rect 7012 41860 7036 41862
rect 7092 41860 7116 41862
rect 7172 41860 7196 41862
rect 7252 41860 7258 41862
rect 6950 41851 7258 41860
rect 11950 41916 12258 41925
rect 11950 41914 11956 41916
rect 12012 41914 12036 41916
rect 12092 41914 12116 41916
rect 12172 41914 12196 41916
rect 12252 41914 12258 41916
rect 12012 41862 12014 41914
rect 12194 41862 12196 41914
rect 11950 41860 11956 41862
rect 12012 41860 12036 41862
rect 12092 41860 12116 41862
rect 12172 41860 12196 41862
rect 12252 41860 12258 41862
rect 11950 41851 12258 41860
rect 16950 41916 17258 41925
rect 16950 41914 16956 41916
rect 17012 41914 17036 41916
rect 17092 41914 17116 41916
rect 17172 41914 17196 41916
rect 17252 41914 17258 41916
rect 17012 41862 17014 41914
rect 17194 41862 17196 41914
rect 16950 41860 16956 41862
rect 17012 41860 17036 41862
rect 17092 41860 17116 41862
rect 17172 41860 17196 41862
rect 17252 41860 17258 41862
rect 16950 41851 17258 41860
rect 21950 41916 22258 41925
rect 21950 41914 21956 41916
rect 22012 41914 22036 41916
rect 22092 41914 22116 41916
rect 22172 41914 22196 41916
rect 22252 41914 22258 41916
rect 22012 41862 22014 41914
rect 22194 41862 22196 41914
rect 21950 41860 21956 41862
rect 22012 41860 22036 41862
rect 22092 41860 22116 41862
rect 22172 41860 22196 41862
rect 22252 41860 22258 41862
rect 21950 41851 22258 41860
rect 26950 41916 27258 41925
rect 26950 41914 26956 41916
rect 27012 41914 27036 41916
rect 27092 41914 27116 41916
rect 27172 41914 27196 41916
rect 27252 41914 27258 41916
rect 27012 41862 27014 41914
rect 27194 41862 27196 41914
rect 26950 41860 26956 41862
rect 27012 41860 27036 41862
rect 27092 41860 27116 41862
rect 27172 41860 27196 41862
rect 27252 41860 27258 41862
rect 26950 41851 27258 41860
rect 31950 41916 32258 41925
rect 31950 41914 31956 41916
rect 32012 41914 32036 41916
rect 32092 41914 32116 41916
rect 32172 41914 32196 41916
rect 32252 41914 32258 41916
rect 32012 41862 32014 41914
rect 32194 41862 32196 41914
rect 31950 41860 31956 41862
rect 32012 41860 32036 41862
rect 32092 41860 32116 41862
rect 32172 41860 32196 41862
rect 32252 41860 32258 41862
rect 31950 41851 32258 41860
rect 36950 41916 37258 41925
rect 36950 41914 36956 41916
rect 37012 41914 37036 41916
rect 37092 41914 37116 41916
rect 37172 41914 37196 41916
rect 37252 41914 37258 41916
rect 37012 41862 37014 41914
rect 37194 41862 37196 41914
rect 36950 41860 36956 41862
rect 37012 41860 37036 41862
rect 37092 41860 37116 41862
rect 37172 41860 37196 41862
rect 37252 41860 37258 41862
rect 36950 41851 37258 41860
rect 41950 41916 42258 41925
rect 41950 41914 41956 41916
rect 42012 41914 42036 41916
rect 42092 41914 42116 41916
rect 42172 41914 42196 41916
rect 42252 41914 42258 41916
rect 42012 41862 42014 41914
rect 42194 41862 42196 41914
rect 41950 41860 41956 41862
rect 42012 41860 42036 41862
rect 42092 41860 42116 41862
rect 42172 41860 42196 41862
rect 42252 41860 42258 41862
rect 41950 41851 42258 41860
rect 46950 41916 47258 41925
rect 46950 41914 46956 41916
rect 47012 41914 47036 41916
rect 47092 41914 47116 41916
rect 47172 41914 47196 41916
rect 47252 41914 47258 41916
rect 47012 41862 47014 41914
rect 47194 41862 47196 41914
rect 46950 41860 46956 41862
rect 47012 41860 47036 41862
rect 47092 41860 47116 41862
rect 47172 41860 47196 41862
rect 47252 41860 47258 41862
rect 46950 41851 47258 41860
rect 51950 41916 52258 41925
rect 51950 41914 51956 41916
rect 52012 41914 52036 41916
rect 52092 41914 52116 41916
rect 52172 41914 52196 41916
rect 52252 41914 52258 41916
rect 52012 41862 52014 41914
rect 52194 41862 52196 41914
rect 51950 41860 51956 41862
rect 52012 41860 52036 41862
rect 52092 41860 52116 41862
rect 52172 41860 52196 41862
rect 52252 41860 52258 41862
rect 51950 41851 52258 41860
rect 56950 41916 57258 41925
rect 56950 41914 56956 41916
rect 57012 41914 57036 41916
rect 57092 41914 57116 41916
rect 57172 41914 57196 41916
rect 57252 41914 57258 41916
rect 57012 41862 57014 41914
rect 57194 41862 57196 41914
rect 56950 41860 56956 41862
rect 57012 41860 57036 41862
rect 57092 41860 57116 41862
rect 57172 41860 57196 41862
rect 57252 41860 57258 41862
rect 56950 41851 57258 41860
rect 58544 41721 58572 41958
rect 58530 41712 58586 41721
rect 58530 41647 58586 41656
rect 2610 41372 2918 41381
rect 2610 41370 2616 41372
rect 2672 41370 2696 41372
rect 2752 41370 2776 41372
rect 2832 41370 2856 41372
rect 2912 41370 2918 41372
rect 2672 41318 2674 41370
rect 2854 41318 2856 41370
rect 2610 41316 2616 41318
rect 2672 41316 2696 41318
rect 2752 41316 2776 41318
rect 2832 41316 2856 41318
rect 2912 41316 2918 41318
rect 2610 41307 2918 41316
rect 7610 41372 7918 41381
rect 7610 41370 7616 41372
rect 7672 41370 7696 41372
rect 7752 41370 7776 41372
rect 7832 41370 7856 41372
rect 7912 41370 7918 41372
rect 7672 41318 7674 41370
rect 7854 41318 7856 41370
rect 7610 41316 7616 41318
rect 7672 41316 7696 41318
rect 7752 41316 7776 41318
rect 7832 41316 7856 41318
rect 7912 41316 7918 41318
rect 7610 41307 7918 41316
rect 12610 41372 12918 41381
rect 12610 41370 12616 41372
rect 12672 41370 12696 41372
rect 12752 41370 12776 41372
rect 12832 41370 12856 41372
rect 12912 41370 12918 41372
rect 12672 41318 12674 41370
rect 12854 41318 12856 41370
rect 12610 41316 12616 41318
rect 12672 41316 12696 41318
rect 12752 41316 12776 41318
rect 12832 41316 12856 41318
rect 12912 41316 12918 41318
rect 12610 41307 12918 41316
rect 17610 41372 17918 41381
rect 17610 41370 17616 41372
rect 17672 41370 17696 41372
rect 17752 41370 17776 41372
rect 17832 41370 17856 41372
rect 17912 41370 17918 41372
rect 17672 41318 17674 41370
rect 17854 41318 17856 41370
rect 17610 41316 17616 41318
rect 17672 41316 17696 41318
rect 17752 41316 17776 41318
rect 17832 41316 17856 41318
rect 17912 41316 17918 41318
rect 17610 41307 17918 41316
rect 22610 41372 22918 41381
rect 22610 41370 22616 41372
rect 22672 41370 22696 41372
rect 22752 41370 22776 41372
rect 22832 41370 22856 41372
rect 22912 41370 22918 41372
rect 22672 41318 22674 41370
rect 22854 41318 22856 41370
rect 22610 41316 22616 41318
rect 22672 41316 22696 41318
rect 22752 41316 22776 41318
rect 22832 41316 22856 41318
rect 22912 41316 22918 41318
rect 22610 41307 22918 41316
rect 27610 41372 27918 41381
rect 27610 41370 27616 41372
rect 27672 41370 27696 41372
rect 27752 41370 27776 41372
rect 27832 41370 27856 41372
rect 27912 41370 27918 41372
rect 27672 41318 27674 41370
rect 27854 41318 27856 41370
rect 27610 41316 27616 41318
rect 27672 41316 27696 41318
rect 27752 41316 27776 41318
rect 27832 41316 27856 41318
rect 27912 41316 27918 41318
rect 27610 41307 27918 41316
rect 32610 41372 32918 41381
rect 32610 41370 32616 41372
rect 32672 41370 32696 41372
rect 32752 41370 32776 41372
rect 32832 41370 32856 41372
rect 32912 41370 32918 41372
rect 32672 41318 32674 41370
rect 32854 41318 32856 41370
rect 32610 41316 32616 41318
rect 32672 41316 32696 41318
rect 32752 41316 32776 41318
rect 32832 41316 32856 41318
rect 32912 41316 32918 41318
rect 32610 41307 32918 41316
rect 37610 41372 37918 41381
rect 37610 41370 37616 41372
rect 37672 41370 37696 41372
rect 37752 41370 37776 41372
rect 37832 41370 37856 41372
rect 37912 41370 37918 41372
rect 37672 41318 37674 41370
rect 37854 41318 37856 41370
rect 37610 41316 37616 41318
rect 37672 41316 37696 41318
rect 37752 41316 37776 41318
rect 37832 41316 37856 41318
rect 37912 41316 37918 41318
rect 37610 41307 37918 41316
rect 42610 41372 42918 41381
rect 42610 41370 42616 41372
rect 42672 41370 42696 41372
rect 42752 41370 42776 41372
rect 42832 41370 42856 41372
rect 42912 41370 42918 41372
rect 42672 41318 42674 41370
rect 42854 41318 42856 41370
rect 42610 41316 42616 41318
rect 42672 41316 42696 41318
rect 42752 41316 42776 41318
rect 42832 41316 42856 41318
rect 42912 41316 42918 41318
rect 42610 41307 42918 41316
rect 47610 41372 47918 41381
rect 47610 41370 47616 41372
rect 47672 41370 47696 41372
rect 47752 41370 47776 41372
rect 47832 41370 47856 41372
rect 47912 41370 47918 41372
rect 47672 41318 47674 41370
rect 47854 41318 47856 41370
rect 47610 41316 47616 41318
rect 47672 41316 47696 41318
rect 47752 41316 47776 41318
rect 47832 41316 47856 41318
rect 47912 41316 47918 41318
rect 47610 41307 47918 41316
rect 52610 41372 52918 41381
rect 52610 41370 52616 41372
rect 52672 41370 52696 41372
rect 52752 41370 52776 41372
rect 52832 41370 52856 41372
rect 52912 41370 52918 41372
rect 52672 41318 52674 41370
rect 52854 41318 52856 41370
rect 52610 41316 52616 41318
rect 52672 41316 52696 41318
rect 52752 41316 52776 41318
rect 52832 41316 52856 41318
rect 52912 41316 52918 41318
rect 52610 41307 52918 41316
rect 57610 41372 57918 41381
rect 57610 41370 57616 41372
rect 57672 41370 57696 41372
rect 57752 41370 57776 41372
rect 57832 41370 57856 41372
rect 57912 41370 57918 41372
rect 57672 41318 57674 41370
rect 57854 41318 57856 41370
rect 57610 41316 57616 41318
rect 57672 41316 57696 41318
rect 57752 41316 57776 41318
rect 57832 41316 57856 41318
rect 57912 41316 57918 41318
rect 57610 41307 57918 41316
rect 58532 40928 58584 40934
rect 58530 40896 58532 40905
rect 58584 40896 58586 40905
rect 1950 40828 2258 40837
rect 1950 40826 1956 40828
rect 2012 40826 2036 40828
rect 2092 40826 2116 40828
rect 2172 40826 2196 40828
rect 2252 40826 2258 40828
rect 2012 40774 2014 40826
rect 2194 40774 2196 40826
rect 1950 40772 1956 40774
rect 2012 40772 2036 40774
rect 2092 40772 2116 40774
rect 2172 40772 2196 40774
rect 2252 40772 2258 40774
rect 1950 40763 2258 40772
rect 6950 40828 7258 40837
rect 6950 40826 6956 40828
rect 7012 40826 7036 40828
rect 7092 40826 7116 40828
rect 7172 40826 7196 40828
rect 7252 40826 7258 40828
rect 7012 40774 7014 40826
rect 7194 40774 7196 40826
rect 6950 40772 6956 40774
rect 7012 40772 7036 40774
rect 7092 40772 7116 40774
rect 7172 40772 7196 40774
rect 7252 40772 7258 40774
rect 6950 40763 7258 40772
rect 11950 40828 12258 40837
rect 11950 40826 11956 40828
rect 12012 40826 12036 40828
rect 12092 40826 12116 40828
rect 12172 40826 12196 40828
rect 12252 40826 12258 40828
rect 12012 40774 12014 40826
rect 12194 40774 12196 40826
rect 11950 40772 11956 40774
rect 12012 40772 12036 40774
rect 12092 40772 12116 40774
rect 12172 40772 12196 40774
rect 12252 40772 12258 40774
rect 11950 40763 12258 40772
rect 16950 40828 17258 40837
rect 16950 40826 16956 40828
rect 17012 40826 17036 40828
rect 17092 40826 17116 40828
rect 17172 40826 17196 40828
rect 17252 40826 17258 40828
rect 17012 40774 17014 40826
rect 17194 40774 17196 40826
rect 16950 40772 16956 40774
rect 17012 40772 17036 40774
rect 17092 40772 17116 40774
rect 17172 40772 17196 40774
rect 17252 40772 17258 40774
rect 16950 40763 17258 40772
rect 21950 40828 22258 40837
rect 21950 40826 21956 40828
rect 22012 40826 22036 40828
rect 22092 40826 22116 40828
rect 22172 40826 22196 40828
rect 22252 40826 22258 40828
rect 22012 40774 22014 40826
rect 22194 40774 22196 40826
rect 21950 40772 21956 40774
rect 22012 40772 22036 40774
rect 22092 40772 22116 40774
rect 22172 40772 22196 40774
rect 22252 40772 22258 40774
rect 21950 40763 22258 40772
rect 26950 40828 27258 40837
rect 26950 40826 26956 40828
rect 27012 40826 27036 40828
rect 27092 40826 27116 40828
rect 27172 40826 27196 40828
rect 27252 40826 27258 40828
rect 27012 40774 27014 40826
rect 27194 40774 27196 40826
rect 26950 40772 26956 40774
rect 27012 40772 27036 40774
rect 27092 40772 27116 40774
rect 27172 40772 27196 40774
rect 27252 40772 27258 40774
rect 26950 40763 27258 40772
rect 31950 40828 32258 40837
rect 31950 40826 31956 40828
rect 32012 40826 32036 40828
rect 32092 40826 32116 40828
rect 32172 40826 32196 40828
rect 32252 40826 32258 40828
rect 32012 40774 32014 40826
rect 32194 40774 32196 40826
rect 31950 40772 31956 40774
rect 32012 40772 32036 40774
rect 32092 40772 32116 40774
rect 32172 40772 32196 40774
rect 32252 40772 32258 40774
rect 31950 40763 32258 40772
rect 36950 40828 37258 40837
rect 36950 40826 36956 40828
rect 37012 40826 37036 40828
rect 37092 40826 37116 40828
rect 37172 40826 37196 40828
rect 37252 40826 37258 40828
rect 37012 40774 37014 40826
rect 37194 40774 37196 40826
rect 36950 40772 36956 40774
rect 37012 40772 37036 40774
rect 37092 40772 37116 40774
rect 37172 40772 37196 40774
rect 37252 40772 37258 40774
rect 36950 40763 37258 40772
rect 41950 40828 42258 40837
rect 41950 40826 41956 40828
rect 42012 40826 42036 40828
rect 42092 40826 42116 40828
rect 42172 40826 42196 40828
rect 42252 40826 42258 40828
rect 42012 40774 42014 40826
rect 42194 40774 42196 40826
rect 41950 40772 41956 40774
rect 42012 40772 42036 40774
rect 42092 40772 42116 40774
rect 42172 40772 42196 40774
rect 42252 40772 42258 40774
rect 41950 40763 42258 40772
rect 46950 40828 47258 40837
rect 46950 40826 46956 40828
rect 47012 40826 47036 40828
rect 47092 40826 47116 40828
rect 47172 40826 47196 40828
rect 47252 40826 47258 40828
rect 47012 40774 47014 40826
rect 47194 40774 47196 40826
rect 46950 40772 46956 40774
rect 47012 40772 47036 40774
rect 47092 40772 47116 40774
rect 47172 40772 47196 40774
rect 47252 40772 47258 40774
rect 46950 40763 47258 40772
rect 51950 40828 52258 40837
rect 51950 40826 51956 40828
rect 52012 40826 52036 40828
rect 52092 40826 52116 40828
rect 52172 40826 52196 40828
rect 52252 40826 52258 40828
rect 52012 40774 52014 40826
rect 52194 40774 52196 40826
rect 51950 40772 51956 40774
rect 52012 40772 52036 40774
rect 52092 40772 52116 40774
rect 52172 40772 52196 40774
rect 52252 40772 52258 40774
rect 51950 40763 52258 40772
rect 56950 40828 57258 40837
rect 58530 40831 58586 40840
rect 56950 40826 56956 40828
rect 57012 40826 57036 40828
rect 57092 40826 57116 40828
rect 57172 40826 57196 40828
rect 57252 40826 57258 40828
rect 57012 40774 57014 40826
rect 57194 40774 57196 40826
rect 56950 40772 56956 40774
rect 57012 40772 57036 40774
rect 57092 40772 57116 40774
rect 57172 40772 57196 40774
rect 57252 40772 57258 40774
rect 56950 40763 57258 40772
rect 58532 40520 58584 40526
rect 58532 40462 58584 40468
rect 2610 40284 2918 40293
rect 2610 40282 2616 40284
rect 2672 40282 2696 40284
rect 2752 40282 2776 40284
rect 2832 40282 2856 40284
rect 2912 40282 2918 40284
rect 2672 40230 2674 40282
rect 2854 40230 2856 40282
rect 2610 40228 2616 40230
rect 2672 40228 2696 40230
rect 2752 40228 2776 40230
rect 2832 40228 2856 40230
rect 2912 40228 2918 40230
rect 2610 40219 2918 40228
rect 7610 40284 7918 40293
rect 7610 40282 7616 40284
rect 7672 40282 7696 40284
rect 7752 40282 7776 40284
rect 7832 40282 7856 40284
rect 7912 40282 7918 40284
rect 7672 40230 7674 40282
rect 7854 40230 7856 40282
rect 7610 40228 7616 40230
rect 7672 40228 7696 40230
rect 7752 40228 7776 40230
rect 7832 40228 7856 40230
rect 7912 40228 7918 40230
rect 7610 40219 7918 40228
rect 12610 40284 12918 40293
rect 12610 40282 12616 40284
rect 12672 40282 12696 40284
rect 12752 40282 12776 40284
rect 12832 40282 12856 40284
rect 12912 40282 12918 40284
rect 12672 40230 12674 40282
rect 12854 40230 12856 40282
rect 12610 40228 12616 40230
rect 12672 40228 12696 40230
rect 12752 40228 12776 40230
rect 12832 40228 12856 40230
rect 12912 40228 12918 40230
rect 12610 40219 12918 40228
rect 17610 40284 17918 40293
rect 17610 40282 17616 40284
rect 17672 40282 17696 40284
rect 17752 40282 17776 40284
rect 17832 40282 17856 40284
rect 17912 40282 17918 40284
rect 17672 40230 17674 40282
rect 17854 40230 17856 40282
rect 17610 40228 17616 40230
rect 17672 40228 17696 40230
rect 17752 40228 17776 40230
rect 17832 40228 17856 40230
rect 17912 40228 17918 40230
rect 17610 40219 17918 40228
rect 22610 40284 22918 40293
rect 22610 40282 22616 40284
rect 22672 40282 22696 40284
rect 22752 40282 22776 40284
rect 22832 40282 22856 40284
rect 22912 40282 22918 40284
rect 22672 40230 22674 40282
rect 22854 40230 22856 40282
rect 22610 40228 22616 40230
rect 22672 40228 22696 40230
rect 22752 40228 22776 40230
rect 22832 40228 22856 40230
rect 22912 40228 22918 40230
rect 22610 40219 22918 40228
rect 27610 40284 27918 40293
rect 27610 40282 27616 40284
rect 27672 40282 27696 40284
rect 27752 40282 27776 40284
rect 27832 40282 27856 40284
rect 27912 40282 27918 40284
rect 27672 40230 27674 40282
rect 27854 40230 27856 40282
rect 27610 40228 27616 40230
rect 27672 40228 27696 40230
rect 27752 40228 27776 40230
rect 27832 40228 27856 40230
rect 27912 40228 27918 40230
rect 27610 40219 27918 40228
rect 32610 40284 32918 40293
rect 32610 40282 32616 40284
rect 32672 40282 32696 40284
rect 32752 40282 32776 40284
rect 32832 40282 32856 40284
rect 32912 40282 32918 40284
rect 32672 40230 32674 40282
rect 32854 40230 32856 40282
rect 32610 40228 32616 40230
rect 32672 40228 32696 40230
rect 32752 40228 32776 40230
rect 32832 40228 32856 40230
rect 32912 40228 32918 40230
rect 32610 40219 32918 40228
rect 37610 40284 37918 40293
rect 37610 40282 37616 40284
rect 37672 40282 37696 40284
rect 37752 40282 37776 40284
rect 37832 40282 37856 40284
rect 37912 40282 37918 40284
rect 37672 40230 37674 40282
rect 37854 40230 37856 40282
rect 37610 40228 37616 40230
rect 37672 40228 37696 40230
rect 37752 40228 37776 40230
rect 37832 40228 37856 40230
rect 37912 40228 37918 40230
rect 37610 40219 37918 40228
rect 42610 40284 42918 40293
rect 42610 40282 42616 40284
rect 42672 40282 42696 40284
rect 42752 40282 42776 40284
rect 42832 40282 42856 40284
rect 42912 40282 42918 40284
rect 42672 40230 42674 40282
rect 42854 40230 42856 40282
rect 42610 40228 42616 40230
rect 42672 40228 42696 40230
rect 42752 40228 42776 40230
rect 42832 40228 42856 40230
rect 42912 40228 42918 40230
rect 42610 40219 42918 40228
rect 47610 40284 47918 40293
rect 47610 40282 47616 40284
rect 47672 40282 47696 40284
rect 47752 40282 47776 40284
rect 47832 40282 47856 40284
rect 47912 40282 47918 40284
rect 47672 40230 47674 40282
rect 47854 40230 47856 40282
rect 47610 40228 47616 40230
rect 47672 40228 47696 40230
rect 47752 40228 47776 40230
rect 47832 40228 47856 40230
rect 47912 40228 47918 40230
rect 47610 40219 47918 40228
rect 52610 40284 52918 40293
rect 52610 40282 52616 40284
rect 52672 40282 52696 40284
rect 52752 40282 52776 40284
rect 52832 40282 52856 40284
rect 52912 40282 52918 40284
rect 52672 40230 52674 40282
rect 52854 40230 52856 40282
rect 52610 40228 52616 40230
rect 52672 40228 52696 40230
rect 52752 40228 52776 40230
rect 52832 40228 52856 40230
rect 52912 40228 52918 40230
rect 52610 40219 52918 40228
rect 57610 40284 57918 40293
rect 57610 40282 57616 40284
rect 57672 40282 57696 40284
rect 57752 40282 57776 40284
rect 57832 40282 57856 40284
rect 57912 40282 57918 40284
rect 57672 40230 57674 40282
rect 57854 40230 57856 40282
rect 57610 40228 57616 40230
rect 57672 40228 57696 40230
rect 57752 40228 57776 40230
rect 57832 40228 57856 40230
rect 57912 40228 57918 40230
rect 57610 40219 57918 40228
rect 58544 40089 58572 40462
rect 58530 40080 58586 40089
rect 58530 40015 58586 40024
rect 1950 39740 2258 39749
rect 1950 39738 1956 39740
rect 2012 39738 2036 39740
rect 2092 39738 2116 39740
rect 2172 39738 2196 39740
rect 2252 39738 2258 39740
rect 2012 39686 2014 39738
rect 2194 39686 2196 39738
rect 1950 39684 1956 39686
rect 2012 39684 2036 39686
rect 2092 39684 2116 39686
rect 2172 39684 2196 39686
rect 2252 39684 2258 39686
rect 1950 39675 2258 39684
rect 6950 39740 7258 39749
rect 6950 39738 6956 39740
rect 7012 39738 7036 39740
rect 7092 39738 7116 39740
rect 7172 39738 7196 39740
rect 7252 39738 7258 39740
rect 7012 39686 7014 39738
rect 7194 39686 7196 39738
rect 6950 39684 6956 39686
rect 7012 39684 7036 39686
rect 7092 39684 7116 39686
rect 7172 39684 7196 39686
rect 7252 39684 7258 39686
rect 6950 39675 7258 39684
rect 11950 39740 12258 39749
rect 11950 39738 11956 39740
rect 12012 39738 12036 39740
rect 12092 39738 12116 39740
rect 12172 39738 12196 39740
rect 12252 39738 12258 39740
rect 12012 39686 12014 39738
rect 12194 39686 12196 39738
rect 11950 39684 11956 39686
rect 12012 39684 12036 39686
rect 12092 39684 12116 39686
rect 12172 39684 12196 39686
rect 12252 39684 12258 39686
rect 11950 39675 12258 39684
rect 16950 39740 17258 39749
rect 16950 39738 16956 39740
rect 17012 39738 17036 39740
rect 17092 39738 17116 39740
rect 17172 39738 17196 39740
rect 17252 39738 17258 39740
rect 17012 39686 17014 39738
rect 17194 39686 17196 39738
rect 16950 39684 16956 39686
rect 17012 39684 17036 39686
rect 17092 39684 17116 39686
rect 17172 39684 17196 39686
rect 17252 39684 17258 39686
rect 16950 39675 17258 39684
rect 21950 39740 22258 39749
rect 21950 39738 21956 39740
rect 22012 39738 22036 39740
rect 22092 39738 22116 39740
rect 22172 39738 22196 39740
rect 22252 39738 22258 39740
rect 22012 39686 22014 39738
rect 22194 39686 22196 39738
rect 21950 39684 21956 39686
rect 22012 39684 22036 39686
rect 22092 39684 22116 39686
rect 22172 39684 22196 39686
rect 22252 39684 22258 39686
rect 21950 39675 22258 39684
rect 26950 39740 27258 39749
rect 26950 39738 26956 39740
rect 27012 39738 27036 39740
rect 27092 39738 27116 39740
rect 27172 39738 27196 39740
rect 27252 39738 27258 39740
rect 27012 39686 27014 39738
rect 27194 39686 27196 39738
rect 26950 39684 26956 39686
rect 27012 39684 27036 39686
rect 27092 39684 27116 39686
rect 27172 39684 27196 39686
rect 27252 39684 27258 39686
rect 26950 39675 27258 39684
rect 31950 39740 32258 39749
rect 31950 39738 31956 39740
rect 32012 39738 32036 39740
rect 32092 39738 32116 39740
rect 32172 39738 32196 39740
rect 32252 39738 32258 39740
rect 32012 39686 32014 39738
rect 32194 39686 32196 39738
rect 31950 39684 31956 39686
rect 32012 39684 32036 39686
rect 32092 39684 32116 39686
rect 32172 39684 32196 39686
rect 32252 39684 32258 39686
rect 31950 39675 32258 39684
rect 36950 39740 37258 39749
rect 36950 39738 36956 39740
rect 37012 39738 37036 39740
rect 37092 39738 37116 39740
rect 37172 39738 37196 39740
rect 37252 39738 37258 39740
rect 37012 39686 37014 39738
rect 37194 39686 37196 39738
rect 36950 39684 36956 39686
rect 37012 39684 37036 39686
rect 37092 39684 37116 39686
rect 37172 39684 37196 39686
rect 37252 39684 37258 39686
rect 36950 39675 37258 39684
rect 41950 39740 42258 39749
rect 41950 39738 41956 39740
rect 42012 39738 42036 39740
rect 42092 39738 42116 39740
rect 42172 39738 42196 39740
rect 42252 39738 42258 39740
rect 42012 39686 42014 39738
rect 42194 39686 42196 39738
rect 41950 39684 41956 39686
rect 42012 39684 42036 39686
rect 42092 39684 42116 39686
rect 42172 39684 42196 39686
rect 42252 39684 42258 39686
rect 41950 39675 42258 39684
rect 46950 39740 47258 39749
rect 46950 39738 46956 39740
rect 47012 39738 47036 39740
rect 47092 39738 47116 39740
rect 47172 39738 47196 39740
rect 47252 39738 47258 39740
rect 47012 39686 47014 39738
rect 47194 39686 47196 39738
rect 46950 39684 46956 39686
rect 47012 39684 47036 39686
rect 47092 39684 47116 39686
rect 47172 39684 47196 39686
rect 47252 39684 47258 39686
rect 46950 39675 47258 39684
rect 51950 39740 52258 39749
rect 51950 39738 51956 39740
rect 52012 39738 52036 39740
rect 52092 39738 52116 39740
rect 52172 39738 52196 39740
rect 52252 39738 52258 39740
rect 52012 39686 52014 39738
rect 52194 39686 52196 39738
rect 51950 39684 51956 39686
rect 52012 39684 52036 39686
rect 52092 39684 52116 39686
rect 52172 39684 52196 39686
rect 52252 39684 52258 39686
rect 51950 39675 52258 39684
rect 56950 39740 57258 39749
rect 56950 39738 56956 39740
rect 57012 39738 57036 39740
rect 57092 39738 57116 39740
rect 57172 39738 57196 39740
rect 57252 39738 57258 39740
rect 57012 39686 57014 39738
rect 57194 39686 57196 39738
rect 56950 39684 56956 39686
rect 57012 39684 57036 39686
rect 57092 39684 57116 39686
rect 57172 39684 57196 39686
rect 57252 39684 57258 39686
rect 56950 39675 57258 39684
rect 58532 39432 58584 39438
rect 58532 39374 58584 39380
rect 58544 39273 58572 39374
rect 58530 39264 58586 39273
rect 2610 39196 2918 39205
rect 2610 39194 2616 39196
rect 2672 39194 2696 39196
rect 2752 39194 2776 39196
rect 2832 39194 2856 39196
rect 2912 39194 2918 39196
rect 2672 39142 2674 39194
rect 2854 39142 2856 39194
rect 2610 39140 2616 39142
rect 2672 39140 2696 39142
rect 2752 39140 2776 39142
rect 2832 39140 2856 39142
rect 2912 39140 2918 39142
rect 2610 39131 2918 39140
rect 7610 39196 7918 39205
rect 7610 39194 7616 39196
rect 7672 39194 7696 39196
rect 7752 39194 7776 39196
rect 7832 39194 7856 39196
rect 7912 39194 7918 39196
rect 7672 39142 7674 39194
rect 7854 39142 7856 39194
rect 7610 39140 7616 39142
rect 7672 39140 7696 39142
rect 7752 39140 7776 39142
rect 7832 39140 7856 39142
rect 7912 39140 7918 39142
rect 7610 39131 7918 39140
rect 12610 39196 12918 39205
rect 12610 39194 12616 39196
rect 12672 39194 12696 39196
rect 12752 39194 12776 39196
rect 12832 39194 12856 39196
rect 12912 39194 12918 39196
rect 12672 39142 12674 39194
rect 12854 39142 12856 39194
rect 12610 39140 12616 39142
rect 12672 39140 12696 39142
rect 12752 39140 12776 39142
rect 12832 39140 12856 39142
rect 12912 39140 12918 39142
rect 12610 39131 12918 39140
rect 17610 39196 17918 39205
rect 17610 39194 17616 39196
rect 17672 39194 17696 39196
rect 17752 39194 17776 39196
rect 17832 39194 17856 39196
rect 17912 39194 17918 39196
rect 17672 39142 17674 39194
rect 17854 39142 17856 39194
rect 17610 39140 17616 39142
rect 17672 39140 17696 39142
rect 17752 39140 17776 39142
rect 17832 39140 17856 39142
rect 17912 39140 17918 39142
rect 17610 39131 17918 39140
rect 22610 39196 22918 39205
rect 22610 39194 22616 39196
rect 22672 39194 22696 39196
rect 22752 39194 22776 39196
rect 22832 39194 22856 39196
rect 22912 39194 22918 39196
rect 22672 39142 22674 39194
rect 22854 39142 22856 39194
rect 22610 39140 22616 39142
rect 22672 39140 22696 39142
rect 22752 39140 22776 39142
rect 22832 39140 22856 39142
rect 22912 39140 22918 39142
rect 22610 39131 22918 39140
rect 27610 39196 27918 39205
rect 27610 39194 27616 39196
rect 27672 39194 27696 39196
rect 27752 39194 27776 39196
rect 27832 39194 27856 39196
rect 27912 39194 27918 39196
rect 27672 39142 27674 39194
rect 27854 39142 27856 39194
rect 27610 39140 27616 39142
rect 27672 39140 27696 39142
rect 27752 39140 27776 39142
rect 27832 39140 27856 39142
rect 27912 39140 27918 39142
rect 27610 39131 27918 39140
rect 32610 39196 32918 39205
rect 32610 39194 32616 39196
rect 32672 39194 32696 39196
rect 32752 39194 32776 39196
rect 32832 39194 32856 39196
rect 32912 39194 32918 39196
rect 32672 39142 32674 39194
rect 32854 39142 32856 39194
rect 32610 39140 32616 39142
rect 32672 39140 32696 39142
rect 32752 39140 32776 39142
rect 32832 39140 32856 39142
rect 32912 39140 32918 39142
rect 32610 39131 32918 39140
rect 37610 39196 37918 39205
rect 37610 39194 37616 39196
rect 37672 39194 37696 39196
rect 37752 39194 37776 39196
rect 37832 39194 37856 39196
rect 37912 39194 37918 39196
rect 37672 39142 37674 39194
rect 37854 39142 37856 39194
rect 37610 39140 37616 39142
rect 37672 39140 37696 39142
rect 37752 39140 37776 39142
rect 37832 39140 37856 39142
rect 37912 39140 37918 39142
rect 37610 39131 37918 39140
rect 42610 39196 42918 39205
rect 42610 39194 42616 39196
rect 42672 39194 42696 39196
rect 42752 39194 42776 39196
rect 42832 39194 42856 39196
rect 42912 39194 42918 39196
rect 42672 39142 42674 39194
rect 42854 39142 42856 39194
rect 42610 39140 42616 39142
rect 42672 39140 42696 39142
rect 42752 39140 42776 39142
rect 42832 39140 42856 39142
rect 42912 39140 42918 39142
rect 42610 39131 42918 39140
rect 47610 39196 47918 39205
rect 47610 39194 47616 39196
rect 47672 39194 47696 39196
rect 47752 39194 47776 39196
rect 47832 39194 47856 39196
rect 47912 39194 47918 39196
rect 47672 39142 47674 39194
rect 47854 39142 47856 39194
rect 47610 39140 47616 39142
rect 47672 39140 47696 39142
rect 47752 39140 47776 39142
rect 47832 39140 47856 39142
rect 47912 39140 47918 39142
rect 47610 39131 47918 39140
rect 52610 39196 52918 39205
rect 52610 39194 52616 39196
rect 52672 39194 52696 39196
rect 52752 39194 52776 39196
rect 52832 39194 52856 39196
rect 52912 39194 52918 39196
rect 52672 39142 52674 39194
rect 52854 39142 52856 39194
rect 52610 39140 52616 39142
rect 52672 39140 52696 39142
rect 52752 39140 52776 39142
rect 52832 39140 52856 39142
rect 52912 39140 52918 39142
rect 52610 39131 52918 39140
rect 57610 39196 57918 39205
rect 58530 39199 58586 39208
rect 57610 39194 57616 39196
rect 57672 39194 57696 39196
rect 57752 39194 57776 39196
rect 57832 39194 57856 39196
rect 57912 39194 57918 39196
rect 57672 39142 57674 39194
rect 57854 39142 57856 39194
rect 57610 39140 57616 39142
rect 57672 39140 57696 39142
rect 57752 39140 57776 39142
rect 57832 39140 57856 39142
rect 57912 39140 57918 39142
rect 57610 39131 57918 39140
rect 58532 38752 58584 38758
rect 58532 38694 58584 38700
rect 1950 38652 2258 38661
rect 1950 38650 1956 38652
rect 2012 38650 2036 38652
rect 2092 38650 2116 38652
rect 2172 38650 2196 38652
rect 2252 38650 2258 38652
rect 2012 38598 2014 38650
rect 2194 38598 2196 38650
rect 1950 38596 1956 38598
rect 2012 38596 2036 38598
rect 2092 38596 2116 38598
rect 2172 38596 2196 38598
rect 2252 38596 2258 38598
rect 1950 38587 2258 38596
rect 6950 38652 7258 38661
rect 6950 38650 6956 38652
rect 7012 38650 7036 38652
rect 7092 38650 7116 38652
rect 7172 38650 7196 38652
rect 7252 38650 7258 38652
rect 7012 38598 7014 38650
rect 7194 38598 7196 38650
rect 6950 38596 6956 38598
rect 7012 38596 7036 38598
rect 7092 38596 7116 38598
rect 7172 38596 7196 38598
rect 7252 38596 7258 38598
rect 6950 38587 7258 38596
rect 11950 38652 12258 38661
rect 11950 38650 11956 38652
rect 12012 38650 12036 38652
rect 12092 38650 12116 38652
rect 12172 38650 12196 38652
rect 12252 38650 12258 38652
rect 12012 38598 12014 38650
rect 12194 38598 12196 38650
rect 11950 38596 11956 38598
rect 12012 38596 12036 38598
rect 12092 38596 12116 38598
rect 12172 38596 12196 38598
rect 12252 38596 12258 38598
rect 11950 38587 12258 38596
rect 16950 38652 17258 38661
rect 16950 38650 16956 38652
rect 17012 38650 17036 38652
rect 17092 38650 17116 38652
rect 17172 38650 17196 38652
rect 17252 38650 17258 38652
rect 17012 38598 17014 38650
rect 17194 38598 17196 38650
rect 16950 38596 16956 38598
rect 17012 38596 17036 38598
rect 17092 38596 17116 38598
rect 17172 38596 17196 38598
rect 17252 38596 17258 38598
rect 16950 38587 17258 38596
rect 21950 38652 22258 38661
rect 21950 38650 21956 38652
rect 22012 38650 22036 38652
rect 22092 38650 22116 38652
rect 22172 38650 22196 38652
rect 22252 38650 22258 38652
rect 22012 38598 22014 38650
rect 22194 38598 22196 38650
rect 21950 38596 21956 38598
rect 22012 38596 22036 38598
rect 22092 38596 22116 38598
rect 22172 38596 22196 38598
rect 22252 38596 22258 38598
rect 21950 38587 22258 38596
rect 26950 38652 27258 38661
rect 26950 38650 26956 38652
rect 27012 38650 27036 38652
rect 27092 38650 27116 38652
rect 27172 38650 27196 38652
rect 27252 38650 27258 38652
rect 27012 38598 27014 38650
rect 27194 38598 27196 38650
rect 26950 38596 26956 38598
rect 27012 38596 27036 38598
rect 27092 38596 27116 38598
rect 27172 38596 27196 38598
rect 27252 38596 27258 38598
rect 26950 38587 27258 38596
rect 31950 38652 32258 38661
rect 31950 38650 31956 38652
rect 32012 38650 32036 38652
rect 32092 38650 32116 38652
rect 32172 38650 32196 38652
rect 32252 38650 32258 38652
rect 32012 38598 32014 38650
rect 32194 38598 32196 38650
rect 31950 38596 31956 38598
rect 32012 38596 32036 38598
rect 32092 38596 32116 38598
rect 32172 38596 32196 38598
rect 32252 38596 32258 38598
rect 31950 38587 32258 38596
rect 36950 38652 37258 38661
rect 36950 38650 36956 38652
rect 37012 38650 37036 38652
rect 37092 38650 37116 38652
rect 37172 38650 37196 38652
rect 37252 38650 37258 38652
rect 37012 38598 37014 38650
rect 37194 38598 37196 38650
rect 36950 38596 36956 38598
rect 37012 38596 37036 38598
rect 37092 38596 37116 38598
rect 37172 38596 37196 38598
rect 37252 38596 37258 38598
rect 36950 38587 37258 38596
rect 41950 38652 42258 38661
rect 41950 38650 41956 38652
rect 42012 38650 42036 38652
rect 42092 38650 42116 38652
rect 42172 38650 42196 38652
rect 42252 38650 42258 38652
rect 42012 38598 42014 38650
rect 42194 38598 42196 38650
rect 41950 38596 41956 38598
rect 42012 38596 42036 38598
rect 42092 38596 42116 38598
rect 42172 38596 42196 38598
rect 42252 38596 42258 38598
rect 41950 38587 42258 38596
rect 46950 38652 47258 38661
rect 46950 38650 46956 38652
rect 47012 38650 47036 38652
rect 47092 38650 47116 38652
rect 47172 38650 47196 38652
rect 47252 38650 47258 38652
rect 47012 38598 47014 38650
rect 47194 38598 47196 38650
rect 46950 38596 46956 38598
rect 47012 38596 47036 38598
rect 47092 38596 47116 38598
rect 47172 38596 47196 38598
rect 47252 38596 47258 38598
rect 46950 38587 47258 38596
rect 51950 38652 52258 38661
rect 51950 38650 51956 38652
rect 52012 38650 52036 38652
rect 52092 38650 52116 38652
rect 52172 38650 52196 38652
rect 52252 38650 52258 38652
rect 52012 38598 52014 38650
rect 52194 38598 52196 38650
rect 51950 38596 51956 38598
rect 52012 38596 52036 38598
rect 52092 38596 52116 38598
rect 52172 38596 52196 38598
rect 52252 38596 52258 38598
rect 51950 38587 52258 38596
rect 56950 38652 57258 38661
rect 56950 38650 56956 38652
rect 57012 38650 57036 38652
rect 57092 38650 57116 38652
rect 57172 38650 57196 38652
rect 57252 38650 57258 38652
rect 57012 38598 57014 38650
rect 57194 38598 57196 38650
rect 56950 38596 56956 38598
rect 57012 38596 57036 38598
rect 57092 38596 57116 38598
rect 57172 38596 57196 38598
rect 57252 38596 57258 38598
rect 56950 38587 57258 38596
rect 58544 38457 58572 38694
rect 58530 38448 58586 38457
rect 58530 38383 58586 38392
rect 2610 38108 2918 38117
rect 2610 38106 2616 38108
rect 2672 38106 2696 38108
rect 2752 38106 2776 38108
rect 2832 38106 2856 38108
rect 2912 38106 2918 38108
rect 2672 38054 2674 38106
rect 2854 38054 2856 38106
rect 2610 38052 2616 38054
rect 2672 38052 2696 38054
rect 2752 38052 2776 38054
rect 2832 38052 2856 38054
rect 2912 38052 2918 38054
rect 2610 38043 2918 38052
rect 7610 38108 7918 38117
rect 7610 38106 7616 38108
rect 7672 38106 7696 38108
rect 7752 38106 7776 38108
rect 7832 38106 7856 38108
rect 7912 38106 7918 38108
rect 7672 38054 7674 38106
rect 7854 38054 7856 38106
rect 7610 38052 7616 38054
rect 7672 38052 7696 38054
rect 7752 38052 7776 38054
rect 7832 38052 7856 38054
rect 7912 38052 7918 38054
rect 7610 38043 7918 38052
rect 12610 38108 12918 38117
rect 12610 38106 12616 38108
rect 12672 38106 12696 38108
rect 12752 38106 12776 38108
rect 12832 38106 12856 38108
rect 12912 38106 12918 38108
rect 12672 38054 12674 38106
rect 12854 38054 12856 38106
rect 12610 38052 12616 38054
rect 12672 38052 12696 38054
rect 12752 38052 12776 38054
rect 12832 38052 12856 38054
rect 12912 38052 12918 38054
rect 12610 38043 12918 38052
rect 17610 38108 17918 38117
rect 17610 38106 17616 38108
rect 17672 38106 17696 38108
rect 17752 38106 17776 38108
rect 17832 38106 17856 38108
rect 17912 38106 17918 38108
rect 17672 38054 17674 38106
rect 17854 38054 17856 38106
rect 17610 38052 17616 38054
rect 17672 38052 17696 38054
rect 17752 38052 17776 38054
rect 17832 38052 17856 38054
rect 17912 38052 17918 38054
rect 17610 38043 17918 38052
rect 22610 38108 22918 38117
rect 22610 38106 22616 38108
rect 22672 38106 22696 38108
rect 22752 38106 22776 38108
rect 22832 38106 22856 38108
rect 22912 38106 22918 38108
rect 22672 38054 22674 38106
rect 22854 38054 22856 38106
rect 22610 38052 22616 38054
rect 22672 38052 22696 38054
rect 22752 38052 22776 38054
rect 22832 38052 22856 38054
rect 22912 38052 22918 38054
rect 22610 38043 22918 38052
rect 27610 38108 27918 38117
rect 27610 38106 27616 38108
rect 27672 38106 27696 38108
rect 27752 38106 27776 38108
rect 27832 38106 27856 38108
rect 27912 38106 27918 38108
rect 27672 38054 27674 38106
rect 27854 38054 27856 38106
rect 27610 38052 27616 38054
rect 27672 38052 27696 38054
rect 27752 38052 27776 38054
rect 27832 38052 27856 38054
rect 27912 38052 27918 38054
rect 27610 38043 27918 38052
rect 32610 38108 32918 38117
rect 32610 38106 32616 38108
rect 32672 38106 32696 38108
rect 32752 38106 32776 38108
rect 32832 38106 32856 38108
rect 32912 38106 32918 38108
rect 32672 38054 32674 38106
rect 32854 38054 32856 38106
rect 32610 38052 32616 38054
rect 32672 38052 32696 38054
rect 32752 38052 32776 38054
rect 32832 38052 32856 38054
rect 32912 38052 32918 38054
rect 32610 38043 32918 38052
rect 37610 38108 37918 38117
rect 37610 38106 37616 38108
rect 37672 38106 37696 38108
rect 37752 38106 37776 38108
rect 37832 38106 37856 38108
rect 37912 38106 37918 38108
rect 37672 38054 37674 38106
rect 37854 38054 37856 38106
rect 37610 38052 37616 38054
rect 37672 38052 37696 38054
rect 37752 38052 37776 38054
rect 37832 38052 37856 38054
rect 37912 38052 37918 38054
rect 37610 38043 37918 38052
rect 42610 38108 42918 38117
rect 42610 38106 42616 38108
rect 42672 38106 42696 38108
rect 42752 38106 42776 38108
rect 42832 38106 42856 38108
rect 42912 38106 42918 38108
rect 42672 38054 42674 38106
rect 42854 38054 42856 38106
rect 42610 38052 42616 38054
rect 42672 38052 42696 38054
rect 42752 38052 42776 38054
rect 42832 38052 42856 38054
rect 42912 38052 42918 38054
rect 42610 38043 42918 38052
rect 47610 38108 47918 38117
rect 47610 38106 47616 38108
rect 47672 38106 47696 38108
rect 47752 38106 47776 38108
rect 47832 38106 47856 38108
rect 47912 38106 47918 38108
rect 47672 38054 47674 38106
rect 47854 38054 47856 38106
rect 47610 38052 47616 38054
rect 47672 38052 47696 38054
rect 47752 38052 47776 38054
rect 47832 38052 47856 38054
rect 47912 38052 47918 38054
rect 47610 38043 47918 38052
rect 52610 38108 52918 38117
rect 52610 38106 52616 38108
rect 52672 38106 52696 38108
rect 52752 38106 52776 38108
rect 52832 38106 52856 38108
rect 52912 38106 52918 38108
rect 52672 38054 52674 38106
rect 52854 38054 52856 38106
rect 52610 38052 52616 38054
rect 52672 38052 52696 38054
rect 52752 38052 52776 38054
rect 52832 38052 52856 38054
rect 52912 38052 52918 38054
rect 52610 38043 52918 38052
rect 57610 38108 57918 38117
rect 57610 38106 57616 38108
rect 57672 38106 57696 38108
rect 57752 38106 57776 38108
rect 57832 38106 57856 38108
rect 57912 38106 57918 38108
rect 57672 38054 57674 38106
rect 57854 38054 57856 38106
rect 57610 38052 57616 38054
rect 57672 38052 57696 38054
rect 57752 38052 57776 38054
rect 57832 38052 57856 38054
rect 57912 38052 57918 38054
rect 57610 38043 57918 38052
rect 58532 37664 58584 37670
rect 58530 37632 58532 37641
rect 58584 37632 58586 37641
rect 1950 37564 2258 37573
rect 1950 37562 1956 37564
rect 2012 37562 2036 37564
rect 2092 37562 2116 37564
rect 2172 37562 2196 37564
rect 2252 37562 2258 37564
rect 2012 37510 2014 37562
rect 2194 37510 2196 37562
rect 1950 37508 1956 37510
rect 2012 37508 2036 37510
rect 2092 37508 2116 37510
rect 2172 37508 2196 37510
rect 2252 37508 2258 37510
rect 1950 37499 2258 37508
rect 6950 37564 7258 37573
rect 6950 37562 6956 37564
rect 7012 37562 7036 37564
rect 7092 37562 7116 37564
rect 7172 37562 7196 37564
rect 7252 37562 7258 37564
rect 7012 37510 7014 37562
rect 7194 37510 7196 37562
rect 6950 37508 6956 37510
rect 7012 37508 7036 37510
rect 7092 37508 7116 37510
rect 7172 37508 7196 37510
rect 7252 37508 7258 37510
rect 6950 37499 7258 37508
rect 11950 37564 12258 37573
rect 11950 37562 11956 37564
rect 12012 37562 12036 37564
rect 12092 37562 12116 37564
rect 12172 37562 12196 37564
rect 12252 37562 12258 37564
rect 12012 37510 12014 37562
rect 12194 37510 12196 37562
rect 11950 37508 11956 37510
rect 12012 37508 12036 37510
rect 12092 37508 12116 37510
rect 12172 37508 12196 37510
rect 12252 37508 12258 37510
rect 11950 37499 12258 37508
rect 16950 37564 17258 37573
rect 16950 37562 16956 37564
rect 17012 37562 17036 37564
rect 17092 37562 17116 37564
rect 17172 37562 17196 37564
rect 17252 37562 17258 37564
rect 17012 37510 17014 37562
rect 17194 37510 17196 37562
rect 16950 37508 16956 37510
rect 17012 37508 17036 37510
rect 17092 37508 17116 37510
rect 17172 37508 17196 37510
rect 17252 37508 17258 37510
rect 16950 37499 17258 37508
rect 21950 37564 22258 37573
rect 21950 37562 21956 37564
rect 22012 37562 22036 37564
rect 22092 37562 22116 37564
rect 22172 37562 22196 37564
rect 22252 37562 22258 37564
rect 22012 37510 22014 37562
rect 22194 37510 22196 37562
rect 21950 37508 21956 37510
rect 22012 37508 22036 37510
rect 22092 37508 22116 37510
rect 22172 37508 22196 37510
rect 22252 37508 22258 37510
rect 21950 37499 22258 37508
rect 26950 37564 27258 37573
rect 26950 37562 26956 37564
rect 27012 37562 27036 37564
rect 27092 37562 27116 37564
rect 27172 37562 27196 37564
rect 27252 37562 27258 37564
rect 27012 37510 27014 37562
rect 27194 37510 27196 37562
rect 26950 37508 26956 37510
rect 27012 37508 27036 37510
rect 27092 37508 27116 37510
rect 27172 37508 27196 37510
rect 27252 37508 27258 37510
rect 26950 37499 27258 37508
rect 31950 37564 32258 37573
rect 31950 37562 31956 37564
rect 32012 37562 32036 37564
rect 32092 37562 32116 37564
rect 32172 37562 32196 37564
rect 32252 37562 32258 37564
rect 32012 37510 32014 37562
rect 32194 37510 32196 37562
rect 31950 37508 31956 37510
rect 32012 37508 32036 37510
rect 32092 37508 32116 37510
rect 32172 37508 32196 37510
rect 32252 37508 32258 37510
rect 31950 37499 32258 37508
rect 36950 37564 37258 37573
rect 36950 37562 36956 37564
rect 37012 37562 37036 37564
rect 37092 37562 37116 37564
rect 37172 37562 37196 37564
rect 37252 37562 37258 37564
rect 37012 37510 37014 37562
rect 37194 37510 37196 37562
rect 36950 37508 36956 37510
rect 37012 37508 37036 37510
rect 37092 37508 37116 37510
rect 37172 37508 37196 37510
rect 37252 37508 37258 37510
rect 36950 37499 37258 37508
rect 41950 37564 42258 37573
rect 41950 37562 41956 37564
rect 42012 37562 42036 37564
rect 42092 37562 42116 37564
rect 42172 37562 42196 37564
rect 42252 37562 42258 37564
rect 42012 37510 42014 37562
rect 42194 37510 42196 37562
rect 41950 37508 41956 37510
rect 42012 37508 42036 37510
rect 42092 37508 42116 37510
rect 42172 37508 42196 37510
rect 42252 37508 42258 37510
rect 41950 37499 42258 37508
rect 46950 37564 47258 37573
rect 46950 37562 46956 37564
rect 47012 37562 47036 37564
rect 47092 37562 47116 37564
rect 47172 37562 47196 37564
rect 47252 37562 47258 37564
rect 47012 37510 47014 37562
rect 47194 37510 47196 37562
rect 46950 37508 46956 37510
rect 47012 37508 47036 37510
rect 47092 37508 47116 37510
rect 47172 37508 47196 37510
rect 47252 37508 47258 37510
rect 46950 37499 47258 37508
rect 51950 37564 52258 37573
rect 51950 37562 51956 37564
rect 52012 37562 52036 37564
rect 52092 37562 52116 37564
rect 52172 37562 52196 37564
rect 52252 37562 52258 37564
rect 52012 37510 52014 37562
rect 52194 37510 52196 37562
rect 51950 37508 51956 37510
rect 52012 37508 52036 37510
rect 52092 37508 52116 37510
rect 52172 37508 52196 37510
rect 52252 37508 52258 37510
rect 51950 37499 52258 37508
rect 56950 37564 57258 37573
rect 58530 37567 58586 37576
rect 56950 37562 56956 37564
rect 57012 37562 57036 37564
rect 57092 37562 57116 37564
rect 57172 37562 57196 37564
rect 57252 37562 57258 37564
rect 57012 37510 57014 37562
rect 57194 37510 57196 37562
rect 56950 37508 56956 37510
rect 57012 37508 57036 37510
rect 57092 37508 57116 37510
rect 57172 37508 57196 37510
rect 57252 37508 57258 37510
rect 56950 37499 57258 37508
rect 58532 37324 58584 37330
rect 58532 37266 58584 37272
rect 2610 37020 2918 37029
rect 2610 37018 2616 37020
rect 2672 37018 2696 37020
rect 2752 37018 2776 37020
rect 2832 37018 2856 37020
rect 2912 37018 2918 37020
rect 2672 36966 2674 37018
rect 2854 36966 2856 37018
rect 2610 36964 2616 36966
rect 2672 36964 2696 36966
rect 2752 36964 2776 36966
rect 2832 36964 2856 36966
rect 2912 36964 2918 36966
rect 2610 36955 2918 36964
rect 7610 37020 7918 37029
rect 7610 37018 7616 37020
rect 7672 37018 7696 37020
rect 7752 37018 7776 37020
rect 7832 37018 7856 37020
rect 7912 37018 7918 37020
rect 7672 36966 7674 37018
rect 7854 36966 7856 37018
rect 7610 36964 7616 36966
rect 7672 36964 7696 36966
rect 7752 36964 7776 36966
rect 7832 36964 7856 36966
rect 7912 36964 7918 36966
rect 7610 36955 7918 36964
rect 12610 37020 12918 37029
rect 12610 37018 12616 37020
rect 12672 37018 12696 37020
rect 12752 37018 12776 37020
rect 12832 37018 12856 37020
rect 12912 37018 12918 37020
rect 12672 36966 12674 37018
rect 12854 36966 12856 37018
rect 12610 36964 12616 36966
rect 12672 36964 12696 36966
rect 12752 36964 12776 36966
rect 12832 36964 12856 36966
rect 12912 36964 12918 36966
rect 12610 36955 12918 36964
rect 17610 37020 17918 37029
rect 17610 37018 17616 37020
rect 17672 37018 17696 37020
rect 17752 37018 17776 37020
rect 17832 37018 17856 37020
rect 17912 37018 17918 37020
rect 17672 36966 17674 37018
rect 17854 36966 17856 37018
rect 17610 36964 17616 36966
rect 17672 36964 17696 36966
rect 17752 36964 17776 36966
rect 17832 36964 17856 36966
rect 17912 36964 17918 36966
rect 17610 36955 17918 36964
rect 22610 37020 22918 37029
rect 22610 37018 22616 37020
rect 22672 37018 22696 37020
rect 22752 37018 22776 37020
rect 22832 37018 22856 37020
rect 22912 37018 22918 37020
rect 22672 36966 22674 37018
rect 22854 36966 22856 37018
rect 22610 36964 22616 36966
rect 22672 36964 22696 36966
rect 22752 36964 22776 36966
rect 22832 36964 22856 36966
rect 22912 36964 22918 36966
rect 22610 36955 22918 36964
rect 27610 37020 27918 37029
rect 27610 37018 27616 37020
rect 27672 37018 27696 37020
rect 27752 37018 27776 37020
rect 27832 37018 27856 37020
rect 27912 37018 27918 37020
rect 27672 36966 27674 37018
rect 27854 36966 27856 37018
rect 27610 36964 27616 36966
rect 27672 36964 27696 36966
rect 27752 36964 27776 36966
rect 27832 36964 27856 36966
rect 27912 36964 27918 36966
rect 27610 36955 27918 36964
rect 32610 37020 32918 37029
rect 32610 37018 32616 37020
rect 32672 37018 32696 37020
rect 32752 37018 32776 37020
rect 32832 37018 32856 37020
rect 32912 37018 32918 37020
rect 32672 36966 32674 37018
rect 32854 36966 32856 37018
rect 32610 36964 32616 36966
rect 32672 36964 32696 36966
rect 32752 36964 32776 36966
rect 32832 36964 32856 36966
rect 32912 36964 32918 36966
rect 32610 36955 32918 36964
rect 37610 37020 37918 37029
rect 37610 37018 37616 37020
rect 37672 37018 37696 37020
rect 37752 37018 37776 37020
rect 37832 37018 37856 37020
rect 37912 37018 37918 37020
rect 37672 36966 37674 37018
rect 37854 36966 37856 37018
rect 37610 36964 37616 36966
rect 37672 36964 37696 36966
rect 37752 36964 37776 36966
rect 37832 36964 37856 36966
rect 37912 36964 37918 36966
rect 37610 36955 37918 36964
rect 42610 37020 42918 37029
rect 42610 37018 42616 37020
rect 42672 37018 42696 37020
rect 42752 37018 42776 37020
rect 42832 37018 42856 37020
rect 42912 37018 42918 37020
rect 42672 36966 42674 37018
rect 42854 36966 42856 37018
rect 42610 36964 42616 36966
rect 42672 36964 42696 36966
rect 42752 36964 42776 36966
rect 42832 36964 42856 36966
rect 42912 36964 42918 36966
rect 42610 36955 42918 36964
rect 47610 37020 47918 37029
rect 47610 37018 47616 37020
rect 47672 37018 47696 37020
rect 47752 37018 47776 37020
rect 47832 37018 47856 37020
rect 47912 37018 47918 37020
rect 47672 36966 47674 37018
rect 47854 36966 47856 37018
rect 47610 36964 47616 36966
rect 47672 36964 47696 36966
rect 47752 36964 47776 36966
rect 47832 36964 47856 36966
rect 47912 36964 47918 36966
rect 47610 36955 47918 36964
rect 52610 37020 52918 37029
rect 52610 37018 52616 37020
rect 52672 37018 52696 37020
rect 52752 37018 52776 37020
rect 52832 37018 52856 37020
rect 52912 37018 52918 37020
rect 52672 36966 52674 37018
rect 52854 36966 52856 37018
rect 52610 36964 52616 36966
rect 52672 36964 52696 36966
rect 52752 36964 52776 36966
rect 52832 36964 52856 36966
rect 52912 36964 52918 36966
rect 52610 36955 52918 36964
rect 57610 37020 57918 37029
rect 57610 37018 57616 37020
rect 57672 37018 57696 37020
rect 57752 37018 57776 37020
rect 57832 37018 57856 37020
rect 57912 37018 57918 37020
rect 57672 36966 57674 37018
rect 57854 36966 57856 37018
rect 57610 36964 57616 36966
rect 57672 36964 57696 36966
rect 57752 36964 57776 36966
rect 57832 36964 57856 36966
rect 57912 36964 57918 36966
rect 57610 36955 57918 36964
rect 58544 36825 58572 37266
rect 58530 36816 58586 36825
rect 58530 36751 58586 36760
rect 1950 36476 2258 36485
rect 1950 36474 1956 36476
rect 2012 36474 2036 36476
rect 2092 36474 2116 36476
rect 2172 36474 2196 36476
rect 2252 36474 2258 36476
rect 2012 36422 2014 36474
rect 2194 36422 2196 36474
rect 1950 36420 1956 36422
rect 2012 36420 2036 36422
rect 2092 36420 2116 36422
rect 2172 36420 2196 36422
rect 2252 36420 2258 36422
rect 1950 36411 2258 36420
rect 6950 36476 7258 36485
rect 6950 36474 6956 36476
rect 7012 36474 7036 36476
rect 7092 36474 7116 36476
rect 7172 36474 7196 36476
rect 7252 36474 7258 36476
rect 7012 36422 7014 36474
rect 7194 36422 7196 36474
rect 6950 36420 6956 36422
rect 7012 36420 7036 36422
rect 7092 36420 7116 36422
rect 7172 36420 7196 36422
rect 7252 36420 7258 36422
rect 6950 36411 7258 36420
rect 11950 36476 12258 36485
rect 11950 36474 11956 36476
rect 12012 36474 12036 36476
rect 12092 36474 12116 36476
rect 12172 36474 12196 36476
rect 12252 36474 12258 36476
rect 12012 36422 12014 36474
rect 12194 36422 12196 36474
rect 11950 36420 11956 36422
rect 12012 36420 12036 36422
rect 12092 36420 12116 36422
rect 12172 36420 12196 36422
rect 12252 36420 12258 36422
rect 11950 36411 12258 36420
rect 16950 36476 17258 36485
rect 16950 36474 16956 36476
rect 17012 36474 17036 36476
rect 17092 36474 17116 36476
rect 17172 36474 17196 36476
rect 17252 36474 17258 36476
rect 17012 36422 17014 36474
rect 17194 36422 17196 36474
rect 16950 36420 16956 36422
rect 17012 36420 17036 36422
rect 17092 36420 17116 36422
rect 17172 36420 17196 36422
rect 17252 36420 17258 36422
rect 16950 36411 17258 36420
rect 21950 36476 22258 36485
rect 21950 36474 21956 36476
rect 22012 36474 22036 36476
rect 22092 36474 22116 36476
rect 22172 36474 22196 36476
rect 22252 36474 22258 36476
rect 22012 36422 22014 36474
rect 22194 36422 22196 36474
rect 21950 36420 21956 36422
rect 22012 36420 22036 36422
rect 22092 36420 22116 36422
rect 22172 36420 22196 36422
rect 22252 36420 22258 36422
rect 21950 36411 22258 36420
rect 26950 36476 27258 36485
rect 26950 36474 26956 36476
rect 27012 36474 27036 36476
rect 27092 36474 27116 36476
rect 27172 36474 27196 36476
rect 27252 36474 27258 36476
rect 27012 36422 27014 36474
rect 27194 36422 27196 36474
rect 26950 36420 26956 36422
rect 27012 36420 27036 36422
rect 27092 36420 27116 36422
rect 27172 36420 27196 36422
rect 27252 36420 27258 36422
rect 26950 36411 27258 36420
rect 31950 36476 32258 36485
rect 31950 36474 31956 36476
rect 32012 36474 32036 36476
rect 32092 36474 32116 36476
rect 32172 36474 32196 36476
rect 32252 36474 32258 36476
rect 32012 36422 32014 36474
rect 32194 36422 32196 36474
rect 31950 36420 31956 36422
rect 32012 36420 32036 36422
rect 32092 36420 32116 36422
rect 32172 36420 32196 36422
rect 32252 36420 32258 36422
rect 31950 36411 32258 36420
rect 36950 36476 37258 36485
rect 36950 36474 36956 36476
rect 37012 36474 37036 36476
rect 37092 36474 37116 36476
rect 37172 36474 37196 36476
rect 37252 36474 37258 36476
rect 37012 36422 37014 36474
rect 37194 36422 37196 36474
rect 36950 36420 36956 36422
rect 37012 36420 37036 36422
rect 37092 36420 37116 36422
rect 37172 36420 37196 36422
rect 37252 36420 37258 36422
rect 36950 36411 37258 36420
rect 41950 36476 42258 36485
rect 41950 36474 41956 36476
rect 42012 36474 42036 36476
rect 42092 36474 42116 36476
rect 42172 36474 42196 36476
rect 42252 36474 42258 36476
rect 42012 36422 42014 36474
rect 42194 36422 42196 36474
rect 41950 36420 41956 36422
rect 42012 36420 42036 36422
rect 42092 36420 42116 36422
rect 42172 36420 42196 36422
rect 42252 36420 42258 36422
rect 41950 36411 42258 36420
rect 46950 36476 47258 36485
rect 46950 36474 46956 36476
rect 47012 36474 47036 36476
rect 47092 36474 47116 36476
rect 47172 36474 47196 36476
rect 47252 36474 47258 36476
rect 47012 36422 47014 36474
rect 47194 36422 47196 36474
rect 46950 36420 46956 36422
rect 47012 36420 47036 36422
rect 47092 36420 47116 36422
rect 47172 36420 47196 36422
rect 47252 36420 47258 36422
rect 46950 36411 47258 36420
rect 51950 36476 52258 36485
rect 51950 36474 51956 36476
rect 52012 36474 52036 36476
rect 52092 36474 52116 36476
rect 52172 36474 52196 36476
rect 52252 36474 52258 36476
rect 52012 36422 52014 36474
rect 52194 36422 52196 36474
rect 51950 36420 51956 36422
rect 52012 36420 52036 36422
rect 52092 36420 52116 36422
rect 52172 36420 52196 36422
rect 52252 36420 52258 36422
rect 51950 36411 52258 36420
rect 56950 36476 57258 36485
rect 56950 36474 56956 36476
rect 57012 36474 57036 36476
rect 57092 36474 57116 36476
rect 57172 36474 57196 36476
rect 57252 36474 57258 36476
rect 57012 36422 57014 36474
rect 57194 36422 57196 36474
rect 56950 36420 56956 36422
rect 57012 36420 57036 36422
rect 57092 36420 57116 36422
rect 57172 36420 57196 36422
rect 57252 36420 57258 36422
rect 56950 36411 57258 36420
rect 58532 36168 58584 36174
rect 58532 36110 58584 36116
rect 58544 36009 58572 36110
rect 58530 36000 58586 36009
rect 2610 35932 2918 35941
rect 2610 35930 2616 35932
rect 2672 35930 2696 35932
rect 2752 35930 2776 35932
rect 2832 35930 2856 35932
rect 2912 35930 2918 35932
rect 2672 35878 2674 35930
rect 2854 35878 2856 35930
rect 2610 35876 2616 35878
rect 2672 35876 2696 35878
rect 2752 35876 2776 35878
rect 2832 35876 2856 35878
rect 2912 35876 2918 35878
rect 2610 35867 2918 35876
rect 7610 35932 7918 35941
rect 7610 35930 7616 35932
rect 7672 35930 7696 35932
rect 7752 35930 7776 35932
rect 7832 35930 7856 35932
rect 7912 35930 7918 35932
rect 7672 35878 7674 35930
rect 7854 35878 7856 35930
rect 7610 35876 7616 35878
rect 7672 35876 7696 35878
rect 7752 35876 7776 35878
rect 7832 35876 7856 35878
rect 7912 35876 7918 35878
rect 7610 35867 7918 35876
rect 12610 35932 12918 35941
rect 12610 35930 12616 35932
rect 12672 35930 12696 35932
rect 12752 35930 12776 35932
rect 12832 35930 12856 35932
rect 12912 35930 12918 35932
rect 12672 35878 12674 35930
rect 12854 35878 12856 35930
rect 12610 35876 12616 35878
rect 12672 35876 12696 35878
rect 12752 35876 12776 35878
rect 12832 35876 12856 35878
rect 12912 35876 12918 35878
rect 12610 35867 12918 35876
rect 17610 35932 17918 35941
rect 17610 35930 17616 35932
rect 17672 35930 17696 35932
rect 17752 35930 17776 35932
rect 17832 35930 17856 35932
rect 17912 35930 17918 35932
rect 17672 35878 17674 35930
rect 17854 35878 17856 35930
rect 17610 35876 17616 35878
rect 17672 35876 17696 35878
rect 17752 35876 17776 35878
rect 17832 35876 17856 35878
rect 17912 35876 17918 35878
rect 17610 35867 17918 35876
rect 22610 35932 22918 35941
rect 22610 35930 22616 35932
rect 22672 35930 22696 35932
rect 22752 35930 22776 35932
rect 22832 35930 22856 35932
rect 22912 35930 22918 35932
rect 22672 35878 22674 35930
rect 22854 35878 22856 35930
rect 22610 35876 22616 35878
rect 22672 35876 22696 35878
rect 22752 35876 22776 35878
rect 22832 35876 22856 35878
rect 22912 35876 22918 35878
rect 22610 35867 22918 35876
rect 27610 35932 27918 35941
rect 27610 35930 27616 35932
rect 27672 35930 27696 35932
rect 27752 35930 27776 35932
rect 27832 35930 27856 35932
rect 27912 35930 27918 35932
rect 27672 35878 27674 35930
rect 27854 35878 27856 35930
rect 27610 35876 27616 35878
rect 27672 35876 27696 35878
rect 27752 35876 27776 35878
rect 27832 35876 27856 35878
rect 27912 35876 27918 35878
rect 27610 35867 27918 35876
rect 32610 35932 32918 35941
rect 32610 35930 32616 35932
rect 32672 35930 32696 35932
rect 32752 35930 32776 35932
rect 32832 35930 32856 35932
rect 32912 35930 32918 35932
rect 32672 35878 32674 35930
rect 32854 35878 32856 35930
rect 32610 35876 32616 35878
rect 32672 35876 32696 35878
rect 32752 35876 32776 35878
rect 32832 35876 32856 35878
rect 32912 35876 32918 35878
rect 32610 35867 32918 35876
rect 37610 35932 37918 35941
rect 37610 35930 37616 35932
rect 37672 35930 37696 35932
rect 37752 35930 37776 35932
rect 37832 35930 37856 35932
rect 37912 35930 37918 35932
rect 37672 35878 37674 35930
rect 37854 35878 37856 35930
rect 37610 35876 37616 35878
rect 37672 35876 37696 35878
rect 37752 35876 37776 35878
rect 37832 35876 37856 35878
rect 37912 35876 37918 35878
rect 37610 35867 37918 35876
rect 42610 35932 42918 35941
rect 42610 35930 42616 35932
rect 42672 35930 42696 35932
rect 42752 35930 42776 35932
rect 42832 35930 42856 35932
rect 42912 35930 42918 35932
rect 42672 35878 42674 35930
rect 42854 35878 42856 35930
rect 42610 35876 42616 35878
rect 42672 35876 42696 35878
rect 42752 35876 42776 35878
rect 42832 35876 42856 35878
rect 42912 35876 42918 35878
rect 42610 35867 42918 35876
rect 47610 35932 47918 35941
rect 47610 35930 47616 35932
rect 47672 35930 47696 35932
rect 47752 35930 47776 35932
rect 47832 35930 47856 35932
rect 47912 35930 47918 35932
rect 47672 35878 47674 35930
rect 47854 35878 47856 35930
rect 47610 35876 47616 35878
rect 47672 35876 47696 35878
rect 47752 35876 47776 35878
rect 47832 35876 47856 35878
rect 47912 35876 47918 35878
rect 47610 35867 47918 35876
rect 52610 35932 52918 35941
rect 52610 35930 52616 35932
rect 52672 35930 52696 35932
rect 52752 35930 52776 35932
rect 52832 35930 52856 35932
rect 52912 35930 52918 35932
rect 52672 35878 52674 35930
rect 52854 35878 52856 35930
rect 52610 35876 52616 35878
rect 52672 35876 52696 35878
rect 52752 35876 52776 35878
rect 52832 35876 52856 35878
rect 52912 35876 52918 35878
rect 52610 35867 52918 35876
rect 57610 35932 57918 35941
rect 58530 35935 58586 35944
rect 57610 35930 57616 35932
rect 57672 35930 57696 35932
rect 57752 35930 57776 35932
rect 57832 35930 57856 35932
rect 57912 35930 57918 35932
rect 57672 35878 57674 35930
rect 57854 35878 57856 35930
rect 57610 35876 57616 35878
rect 57672 35876 57696 35878
rect 57752 35876 57776 35878
rect 57832 35876 57856 35878
rect 57912 35876 57918 35878
rect 57610 35867 57918 35876
rect 58532 35488 58584 35494
rect 58532 35430 58584 35436
rect 1950 35388 2258 35397
rect 1950 35386 1956 35388
rect 2012 35386 2036 35388
rect 2092 35386 2116 35388
rect 2172 35386 2196 35388
rect 2252 35386 2258 35388
rect 2012 35334 2014 35386
rect 2194 35334 2196 35386
rect 1950 35332 1956 35334
rect 2012 35332 2036 35334
rect 2092 35332 2116 35334
rect 2172 35332 2196 35334
rect 2252 35332 2258 35334
rect 1950 35323 2258 35332
rect 6950 35388 7258 35397
rect 6950 35386 6956 35388
rect 7012 35386 7036 35388
rect 7092 35386 7116 35388
rect 7172 35386 7196 35388
rect 7252 35386 7258 35388
rect 7012 35334 7014 35386
rect 7194 35334 7196 35386
rect 6950 35332 6956 35334
rect 7012 35332 7036 35334
rect 7092 35332 7116 35334
rect 7172 35332 7196 35334
rect 7252 35332 7258 35334
rect 6950 35323 7258 35332
rect 11950 35388 12258 35397
rect 11950 35386 11956 35388
rect 12012 35386 12036 35388
rect 12092 35386 12116 35388
rect 12172 35386 12196 35388
rect 12252 35386 12258 35388
rect 12012 35334 12014 35386
rect 12194 35334 12196 35386
rect 11950 35332 11956 35334
rect 12012 35332 12036 35334
rect 12092 35332 12116 35334
rect 12172 35332 12196 35334
rect 12252 35332 12258 35334
rect 11950 35323 12258 35332
rect 16950 35388 17258 35397
rect 16950 35386 16956 35388
rect 17012 35386 17036 35388
rect 17092 35386 17116 35388
rect 17172 35386 17196 35388
rect 17252 35386 17258 35388
rect 17012 35334 17014 35386
rect 17194 35334 17196 35386
rect 16950 35332 16956 35334
rect 17012 35332 17036 35334
rect 17092 35332 17116 35334
rect 17172 35332 17196 35334
rect 17252 35332 17258 35334
rect 16950 35323 17258 35332
rect 21950 35388 22258 35397
rect 21950 35386 21956 35388
rect 22012 35386 22036 35388
rect 22092 35386 22116 35388
rect 22172 35386 22196 35388
rect 22252 35386 22258 35388
rect 22012 35334 22014 35386
rect 22194 35334 22196 35386
rect 21950 35332 21956 35334
rect 22012 35332 22036 35334
rect 22092 35332 22116 35334
rect 22172 35332 22196 35334
rect 22252 35332 22258 35334
rect 21950 35323 22258 35332
rect 26950 35388 27258 35397
rect 26950 35386 26956 35388
rect 27012 35386 27036 35388
rect 27092 35386 27116 35388
rect 27172 35386 27196 35388
rect 27252 35386 27258 35388
rect 27012 35334 27014 35386
rect 27194 35334 27196 35386
rect 26950 35332 26956 35334
rect 27012 35332 27036 35334
rect 27092 35332 27116 35334
rect 27172 35332 27196 35334
rect 27252 35332 27258 35334
rect 26950 35323 27258 35332
rect 31950 35388 32258 35397
rect 31950 35386 31956 35388
rect 32012 35386 32036 35388
rect 32092 35386 32116 35388
rect 32172 35386 32196 35388
rect 32252 35386 32258 35388
rect 32012 35334 32014 35386
rect 32194 35334 32196 35386
rect 31950 35332 31956 35334
rect 32012 35332 32036 35334
rect 32092 35332 32116 35334
rect 32172 35332 32196 35334
rect 32252 35332 32258 35334
rect 31950 35323 32258 35332
rect 36950 35388 37258 35397
rect 36950 35386 36956 35388
rect 37012 35386 37036 35388
rect 37092 35386 37116 35388
rect 37172 35386 37196 35388
rect 37252 35386 37258 35388
rect 37012 35334 37014 35386
rect 37194 35334 37196 35386
rect 36950 35332 36956 35334
rect 37012 35332 37036 35334
rect 37092 35332 37116 35334
rect 37172 35332 37196 35334
rect 37252 35332 37258 35334
rect 36950 35323 37258 35332
rect 41950 35388 42258 35397
rect 41950 35386 41956 35388
rect 42012 35386 42036 35388
rect 42092 35386 42116 35388
rect 42172 35386 42196 35388
rect 42252 35386 42258 35388
rect 42012 35334 42014 35386
rect 42194 35334 42196 35386
rect 41950 35332 41956 35334
rect 42012 35332 42036 35334
rect 42092 35332 42116 35334
rect 42172 35332 42196 35334
rect 42252 35332 42258 35334
rect 41950 35323 42258 35332
rect 46950 35388 47258 35397
rect 46950 35386 46956 35388
rect 47012 35386 47036 35388
rect 47092 35386 47116 35388
rect 47172 35386 47196 35388
rect 47252 35386 47258 35388
rect 47012 35334 47014 35386
rect 47194 35334 47196 35386
rect 46950 35332 46956 35334
rect 47012 35332 47036 35334
rect 47092 35332 47116 35334
rect 47172 35332 47196 35334
rect 47252 35332 47258 35334
rect 46950 35323 47258 35332
rect 51950 35388 52258 35397
rect 51950 35386 51956 35388
rect 52012 35386 52036 35388
rect 52092 35386 52116 35388
rect 52172 35386 52196 35388
rect 52252 35386 52258 35388
rect 52012 35334 52014 35386
rect 52194 35334 52196 35386
rect 51950 35332 51956 35334
rect 52012 35332 52036 35334
rect 52092 35332 52116 35334
rect 52172 35332 52196 35334
rect 52252 35332 52258 35334
rect 51950 35323 52258 35332
rect 56950 35388 57258 35397
rect 56950 35386 56956 35388
rect 57012 35386 57036 35388
rect 57092 35386 57116 35388
rect 57172 35386 57196 35388
rect 57252 35386 57258 35388
rect 57012 35334 57014 35386
rect 57194 35334 57196 35386
rect 56950 35332 56956 35334
rect 57012 35332 57036 35334
rect 57092 35332 57116 35334
rect 57172 35332 57196 35334
rect 57252 35332 57258 35334
rect 56950 35323 57258 35332
rect 58544 35193 58572 35430
rect 58530 35184 58586 35193
rect 58530 35119 58586 35128
rect 2610 34844 2918 34853
rect 2610 34842 2616 34844
rect 2672 34842 2696 34844
rect 2752 34842 2776 34844
rect 2832 34842 2856 34844
rect 2912 34842 2918 34844
rect 2672 34790 2674 34842
rect 2854 34790 2856 34842
rect 2610 34788 2616 34790
rect 2672 34788 2696 34790
rect 2752 34788 2776 34790
rect 2832 34788 2856 34790
rect 2912 34788 2918 34790
rect 2610 34779 2918 34788
rect 7610 34844 7918 34853
rect 7610 34842 7616 34844
rect 7672 34842 7696 34844
rect 7752 34842 7776 34844
rect 7832 34842 7856 34844
rect 7912 34842 7918 34844
rect 7672 34790 7674 34842
rect 7854 34790 7856 34842
rect 7610 34788 7616 34790
rect 7672 34788 7696 34790
rect 7752 34788 7776 34790
rect 7832 34788 7856 34790
rect 7912 34788 7918 34790
rect 7610 34779 7918 34788
rect 12610 34844 12918 34853
rect 12610 34842 12616 34844
rect 12672 34842 12696 34844
rect 12752 34842 12776 34844
rect 12832 34842 12856 34844
rect 12912 34842 12918 34844
rect 12672 34790 12674 34842
rect 12854 34790 12856 34842
rect 12610 34788 12616 34790
rect 12672 34788 12696 34790
rect 12752 34788 12776 34790
rect 12832 34788 12856 34790
rect 12912 34788 12918 34790
rect 12610 34779 12918 34788
rect 17610 34844 17918 34853
rect 17610 34842 17616 34844
rect 17672 34842 17696 34844
rect 17752 34842 17776 34844
rect 17832 34842 17856 34844
rect 17912 34842 17918 34844
rect 17672 34790 17674 34842
rect 17854 34790 17856 34842
rect 17610 34788 17616 34790
rect 17672 34788 17696 34790
rect 17752 34788 17776 34790
rect 17832 34788 17856 34790
rect 17912 34788 17918 34790
rect 17610 34779 17918 34788
rect 22610 34844 22918 34853
rect 22610 34842 22616 34844
rect 22672 34842 22696 34844
rect 22752 34842 22776 34844
rect 22832 34842 22856 34844
rect 22912 34842 22918 34844
rect 22672 34790 22674 34842
rect 22854 34790 22856 34842
rect 22610 34788 22616 34790
rect 22672 34788 22696 34790
rect 22752 34788 22776 34790
rect 22832 34788 22856 34790
rect 22912 34788 22918 34790
rect 22610 34779 22918 34788
rect 27610 34844 27918 34853
rect 27610 34842 27616 34844
rect 27672 34842 27696 34844
rect 27752 34842 27776 34844
rect 27832 34842 27856 34844
rect 27912 34842 27918 34844
rect 27672 34790 27674 34842
rect 27854 34790 27856 34842
rect 27610 34788 27616 34790
rect 27672 34788 27696 34790
rect 27752 34788 27776 34790
rect 27832 34788 27856 34790
rect 27912 34788 27918 34790
rect 27610 34779 27918 34788
rect 32610 34844 32918 34853
rect 32610 34842 32616 34844
rect 32672 34842 32696 34844
rect 32752 34842 32776 34844
rect 32832 34842 32856 34844
rect 32912 34842 32918 34844
rect 32672 34790 32674 34842
rect 32854 34790 32856 34842
rect 32610 34788 32616 34790
rect 32672 34788 32696 34790
rect 32752 34788 32776 34790
rect 32832 34788 32856 34790
rect 32912 34788 32918 34790
rect 32610 34779 32918 34788
rect 37610 34844 37918 34853
rect 37610 34842 37616 34844
rect 37672 34842 37696 34844
rect 37752 34842 37776 34844
rect 37832 34842 37856 34844
rect 37912 34842 37918 34844
rect 37672 34790 37674 34842
rect 37854 34790 37856 34842
rect 37610 34788 37616 34790
rect 37672 34788 37696 34790
rect 37752 34788 37776 34790
rect 37832 34788 37856 34790
rect 37912 34788 37918 34790
rect 37610 34779 37918 34788
rect 42610 34844 42918 34853
rect 42610 34842 42616 34844
rect 42672 34842 42696 34844
rect 42752 34842 42776 34844
rect 42832 34842 42856 34844
rect 42912 34842 42918 34844
rect 42672 34790 42674 34842
rect 42854 34790 42856 34842
rect 42610 34788 42616 34790
rect 42672 34788 42696 34790
rect 42752 34788 42776 34790
rect 42832 34788 42856 34790
rect 42912 34788 42918 34790
rect 42610 34779 42918 34788
rect 47610 34844 47918 34853
rect 47610 34842 47616 34844
rect 47672 34842 47696 34844
rect 47752 34842 47776 34844
rect 47832 34842 47856 34844
rect 47912 34842 47918 34844
rect 47672 34790 47674 34842
rect 47854 34790 47856 34842
rect 47610 34788 47616 34790
rect 47672 34788 47696 34790
rect 47752 34788 47776 34790
rect 47832 34788 47856 34790
rect 47912 34788 47918 34790
rect 47610 34779 47918 34788
rect 52610 34844 52918 34853
rect 52610 34842 52616 34844
rect 52672 34842 52696 34844
rect 52752 34842 52776 34844
rect 52832 34842 52856 34844
rect 52912 34842 52918 34844
rect 52672 34790 52674 34842
rect 52854 34790 52856 34842
rect 52610 34788 52616 34790
rect 52672 34788 52696 34790
rect 52752 34788 52776 34790
rect 52832 34788 52856 34790
rect 52912 34788 52918 34790
rect 52610 34779 52918 34788
rect 57610 34844 57918 34853
rect 57610 34842 57616 34844
rect 57672 34842 57696 34844
rect 57752 34842 57776 34844
rect 57832 34842 57856 34844
rect 57912 34842 57918 34844
rect 57672 34790 57674 34842
rect 57854 34790 57856 34842
rect 57610 34788 57616 34790
rect 57672 34788 57696 34790
rect 57752 34788 57776 34790
rect 57832 34788 57856 34790
rect 57912 34788 57918 34790
rect 57610 34779 57918 34788
rect 58532 34400 58584 34406
rect 58530 34368 58532 34377
rect 58584 34368 58586 34377
rect 1950 34300 2258 34309
rect 1950 34298 1956 34300
rect 2012 34298 2036 34300
rect 2092 34298 2116 34300
rect 2172 34298 2196 34300
rect 2252 34298 2258 34300
rect 2012 34246 2014 34298
rect 2194 34246 2196 34298
rect 1950 34244 1956 34246
rect 2012 34244 2036 34246
rect 2092 34244 2116 34246
rect 2172 34244 2196 34246
rect 2252 34244 2258 34246
rect 1950 34235 2258 34244
rect 6950 34300 7258 34309
rect 6950 34298 6956 34300
rect 7012 34298 7036 34300
rect 7092 34298 7116 34300
rect 7172 34298 7196 34300
rect 7252 34298 7258 34300
rect 7012 34246 7014 34298
rect 7194 34246 7196 34298
rect 6950 34244 6956 34246
rect 7012 34244 7036 34246
rect 7092 34244 7116 34246
rect 7172 34244 7196 34246
rect 7252 34244 7258 34246
rect 6950 34235 7258 34244
rect 11950 34300 12258 34309
rect 11950 34298 11956 34300
rect 12012 34298 12036 34300
rect 12092 34298 12116 34300
rect 12172 34298 12196 34300
rect 12252 34298 12258 34300
rect 12012 34246 12014 34298
rect 12194 34246 12196 34298
rect 11950 34244 11956 34246
rect 12012 34244 12036 34246
rect 12092 34244 12116 34246
rect 12172 34244 12196 34246
rect 12252 34244 12258 34246
rect 11950 34235 12258 34244
rect 16950 34300 17258 34309
rect 16950 34298 16956 34300
rect 17012 34298 17036 34300
rect 17092 34298 17116 34300
rect 17172 34298 17196 34300
rect 17252 34298 17258 34300
rect 17012 34246 17014 34298
rect 17194 34246 17196 34298
rect 16950 34244 16956 34246
rect 17012 34244 17036 34246
rect 17092 34244 17116 34246
rect 17172 34244 17196 34246
rect 17252 34244 17258 34246
rect 16950 34235 17258 34244
rect 21950 34300 22258 34309
rect 21950 34298 21956 34300
rect 22012 34298 22036 34300
rect 22092 34298 22116 34300
rect 22172 34298 22196 34300
rect 22252 34298 22258 34300
rect 22012 34246 22014 34298
rect 22194 34246 22196 34298
rect 21950 34244 21956 34246
rect 22012 34244 22036 34246
rect 22092 34244 22116 34246
rect 22172 34244 22196 34246
rect 22252 34244 22258 34246
rect 21950 34235 22258 34244
rect 26950 34300 27258 34309
rect 26950 34298 26956 34300
rect 27012 34298 27036 34300
rect 27092 34298 27116 34300
rect 27172 34298 27196 34300
rect 27252 34298 27258 34300
rect 27012 34246 27014 34298
rect 27194 34246 27196 34298
rect 26950 34244 26956 34246
rect 27012 34244 27036 34246
rect 27092 34244 27116 34246
rect 27172 34244 27196 34246
rect 27252 34244 27258 34246
rect 26950 34235 27258 34244
rect 31950 34300 32258 34309
rect 31950 34298 31956 34300
rect 32012 34298 32036 34300
rect 32092 34298 32116 34300
rect 32172 34298 32196 34300
rect 32252 34298 32258 34300
rect 32012 34246 32014 34298
rect 32194 34246 32196 34298
rect 31950 34244 31956 34246
rect 32012 34244 32036 34246
rect 32092 34244 32116 34246
rect 32172 34244 32196 34246
rect 32252 34244 32258 34246
rect 31950 34235 32258 34244
rect 36950 34300 37258 34309
rect 36950 34298 36956 34300
rect 37012 34298 37036 34300
rect 37092 34298 37116 34300
rect 37172 34298 37196 34300
rect 37252 34298 37258 34300
rect 37012 34246 37014 34298
rect 37194 34246 37196 34298
rect 36950 34244 36956 34246
rect 37012 34244 37036 34246
rect 37092 34244 37116 34246
rect 37172 34244 37196 34246
rect 37252 34244 37258 34246
rect 36950 34235 37258 34244
rect 41950 34300 42258 34309
rect 41950 34298 41956 34300
rect 42012 34298 42036 34300
rect 42092 34298 42116 34300
rect 42172 34298 42196 34300
rect 42252 34298 42258 34300
rect 42012 34246 42014 34298
rect 42194 34246 42196 34298
rect 41950 34244 41956 34246
rect 42012 34244 42036 34246
rect 42092 34244 42116 34246
rect 42172 34244 42196 34246
rect 42252 34244 42258 34246
rect 41950 34235 42258 34244
rect 46950 34300 47258 34309
rect 46950 34298 46956 34300
rect 47012 34298 47036 34300
rect 47092 34298 47116 34300
rect 47172 34298 47196 34300
rect 47252 34298 47258 34300
rect 47012 34246 47014 34298
rect 47194 34246 47196 34298
rect 46950 34244 46956 34246
rect 47012 34244 47036 34246
rect 47092 34244 47116 34246
rect 47172 34244 47196 34246
rect 47252 34244 47258 34246
rect 46950 34235 47258 34244
rect 51950 34300 52258 34309
rect 51950 34298 51956 34300
rect 52012 34298 52036 34300
rect 52092 34298 52116 34300
rect 52172 34298 52196 34300
rect 52252 34298 52258 34300
rect 52012 34246 52014 34298
rect 52194 34246 52196 34298
rect 51950 34244 51956 34246
rect 52012 34244 52036 34246
rect 52092 34244 52116 34246
rect 52172 34244 52196 34246
rect 52252 34244 52258 34246
rect 51950 34235 52258 34244
rect 56950 34300 57258 34309
rect 58530 34303 58586 34312
rect 56950 34298 56956 34300
rect 57012 34298 57036 34300
rect 57092 34298 57116 34300
rect 57172 34298 57196 34300
rect 57252 34298 57258 34300
rect 57012 34246 57014 34298
rect 57194 34246 57196 34298
rect 56950 34244 56956 34246
rect 57012 34244 57036 34246
rect 57092 34244 57116 34246
rect 57172 34244 57196 34246
rect 57252 34244 57258 34246
rect 56950 34235 57258 34244
rect 58532 33992 58584 33998
rect 58532 33934 58584 33940
rect 2610 33756 2918 33765
rect 2610 33754 2616 33756
rect 2672 33754 2696 33756
rect 2752 33754 2776 33756
rect 2832 33754 2856 33756
rect 2912 33754 2918 33756
rect 2672 33702 2674 33754
rect 2854 33702 2856 33754
rect 2610 33700 2616 33702
rect 2672 33700 2696 33702
rect 2752 33700 2776 33702
rect 2832 33700 2856 33702
rect 2912 33700 2918 33702
rect 2610 33691 2918 33700
rect 7610 33756 7918 33765
rect 7610 33754 7616 33756
rect 7672 33754 7696 33756
rect 7752 33754 7776 33756
rect 7832 33754 7856 33756
rect 7912 33754 7918 33756
rect 7672 33702 7674 33754
rect 7854 33702 7856 33754
rect 7610 33700 7616 33702
rect 7672 33700 7696 33702
rect 7752 33700 7776 33702
rect 7832 33700 7856 33702
rect 7912 33700 7918 33702
rect 7610 33691 7918 33700
rect 12610 33756 12918 33765
rect 12610 33754 12616 33756
rect 12672 33754 12696 33756
rect 12752 33754 12776 33756
rect 12832 33754 12856 33756
rect 12912 33754 12918 33756
rect 12672 33702 12674 33754
rect 12854 33702 12856 33754
rect 12610 33700 12616 33702
rect 12672 33700 12696 33702
rect 12752 33700 12776 33702
rect 12832 33700 12856 33702
rect 12912 33700 12918 33702
rect 12610 33691 12918 33700
rect 17610 33756 17918 33765
rect 17610 33754 17616 33756
rect 17672 33754 17696 33756
rect 17752 33754 17776 33756
rect 17832 33754 17856 33756
rect 17912 33754 17918 33756
rect 17672 33702 17674 33754
rect 17854 33702 17856 33754
rect 17610 33700 17616 33702
rect 17672 33700 17696 33702
rect 17752 33700 17776 33702
rect 17832 33700 17856 33702
rect 17912 33700 17918 33702
rect 17610 33691 17918 33700
rect 22610 33756 22918 33765
rect 22610 33754 22616 33756
rect 22672 33754 22696 33756
rect 22752 33754 22776 33756
rect 22832 33754 22856 33756
rect 22912 33754 22918 33756
rect 22672 33702 22674 33754
rect 22854 33702 22856 33754
rect 22610 33700 22616 33702
rect 22672 33700 22696 33702
rect 22752 33700 22776 33702
rect 22832 33700 22856 33702
rect 22912 33700 22918 33702
rect 22610 33691 22918 33700
rect 27610 33756 27918 33765
rect 27610 33754 27616 33756
rect 27672 33754 27696 33756
rect 27752 33754 27776 33756
rect 27832 33754 27856 33756
rect 27912 33754 27918 33756
rect 27672 33702 27674 33754
rect 27854 33702 27856 33754
rect 27610 33700 27616 33702
rect 27672 33700 27696 33702
rect 27752 33700 27776 33702
rect 27832 33700 27856 33702
rect 27912 33700 27918 33702
rect 27610 33691 27918 33700
rect 32610 33756 32918 33765
rect 32610 33754 32616 33756
rect 32672 33754 32696 33756
rect 32752 33754 32776 33756
rect 32832 33754 32856 33756
rect 32912 33754 32918 33756
rect 32672 33702 32674 33754
rect 32854 33702 32856 33754
rect 32610 33700 32616 33702
rect 32672 33700 32696 33702
rect 32752 33700 32776 33702
rect 32832 33700 32856 33702
rect 32912 33700 32918 33702
rect 32610 33691 32918 33700
rect 37610 33756 37918 33765
rect 37610 33754 37616 33756
rect 37672 33754 37696 33756
rect 37752 33754 37776 33756
rect 37832 33754 37856 33756
rect 37912 33754 37918 33756
rect 37672 33702 37674 33754
rect 37854 33702 37856 33754
rect 37610 33700 37616 33702
rect 37672 33700 37696 33702
rect 37752 33700 37776 33702
rect 37832 33700 37856 33702
rect 37912 33700 37918 33702
rect 37610 33691 37918 33700
rect 42610 33756 42918 33765
rect 42610 33754 42616 33756
rect 42672 33754 42696 33756
rect 42752 33754 42776 33756
rect 42832 33754 42856 33756
rect 42912 33754 42918 33756
rect 42672 33702 42674 33754
rect 42854 33702 42856 33754
rect 42610 33700 42616 33702
rect 42672 33700 42696 33702
rect 42752 33700 42776 33702
rect 42832 33700 42856 33702
rect 42912 33700 42918 33702
rect 42610 33691 42918 33700
rect 47610 33756 47918 33765
rect 47610 33754 47616 33756
rect 47672 33754 47696 33756
rect 47752 33754 47776 33756
rect 47832 33754 47856 33756
rect 47912 33754 47918 33756
rect 47672 33702 47674 33754
rect 47854 33702 47856 33754
rect 47610 33700 47616 33702
rect 47672 33700 47696 33702
rect 47752 33700 47776 33702
rect 47832 33700 47856 33702
rect 47912 33700 47918 33702
rect 47610 33691 47918 33700
rect 52610 33756 52918 33765
rect 52610 33754 52616 33756
rect 52672 33754 52696 33756
rect 52752 33754 52776 33756
rect 52832 33754 52856 33756
rect 52912 33754 52918 33756
rect 52672 33702 52674 33754
rect 52854 33702 52856 33754
rect 52610 33700 52616 33702
rect 52672 33700 52696 33702
rect 52752 33700 52776 33702
rect 52832 33700 52856 33702
rect 52912 33700 52918 33702
rect 52610 33691 52918 33700
rect 57610 33756 57918 33765
rect 57610 33754 57616 33756
rect 57672 33754 57696 33756
rect 57752 33754 57776 33756
rect 57832 33754 57856 33756
rect 57912 33754 57918 33756
rect 57672 33702 57674 33754
rect 57854 33702 57856 33754
rect 57610 33700 57616 33702
rect 57672 33700 57696 33702
rect 57752 33700 57776 33702
rect 57832 33700 57856 33702
rect 57912 33700 57918 33702
rect 57610 33691 57918 33700
rect 58544 33561 58572 33934
rect 58530 33552 58586 33561
rect 58530 33487 58586 33496
rect 1950 33212 2258 33221
rect 1950 33210 1956 33212
rect 2012 33210 2036 33212
rect 2092 33210 2116 33212
rect 2172 33210 2196 33212
rect 2252 33210 2258 33212
rect 2012 33158 2014 33210
rect 2194 33158 2196 33210
rect 1950 33156 1956 33158
rect 2012 33156 2036 33158
rect 2092 33156 2116 33158
rect 2172 33156 2196 33158
rect 2252 33156 2258 33158
rect 1950 33147 2258 33156
rect 6950 33212 7258 33221
rect 6950 33210 6956 33212
rect 7012 33210 7036 33212
rect 7092 33210 7116 33212
rect 7172 33210 7196 33212
rect 7252 33210 7258 33212
rect 7012 33158 7014 33210
rect 7194 33158 7196 33210
rect 6950 33156 6956 33158
rect 7012 33156 7036 33158
rect 7092 33156 7116 33158
rect 7172 33156 7196 33158
rect 7252 33156 7258 33158
rect 6950 33147 7258 33156
rect 11950 33212 12258 33221
rect 11950 33210 11956 33212
rect 12012 33210 12036 33212
rect 12092 33210 12116 33212
rect 12172 33210 12196 33212
rect 12252 33210 12258 33212
rect 12012 33158 12014 33210
rect 12194 33158 12196 33210
rect 11950 33156 11956 33158
rect 12012 33156 12036 33158
rect 12092 33156 12116 33158
rect 12172 33156 12196 33158
rect 12252 33156 12258 33158
rect 11950 33147 12258 33156
rect 16950 33212 17258 33221
rect 16950 33210 16956 33212
rect 17012 33210 17036 33212
rect 17092 33210 17116 33212
rect 17172 33210 17196 33212
rect 17252 33210 17258 33212
rect 17012 33158 17014 33210
rect 17194 33158 17196 33210
rect 16950 33156 16956 33158
rect 17012 33156 17036 33158
rect 17092 33156 17116 33158
rect 17172 33156 17196 33158
rect 17252 33156 17258 33158
rect 16950 33147 17258 33156
rect 21950 33212 22258 33221
rect 21950 33210 21956 33212
rect 22012 33210 22036 33212
rect 22092 33210 22116 33212
rect 22172 33210 22196 33212
rect 22252 33210 22258 33212
rect 22012 33158 22014 33210
rect 22194 33158 22196 33210
rect 21950 33156 21956 33158
rect 22012 33156 22036 33158
rect 22092 33156 22116 33158
rect 22172 33156 22196 33158
rect 22252 33156 22258 33158
rect 21950 33147 22258 33156
rect 26950 33212 27258 33221
rect 26950 33210 26956 33212
rect 27012 33210 27036 33212
rect 27092 33210 27116 33212
rect 27172 33210 27196 33212
rect 27252 33210 27258 33212
rect 27012 33158 27014 33210
rect 27194 33158 27196 33210
rect 26950 33156 26956 33158
rect 27012 33156 27036 33158
rect 27092 33156 27116 33158
rect 27172 33156 27196 33158
rect 27252 33156 27258 33158
rect 26950 33147 27258 33156
rect 31950 33212 32258 33221
rect 31950 33210 31956 33212
rect 32012 33210 32036 33212
rect 32092 33210 32116 33212
rect 32172 33210 32196 33212
rect 32252 33210 32258 33212
rect 32012 33158 32014 33210
rect 32194 33158 32196 33210
rect 31950 33156 31956 33158
rect 32012 33156 32036 33158
rect 32092 33156 32116 33158
rect 32172 33156 32196 33158
rect 32252 33156 32258 33158
rect 31950 33147 32258 33156
rect 36950 33212 37258 33221
rect 36950 33210 36956 33212
rect 37012 33210 37036 33212
rect 37092 33210 37116 33212
rect 37172 33210 37196 33212
rect 37252 33210 37258 33212
rect 37012 33158 37014 33210
rect 37194 33158 37196 33210
rect 36950 33156 36956 33158
rect 37012 33156 37036 33158
rect 37092 33156 37116 33158
rect 37172 33156 37196 33158
rect 37252 33156 37258 33158
rect 36950 33147 37258 33156
rect 41950 33212 42258 33221
rect 41950 33210 41956 33212
rect 42012 33210 42036 33212
rect 42092 33210 42116 33212
rect 42172 33210 42196 33212
rect 42252 33210 42258 33212
rect 42012 33158 42014 33210
rect 42194 33158 42196 33210
rect 41950 33156 41956 33158
rect 42012 33156 42036 33158
rect 42092 33156 42116 33158
rect 42172 33156 42196 33158
rect 42252 33156 42258 33158
rect 41950 33147 42258 33156
rect 46950 33212 47258 33221
rect 46950 33210 46956 33212
rect 47012 33210 47036 33212
rect 47092 33210 47116 33212
rect 47172 33210 47196 33212
rect 47252 33210 47258 33212
rect 47012 33158 47014 33210
rect 47194 33158 47196 33210
rect 46950 33156 46956 33158
rect 47012 33156 47036 33158
rect 47092 33156 47116 33158
rect 47172 33156 47196 33158
rect 47252 33156 47258 33158
rect 46950 33147 47258 33156
rect 51950 33212 52258 33221
rect 51950 33210 51956 33212
rect 52012 33210 52036 33212
rect 52092 33210 52116 33212
rect 52172 33210 52196 33212
rect 52252 33210 52258 33212
rect 52012 33158 52014 33210
rect 52194 33158 52196 33210
rect 51950 33156 51956 33158
rect 52012 33156 52036 33158
rect 52092 33156 52116 33158
rect 52172 33156 52196 33158
rect 52252 33156 52258 33158
rect 51950 33147 52258 33156
rect 56950 33212 57258 33221
rect 56950 33210 56956 33212
rect 57012 33210 57036 33212
rect 57092 33210 57116 33212
rect 57172 33210 57196 33212
rect 57252 33210 57258 33212
rect 57012 33158 57014 33210
rect 57194 33158 57196 33210
rect 56950 33156 56956 33158
rect 57012 33156 57036 33158
rect 57092 33156 57116 33158
rect 57172 33156 57196 33158
rect 57252 33156 57258 33158
rect 56950 33147 57258 33156
rect 58532 32904 58584 32910
rect 58532 32846 58584 32852
rect 58544 32745 58572 32846
rect 58530 32736 58586 32745
rect 2610 32668 2918 32677
rect 2610 32666 2616 32668
rect 2672 32666 2696 32668
rect 2752 32666 2776 32668
rect 2832 32666 2856 32668
rect 2912 32666 2918 32668
rect 2672 32614 2674 32666
rect 2854 32614 2856 32666
rect 2610 32612 2616 32614
rect 2672 32612 2696 32614
rect 2752 32612 2776 32614
rect 2832 32612 2856 32614
rect 2912 32612 2918 32614
rect 2610 32603 2918 32612
rect 7610 32668 7918 32677
rect 7610 32666 7616 32668
rect 7672 32666 7696 32668
rect 7752 32666 7776 32668
rect 7832 32666 7856 32668
rect 7912 32666 7918 32668
rect 7672 32614 7674 32666
rect 7854 32614 7856 32666
rect 7610 32612 7616 32614
rect 7672 32612 7696 32614
rect 7752 32612 7776 32614
rect 7832 32612 7856 32614
rect 7912 32612 7918 32614
rect 7610 32603 7918 32612
rect 12610 32668 12918 32677
rect 12610 32666 12616 32668
rect 12672 32666 12696 32668
rect 12752 32666 12776 32668
rect 12832 32666 12856 32668
rect 12912 32666 12918 32668
rect 12672 32614 12674 32666
rect 12854 32614 12856 32666
rect 12610 32612 12616 32614
rect 12672 32612 12696 32614
rect 12752 32612 12776 32614
rect 12832 32612 12856 32614
rect 12912 32612 12918 32614
rect 12610 32603 12918 32612
rect 17610 32668 17918 32677
rect 17610 32666 17616 32668
rect 17672 32666 17696 32668
rect 17752 32666 17776 32668
rect 17832 32666 17856 32668
rect 17912 32666 17918 32668
rect 17672 32614 17674 32666
rect 17854 32614 17856 32666
rect 17610 32612 17616 32614
rect 17672 32612 17696 32614
rect 17752 32612 17776 32614
rect 17832 32612 17856 32614
rect 17912 32612 17918 32614
rect 17610 32603 17918 32612
rect 22610 32668 22918 32677
rect 22610 32666 22616 32668
rect 22672 32666 22696 32668
rect 22752 32666 22776 32668
rect 22832 32666 22856 32668
rect 22912 32666 22918 32668
rect 22672 32614 22674 32666
rect 22854 32614 22856 32666
rect 22610 32612 22616 32614
rect 22672 32612 22696 32614
rect 22752 32612 22776 32614
rect 22832 32612 22856 32614
rect 22912 32612 22918 32614
rect 22610 32603 22918 32612
rect 27610 32668 27918 32677
rect 27610 32666 27616 32668
rect 27672 32666 27696 32668
rect 27752 32666 27776 32668
rect 27832 32666 27856 32668
rect 27912 32666 27918 32668
rect 27672 32614 27674 32666
rect 27854 32614 27856 32666
rect 27610 32612 27616 32614
rect 27672 32612 27696 32614
rect 27752 32612 27776 32614
rect 27832 32612 27856 32614
rect 27912 32612 27918 32614
rect 27610 32603 27918 32612
rect 32610 32668 32918 32677
rect 32610 32666 32616 32668
rect 32672 32666 32696 32668
rect 32752 32666 32776 32668
rect 32832 32666 32856 32668
rect 32912 32666 32918 32668
rect 32672 32614 32674 32666
rect 32854 32614 32856 32666
rect 32610 32612 32616 32614
rect 32672 32612 32696 32614
rect 32752 32612 32776 32614
rect 32832 32612 32856 32614
rect 32912 32612 32918 32614
rect 32610 32603 32918 32612
rect 37610 32668 37918 32677
rect 37610 32666 37616 32668
rect 37672 32666 37696 32668
rect 37752 32666 37776 32668
rect 37832 32666 37856 32668
rect 37912 32666 37918 32668
rect 37672 32614 37674 32666
rect 37854 32614 37856 32666
rect 37610 32612 37616 32614
rect 37672 32612 37696 32614
rect 37752 32612 37776 32614
rect 37832 32612 37856 32614
rect 37912 32612 37918 32614
rect 37610 32603 37918 32612
rect 42610 32668 42918 32677
rect 42610 32666 42616 32668
rect 42672 32666 42696 32668
rect 42752 32666 42776 32668
rect 42832 32666 42856 32668
rect 42912 32666 42918 32668
rect 42672 32614 42674 32666
rect 42854 32614 42856 32666
rect 42610 32612 42616 32614
rect 42672 32612 42696 32614
rect 42752 32612 42776 32614
rect 42832 32612 42856 32614
rect 42912 32612 42918 32614
rect 42610 32603 42918 32612
rect 47610 32668 47918 32677
rect 47610 32666 47616 32668
rect 47672 32666 47696 32668
rect 47752 32666 47776 32668
rect 47832 32666 47856 32668
rect 47912 32666 47918 32668
rect 47672 32614 47674 32666
rect 47854 32614 47856 32666
rect 47610 32612 47616 32614
rect 47672 32612 47696 32614
rect 47752 32612 47776 32614
rect 47832 32612 47856 32614
rect 47912 32612 47918 32614
rect 47610 32603 47918 32612
rect 52610 32668 52918 32677
rect 52610 32666 52616 32668
rect 52672 32666 52696 32668
rect 52752 32666 52776 32668
rect 52832 32666 52856 32668
rect 52912 32666 52918 32668
rect 52672 32614 52674 32666
rect 52854 32614 52856 32666
rect 52610 32612 52616 32614
rect 52672 32612 52696 32614
rect 52752 32612 52776 32614
rect 52832 32612 52856 32614
rect 52912 32612 52918 32614
rect 52610 32603 52918 32612
rect 57610 32668 57918 32677
rect 58530 32671 58586 32680
rect 57610 32666 57616 32668
rect 57672 32666 57696 32668
rect 57752 32666 57776 32668
rect 57832 32666 57856 32668
rect 57912 32666 57918 32668
rect 57672 32614 57674 32666
rect 57854 32614 57856 32666
rect 57610 32612 57616 32614
rect 57672 32612 57696 32614
rect 57752 32612 57776 32614
rect 57832 32612 57856 32614
rect 57912 32612 57918 32614
rect 57610 32603 57918 32612
rect 58532 32224 58584 32230
rect 58532 32166 58584 32172
rect 1950 32124 2258 32133
rect 1950 32122 1956 32124
rect 2012 32122 2036 32124
rect 2092 32122 2116 32124
rect 2172 32122 2196 32124
rect 2252 32122 2258 32124
rect 2012 32070 2014 32122
rect 2194 32070 2196 32122
rect 1950 32068 1956 32070
rect 2012 32068 2036 32070
rect 2092 32068 2116 32070
rect 2172 32068 2196 32070
rect 2252 32068 2258 32070
rect 1950 32059 2258 32068
rect 6950 32124 7258 32133
rect 6950 32122 6956 32124
rect 7012 32122 7036 32124
rect 7092 32122 7116 32124
rect 7172 32122 7196 32124
rect 7252 32122 7258 32124
rect 7012 32070 7014 32122
rect 7194 32070 7196 32122
rect 6950 32068 6956 32070
rect 7012 32068 7036 32070
rect 7092 32068 7116 32070
rect 7172 32068 7196 32070
rect 7252 32068 7258 32070
rect 6950 32059 7258 32068
rect 11950 32124 12258 32133
rect 11950 32122 11956 32124
rect 12012 32122 12036 32124
rect 12092 32122 12116 32124
rect 12172 32122 12196 32124
rect 12252 32122 12258 32124
rect 12012 32070 12014 32122
rect 12194 32070 12196 32122
rect 11950 32068 11956 32070
rect 12012 32068 12036 32070
rect 12092 32068 12116 32070
rect 12172 32068 12196 32070
rect 12252 32068 12258 32070
rect 11950 32059 12258 32068
rect 16950 32124 17258 32133
rect 16950 32122 16956 32124
rect 17012 32122 17036 32124
rect 17092 32122 17116 32124
rect 17172 32122 17196 32124
rect 17252 32122 17258 32124
rect 17012 32070 17014 32122
rect 17194 32070 17196 32122
rect 16950 32068 16956 32070
rect 17012 32068 17036 32070
rect 17092 32068 17116 32070
rect 17172 32068 17196 32070
rect 17252 32068 17258 32070
rect 16950 32059 17258 32068
rect 21950 32124 22258 32133
rect 21950 32122 21956 32124
rect 22012 32122 22036 32124
rect 22092 32122 22116 32124
rect 22172 32122 22196 32124
rect 22252 32122 22258 32124
rect 22012 32070 22014 32122
rect 22194 32070 22196 32122
rect 21950 32068 21956 32070
rect 22012 32068 22036 32070
rect 22092 32068 22116 32070
rect 22172 32068 22196 32070
rect 22252 32068 22258 32070
rect 21950 32059 22258 32068
rect 26950 32124 27258 32133
rect 26950 32122 26956 32124
rect 27012 32122 27036 32124
rect 27092 32122 27116 32124
rect 27172 32122 27196 32124
rect 27252 32122 27258 32124
rect 27012 32070 27014 32122
rect 27194 32070 27196 32122
rect 26950 32068 26956 32070
rect 27012 32068 27036 32070
rect 27092 32068 27116 32070
rect 27172 32068 27196 32070
rect 27252 32068 27258 32070
rect 26950 32059 27258 32068
rect 31950 32124 32258 32133
rect 31950 32122 31956 32124
rect 32012 32122 32036 32124
rect 32092 32122 32116 32124
rect 32172 32122 32196 32124
rect 32252 32122 32258 32124
rect 32012 32070 32014 32122
rect 32194 32070 32196 32122
rect 31950 32068 31956 32070
rect 32012 32068 32036 32070
rect 32092 32068 32116 32070
rect 32172 32068 32196 32070
rect 32252 32068 32258 32070
rect 31950 32059 32258 32068
rect 36950 32124 37258 32133
rect 36950 32122 36956 32124
rect 37012 32122 37036 32124
rect 37092 32122 37116 32124
rect 37172 32122 37196 32124
rect 37252 32122 37258 32124
rect 37012 32070 37014 32122
rect 37194 32070 37196 32122
rect 36950 32068 36956 32070
rect 37012 32068 37036 32070
rect 37092 32068 37116 32070
rect 37172 32068 37196 32070
rect 37252 32068 37258 32070
rect 36950 32059 37258 32068
rect 41950 32124 42258 32133
rect 41950 32122 41956 32124
rect 42012 32122 42036 32124
rect 42092 32122 42116 32124
rect 42172 32122 42196 32124
rect 42252 32122 42258 32124
rect 42012 32070 42014 32122
rect 42194 32070 42196 32122
rect 41950 32068 41956 32070
rect 42012 32068 42036 32070
rect 42092 32068 42116 32070
rect 42172 32068 42196 32070
rect 42252 32068 42258 32070
rect 41950 32059 42258 32068
rect 46950 32124 47258 32133
rect 46950 32122 46956 32124
rect 47012 32122 47036 32124
rect 47092 32122 47116 32124
rect 47172 32122 47196 32124
rect 47252 32122 47258 32124
rect 47012 32070 47014 32122
rect 47194 32070 47196 32122
rect 46950 32068 46956 32070
rect 47012 32068 47036 32070
rect 47092 32068 47116 32070
rect 47172 32068 47196 32070
rect 47252 32068 47258 32070
rect 46950 32059 47258 32068
rect 51950 32124 52258 32133
rect 51950 32122 51956 32124
rect 52012 32122 52036 32124
rect 52092 32122 52116 32124
rect 52172 32122 52196 32124
rect 52252 32122 52258 32124
rect 52012 32070 52014 32122
rect 52194 32070 52196 32122
rect 51950 32068 51956 32070
rect 52012 32068 52036 32070
rect 52092 32068 52116 32070
rect 52172 32068 52196 32070
rect 52252 32068 52258 32070
rect 51950 32059 52258 32068
rect 56950 32124 57258 32133
rect 56950 32122 56956 32124
rect 57012 32122 57036 32124
rect 57092 32122 57116 32124
rect 57172 32122 57196 32124
rect 57252 32122 57258 32124
rect 57012 32070 57014 32122
rect 57194 32070 57196 32122
rect 56950 32068 56956 32070
rect 57012 32068 57036 32070
rect 57092 32068 57116 32070
rect 57172 32068 57196 32070
rect 57252 32068 57258 32070
rect 56950 32059 57258 32068
rect 58544 31929 58572 32166
rect 58530 31920 58586 31929
rect 58530 31855 58586 31864
rect 2610 31580 2918 31589
rect 2610 31578 2616 31580
rect 2672 31578 2696 31580
rect 2752 31578 2776 31580
rect 2832 31578 2856 31580
rect 2912 31578 2918 31580
rect 2672 31526 2674 31578
rect 2854 31526 2856 31578
rect 2610 31524 2616 31526
rect 2672 31524 2696 31526
rect 2752 31524 2776 31526
rect 2832 31524 2856 31526
rect 2912 31524 2918 31526
rect 2610 31515 2918 31524
rect 7610 31580 7918 31589
rect 7610 31578 7616 31580
rect 7672 31578 7696 31580
rect 7752 31578 7776 31580
rect 7832 31578 7856 31580
rect 7912 31578 7918 31580
rect 7672 31526 7674 31578
rect 7854 31526 7856 31578
rect 7610 31524 7616 31526
rect 7672 31524 7696 31526
rect 7752 31524 7776 31526
rect 7832 31524 7856 31526
rect 7912 31524 7918 31526
rect 7610 31515 7918 31524
rect 12610 31580 12918 31589
rect 12610 31578 12616 31580
rect 12672 31578 12696 31580
rect 12752 31578 12776 31580
rect 12832 31578 12856 31580
rect 12912 31578 12918 31580
rect 12672 31526 12674 31578
rect 12854 31526 12856 31578
rect 12610 31524 12616 31526
rect 12672 31524 12696 31526
rect 12752 31524 12776 31526
rect 12832 31524 12856 31526
rect 12912 31524 12918 31526
rect 12610 31515 12918 31524
rect 17610 31580 17918 31589
rect 17610 31578 17616 31580
rect 17672 31578 17696 31580
rect 17752 31578 17776 31580
rect 17832 31578 17856 31580
rect 17912 31578 17918 31580
rect 17672 31526 17674 31578
rect 17854 31526 17856 31578
rect 17610 31524 17616 31526
rect 17672 31524 17696 31526
rect 17752 31524 17776 31526
rect 17832 31524 17856 31526
rect 17912 31524 17918 31526
rect 17610 31515 17918 31524
rect 22610 31580 22918 31589
rect 22610 31578 22616 31580
rect 22672 31578 22696 31580
rect 22752 31578 22776 31580
rect 22832 31578 22856 31580
rect 22912 31578 22918 31580
rect 22672 31526 22674 31578
rect 22854 31526 22856 31578
rect 22610 31524 22616 31526
rect 22672 31524 22696 31526
rect 22752 31524 22776 31526
rect 22832 31524 22856 31526
rect 22912 31524 22918 31526
rect 22610 31515 22918 31524
rect 27610 31580 27918 31589
rect 27610 31578 27616 31580
rect 27672 31578 27696 31580
rect 27752 31578 27776 31580
rect 27832 31578 27856 31580
rect 27912 31578 27918 31580
rect 27672 31526 27674 31578
rect 27854 31526 27856 31578
rect 27610 31524 27616 31526
rect 27672 31524 27696 31526
rect 27752 31524 27776 31526
rect 27832 31524 27856 31526
rect 27912 31524 27918 31526
rect 27610 31515 27918 31524
rect 32610 31580 32918 31589
rect 32610 31578 32616 31580
rect 32672 31578 32696 31580
rect 32752 31578 32776 31580
rect 32832 31578 32856 31580
rect 32912 31578 32918 31580
rect 32672 31526 32674 31578
rect 32854 31526 32856 31578
rect 32610 31524 32616 31526
rect 32672 31524 32696 31526
rect 32752 31524 32776 31526
rect 32832 31524 32856 31526
rect 32912 31524 32918 31526
rect 32610 31515 32918 31524
rect 37610 31580 37918 31589
rect 37610 31578 37616 31580
rect 37672 31578 37696 31580
rect 37752 31578 37776 31580
rect 37832 31578 37856 31580
rect 37912 31578 37918 31580
rect 37672 31526 37674 31578
rect 37854 31526 37856 31578
rect 37610 31524 37616 31526
rect 37672 31524 37696 31526
rect 37752 31524 37776 31526
rect 37832 31524 37856 31526
rect 37912 31524 37918 31526
rect 37610 31515 37918 31524
rect 42610 31580 42918 31589
rect 42610 31578 42616 31580
rect 42672 31578 42696 31580
rect 42752 31578 42776 31580
rect 42832 31578 42856 31580
rect 42912 31578 42918 31580
rect 42672 31526 42674 31578
rect 42854 31526 42856 31578
rect 42610 31524 42616 31526
rect 42672 31524 42696 31526
rect 42752 31524 42776 31526
rect 42832 31524 42856 31526
rect 42912 31524 42918 31526
rect 42610 31515 42918 31524
rect 47610 31580 47918 31589
rect 47610 31578 47616 31580
rect 47672 31578 47696 31580
rect 47752 31578 47776 31580
rect 47832 31578 47856 31580
rect 47912 31578 47918 31580
rect 47672 31526 47674 31578
rect 47854 31526 47856 31578
rect 47610 31524 47616 31526
rect 47672 31524 47696 31526
rect 47752 31524 47776 31526
rect 47832 31524 47856 31526
rect 47912 31524 47918 31526
rect 47610 31515 47918 31524
rect 52610 31580 52918 31589
rect 52610 31578 52616 31580
rect 52672 31578 52696 31580
rect 52752 31578 52776 31580
rect 52832 31578 52856 31580
rect 52912 31578 52918 31580
rect 52672 31526 52674 31578
rect 52854 31526 52856 31578
rect 52610 31524 52616 31526
rect 52672 31524 52696 31526
rect 52752 31524 52776 31526
rect 52832 31524 52856 31526
rect 52912 31524 52918 31526
rect 52610 31515 52918 31524
rect 57610 31580 57918 31589
rect 57610 31578 57616 31580
rect 57672 31578 57696 31580
rect 57752 31578 57776 31580
rect 57832 31578 57856 31580
rect 57912 31578 57918 31580
rect 57672 31526 57674 31578
rect 57854 31526 57856 31578
rect 57610 31524 57616 31526
rect 57672 31524 57696 31526
rect 57752 31524 57776 31526
rect 57832 31524 57856 31526
rect 57912 31524 57918 31526
rect 57610 31515 57918 31524
rect 58532 31136 58584 31142
rect 58530 31104 58532 31113
rect 58584 31104 58586 31113
rect 1950 31036 2258 31045
rect 1950 31034 1956 31036
rect 2012 31034 2036 31036
rect 2092 31034 2116 31036
rect 2172 31034 2196 31036
rect 2252 31034 2258 31036
rect 2012 30982 2014 31034
rect 2194 30982 2196 31034
rect 1950 30980 1956 30982
rect 2012 30980 2036 30982
rect 2092 30980 2116 30982
rect 2172 30980 2196 30982
rect 2252 30980 2258 30982
rect 1950 30971 2258 30980
rect 6950 31036 7258 31045
rect 6950 31034 6956 31036
rect 7012 31034 7036 31036
rect 7092 31034 7116 31036
rect 7172 31034 7196 31036
rect 7252 31034 7258 31036
rect 7012 30982 7014 31034
rect 7194 30982 7196 31034
rect 6950 30980 6956 30982
rect 7012 30980 7036 30982
rect 7092 30980 7116 30982
rect 7172 30980 7196 30982
rect 7252 30980 7258 30982
rect 6950 30971 7258 30980
rect 11950 31036 12258 31045
rect 11950 31034 11956 31036
rect 12012 31034 12036 31036
rect 12092 31034 12116 31036
rect 12172 31034 12196 31036
rect 12252 31034 12258 31036
rect 12012 30982 12014 31034
rect 12194 30982 12196 31034
rect 11950 30980 11956 30982
rect 12012 30980 12036 30982
rect 12092 30980 12116 30982
rect 12172 30980 12196 30982
rect 12252 30980 12258 30982
rect 11950 30971 12258 30980
rect 16950 31036 17258 31045
rect 16950 31034 16956 31036
rect 17012 31034 17036 31036
rect 17092 31034 17116 31036
rect 17172 31034 17196 31036
rect 17252 31034 17258 31036
rect 17012 30982 17014 31034
rect 17194 30982 17196 31034
rect 16950 30980 16956 30982
rect 17012 30980 17036 30982
rect 17092 30980 17116 30982
rect 17172 30980 17196 30982
rect 17252 30980 17258 30982
rect 16950 30971 17258 30980
rect 21950 31036 22258 31045
rect 21950 31034 21956 31036
rect 22012 31034 22036 31036
rect 22092 31034 22116 31036
rect 22172 31034 22196 31036
rect 22252 31034 22258 31036
rect 22012 30982 22014 31034
rect 22194 30982 22196 31034
rect 21950 30980 21956 30982
rect 22012 30980 22036 30982
rect 22092 30980 22116 30982
rect 22172 30980 22196 30982
rect 22252 30980 22258 30982
rect 21950 30971 22258 30980
rect 26950 31036 27258 31045
rect 26950 31034 26956 31036
rect 27012 31034 27036 31036
rect 27092 31034 27116 31036
rect 27172 31034 27196 31036
rect 27252 31034 27258 31036
rect 27012 30982 27014 31034
rect 27194 30982 27196 31034
rect 26950 30980 26956 30982
rect 27012 30980 27036 30982
rect 27092 30980 27116 30982
rect 27172 30980 27196 30982
rect 27252 30980 27258 30982
rect 26950 30971 27258 30980
rect 31950 31036 32258 31045
rect 31950 31034 31956 31036
rect 32012 31034 32036 31036
rect 32092 31034 32116 31036
rect 32172 31034 32196 31036
rect 32252 31034 32258 31036
rect 32012 30982 32014 31034
rect 32194 30982 32196 31034
rect 31950 30980 31956 30982
rect 32012 30980 32036 30982
rect 32092 30980 32116 30982
rect 32172 30980 32196 30982
rect 32252 30980 32258 30982
rect 31950 30971 32258 30980
rect 36950 31036 37258 31045
rect 36950 31034 36956 31036
rect 37012 31034 37036 31036
rect 37092 31034 37116 31036
rect 37172 31034 37196 31036
rect 37252 31034 37258 31036
rect 37012 30982 37014 31034
rect 37194 30982 37196 31034
rect 36950 30980 36956 30982
rect 37012 30980 37036 30982
rect 37092 30980 37116 30982
rect 37172 30980 37196 30982
rect 37252 30980 37258 30982
rect 36950 30971 37258 30980
rect 41950 31036 42258 31045
rect 41950 31034 41956 31036
rect 42012 31034 42036 31036
rect 42092 31034 42116 31036
rect 42172 31034 42196 31036
rect 42252 31034 42258 31036
rect 42012 30982 42014 31034
rect 42194 30982 42196 31034
rect 41950 30980 41956 30982
rect 42012 30980 42036 30982
rect 42092 30980 42116 30982
rect 42172 30980 42196 30982
rect 42252 30980 42258 30982
rect 41950 30971 42258 30980
rect 46950 31036 47258 31045
rect 46950 31034 46956 31036
rect 47012 31034 47036 31036
rect 47092 31034 47116 31036
rect 47172 31034 47196 31036
rect 47252 31034 47258 31036
rect 47012 30982 47014 31034
rect 47194 30982 47196 31034
rect 46950 30980 46956 30982
rect 47012 30980 47036 30982
rect 47092 30980 47116 30982
rect 47172 30980 47196 30982
rect 47252 30980 47258 30982
rect 46950 30971 47258 30980
rect 51950 31036 52258 31045
rect 51950 31034 51956 31036
rect 52012 31034 52036 31036
rect 52092 31034 52116 31036
rect 52172 31034 52196 31036
rect 52252 31034 52258 31036
rect 52012 30982 52014 31034
rect 52194 30982 52196 31034
rect 51950 30980 51956 30982
rect 52012 30980 52036 30982
rect 52092 30980 52116 30982
rect 52172 30980 52196 30982
rect 52252 30980 52258 30982
rect 51950 30971 52258 30980
rect 56950 31036 57258 31045
rect 58530 31039 58586 31048
rect 56950 31034 56956 31036
rect 57012 31034 57036 31036
rect 57092 31034 57116 31036
rect 57172 31034 57196 31036
rect 57252 31034 57258 31036
rect 57012 30982 57014 31034
rect 57194 30982 57196 31034
rect 56950 30980 56956 30982
rect 57012 30980 57036 30982
rect 57092 30980 57116 30982
rect 57172 30980 57196 30982
rect 57252 30980 57258 30982
rect 56950 30971 57258 30980
rect 58532 30728 58584 30734
rect 58532 30670 58584 30676
rect 2610 30492 2918 30501
rect 2610 30490 2616 30492
rect 2672 30490 2696 30492
rect 2752 30490 2776 30492
rect 2832 30490 2856 30492
rect 2912 30490 2918 30492
rect 2672 30438 2674 30490
rect 2854 30438 2856 30490
rect 2610 30436 2616 30438
rect 2672 30436 2696 30438
rect 2752 30436 2776 30438
rect 2832 30436 2856 30438
rect 2912 30436 2918 30438
rect 2610 30427 2918 30436
rect 7610 30492 7918 30501
rect 7610 30490 7616 30492
rect 7672 30490 7696 30492
rect 7752 30490 7776 30492
rect 7832 30490 7856 30492
rect 7912 30490 7918 30492
rect 7672 30438 7674 30490
rect 7854 30438 7856 30490
rect 7610 30436 7616 30438
rect 7672 30436 7696 30438
rect 7752 30436 7776 30438
rect 7832 30436 7856 30438
rect 7912 30436 7918 30438
rect 7610 30427 7918 30436
rect 12610 30492 12918 30501
rect 12610 30490 12616 30492
rect 12672 30490 12696 30492
rect 12752 30490 12776 30492
rect 12832 30490 12856 30492
rect 12912 30490 12918 30492
rect 12672 30438 12674 30490
rect 12854 30438 12856 30490
rect 12610 30436 12616 30438
rect 12672 30436 12696 30438
rect 12752 30436 12776 30438
rect 12832 30436 12856 30438
rect 12912 30436 12918 30438
rect 12610 30427 12918 30436
rect 17610 30492 17918 30501
rect 17610 30490 17616 30492
rect 17672 30490 17696 30492
rect 17752 30490 17776 30492
rect 17832 30490 17856 30492
rect 17912 30490 17918 30492
rect 17672 30438 17674 30490
rect 17854 30438 17856 30490
rect 17610 30436 17616 30438
rect 17672 30436 17696 30438
rect 17752 30436 17776 30438
rect 17832 30436 17856 30438
rect 17912 30436 17918 30438
rect 17610 30427 17918 30436
rect 22610 30492 22918 30501
rect 22610 30490 22616 30492
rect 22672 30490 22696 30492
rect 22752 30490 22776 30492
rect 22832 30490 22856 30492
rect 22912 30490 22918 30492
rect 22672 30438 22674 30490
rect 22854 30438 22856 30490
rect 22610 30436 22616 30438
rect 22672 30436 22696 30438
rect 22752 30436 22776 30438
rect 22832 30436 22856 30438
rect 22912 30436 22918 30438
rect 22610 30427 22918 30436
rect 27610 30492 27918 30501
rect 27610 30490 27616 30492
rect 27672 30490 27696 30492
rect 27752 30490 27776 30492
rect 27832 30490 27856 30492
rect 27912 30490 27918 30492
rect 27672 30438 27674 30490
rect 27854 30438 27856 30490
rect 27610 30436 27616 30438
rect 27672 30436 27696 30438
rect 27752 30436 27776 30438
rect 27832 30436 27856 30438
rect 27912 30436 27918 30438
rect 27610 30427 27918 30436
rect 32610 30492 32918 30501
rect 32610 30490 32616 30492
rect 32672 30490 32696 30492
rect 32752 30490 32776 30492
rect 32832 30490 32856 30492
rect 32912 30490 32918 30492
rect 32672 30438 32674 30490
rect 32854 30438 32856 30490
rect 32610 30436 32616 30438
rect 32672 30436 32696 30438
rect 32752 30436 32776 30438
rect 32832 30436 32856 30438
rect 32912 30436 32918 30438
rect 32610 30427 32918 30436
rect 37610 30492 37918 30501
rect 37610 30490 37616 30492
rect 37672 30490 37696 30492
rect 37752 30490 37776 30492
rect 37832 30490 37856 30492
rect 37912 30490 37918 30492
rect 37672 30438 37674 30490
rect 37854 30438 37856 30490
rect 37610 30436 37616 30438
rect 37672 30436 37696 30438
rect 37752 30436 37776 30438
rect 37832 30436 37856 30438
rect 37912 30436 37918 30438
rect 37610 30427 37918 30436
rect 42610 30492 42918 30501
rect 42610 30490 42616 30492
rect 42672 30490 42696 30492
rect 42752 30490 42776 30492
rect 42832 30490 42856 30492
rect 42912 30490 42918 30492
rect 42672 30438 42674 30490
rect 42854 30438 42856 30490
rect 42610 30436 42616 30438
rect 42672 30436 42696 30438
rect 42752 30436 42776 30438
rect 42832 30436 42856 30438
rect 42912 30436 42918 30438
rect 42610 30427 42918 30436
rect 47610 30492 47918 30501
rect 47610 30490 47616 30492
rect 47672 30490 47696 30492
rect 47752 30490 47776 30492
rect 47832 30490 47856 30492
rect 47912 30490 47918 30492
rect 47672 30438 47674 30490
rect 47854 30438 47856 30490
rect 47610 30436 47616 30438
rect 47672 30436 47696 30438
rect 47752 30436 47776 30438
rect 47832 30436 47856 30438
rect 47912 30436 47918 30438
rect 47610 30427 47918 30436
rect 52610 30492 52918 30501
rect 52610 30490 52616 30492
rect 52672 30490 52696 30492
rect 52752 30490 52776 30492
rect 52832 30490 52856 30492
rect 52912 30490 52918 30492
rect 52672 30438 52674 30490
rect 52854 30438 52856 30490
rect 52610 30436 52616 30438
rect 52672 30436 52696 30438
rect 52752 30436 52776 30438
rect 52832 30436 52856 30438
rect 52912 30436 52918 30438
rect 52610 30427 52918 30436
rect 57610 30492 57918 30501
rect 57610 30490 57616 30492
rect 57672 30490 57696 30492
rect 57752 30490 57776 30492
rect 57832 30490 57856 30492
rect 57912 30490 57918 30492
rect 57672 30438 57674 30490
rect 57854 30438 57856 30490
rect 57610 30436 57616 30438
rect 57672 30436 57696 30438
rect 57752 30436 57776 30438
rect 57832 30436 57856 30438
rect 57912 30436 57918 30438
rect 57610 30427 57918 30436
rect 58544 30297 58572 30670
rect 58530 30288 58586 30297
rect 58530 30223 58586 30232
rect 1950 29948 2258 29957
rect 1950 29946 1956 29948
rect 2012 29946 2036 29948
rect 2092 29946 2116 29948
rect 2172 29946 2196 29948
rect 2252 29946 2258 29948
rect 2012 29894 2014 29946
rect 2194 29894 2196 29946
rect 1950 29892 1956 29894
rect 2012 29892 2036 29894
rect 2092 29892 2116 29894
rect 2172 29892 2196 29894
rect 2252 29892 2258 29894
rect 1950 29883 2258 29892
rect 6950 29948 7258 29957
rect 6950 29946 6956 29948
rect 7012 29946 7036 29948
rect 7092 29946 7116 29948
rect 7172 29946 7196 29948
rect 7252 29946 7258 29948
rect 7012 29894 7014 29946
rect 7194 29894 7196 29946
rect 6950 29892 6956 29894
rect 7012 29892 7036 29894
rect 7092 29892 7116 29894
rect 7172 29892 7196 29894
rect 7252 29892 7258 29894
rect 6950 29883 7258 29892
rect 11950 29948 12258 29957
rect 11950 29946 11956 29948
rect 12012 29946 12036 29948
rect 12092 29946 12116 29948
rect 12172 29946 12196 29948
rect 12252 29946 12258 29948
rect 12012 29894 12014 29946
rect 12194 29894 12196 29946
rect 11950 29892 11956 29894
rect 12012 29892 12036 29894
rect 12092 29892 12116 29894
rect 12172 29892 12196 29894
rect 12252 29892 12258 29894
rect 11950 29883 12258 29892
rect 16950 29948 17258 29957
rect 16950 29946 16956 29948
rect 17012 29946 17036 29948
rect 17092 29946 17116 29948
rect 17172 29946 17196 29948
rect 17252 29946 17258 29948
rect 17012 29894 17014 29946
rect 17194 29894 17196 29946
rect 16950 29892 16956 29894
rect 17012 29892 17036 29894
rect 17092 29892 17116 29894
rect 17172 29892 17196 29894
rect 17252 29892 17258 29894
rect 16950 29883 17258 29892
rect 21950 29948 22258 29957
rect 21950 29946 21956 29948
rect 22012 29946 22036 29948
rect 22092 29946 22116 29948
rect 22172 29946 22196 29948
rect 22252 29946 22258 29948
rect 22012 29894 22014 29946
rect 22194 29894 22196 29946
rect 21950 29892 21956 29894
rect 22012 29892 22036 29894
rect 22092 29892 22116 29894
rect 22172 29892 22196 29894
rect 22252 29892 22258 29894
rect 21950 29883 22258 29892
rect 26950 29948 27258 29957
rect 26950 29946 26956 29948
rect 27012 29946 27036 29948
rect 27092 29946 27116 29948
rect 27172 29946 27196 29948
rect 27252 29946 27258 29948
rect 27012 29894 27014 29946
rect 27194 29894 27196 29946
rect 26950 29892 26956 29894
rect 27012 29892 27036 29894
rect 27092 29892 27116 29894
rect 27172 29892 27196 29894
rect 27252 29892 27258 29894
rect 26950 29883 27258 29892
rect 31950 29948 32258 29957
rect 31950 29946 31956 29948
rect 32012 29946 32036 29948
rect 32092 29946 32116 29948
rect 32172 29946 32196 29948
rect 32252 29946 32258 29948
rect 32012 29894 32014 29946
rect 32194 29894 32196 29946
rect 31950 29892 31956 29894
rect 32012 29892 32036 29894
rect 32092 29892 32116 29894
rect 32172 29892 32196 29894
rect 32252 29892 32258 29894
rect 31950 29883 32258 29892
rect 36950 29948 37258 29957
rect 36950 29946 36956 29948
rect 37012 29946 37036 29948
rect 37092 29946 37116 29948
rect 37172 29946 37196 29948
rect 37252 29946 37258 29948
rect 37012 29894 37014 29946
rect 37194 29894 37196 29946
rect 36950 29892 36956 29894
rect 37012 29892 37036 29894
rect 37092 29892 37116 29894
rect 37172 29892 37196 29894
rect 37252 29892 37258 29894
rect 36950 29883 37258 29892
rect 41950 29948 42258 29957
rect 41950 29946 41956 29948
rect 42012 29946 42036 29948
rect 42092 29946 42116 29948
rect 42172 29946 42196 29948
rect 42252 29946 42258 29948
rect 42012 29894 42014 29946
rect 42194 29894 42196 29946
rect 41950 29892 41956 29894
rect 42012 29892 42036 29894
rect 42092 29892 42116 29894
rect 42172 29892 42196 29894
rect 42252 29892 42258 29894
rect 41950 29883 42258 29892
rect 46950 29948 47258 29957
rect 46950 29946 46956 29948
rect 47012 29946 47036 29948
rect 47092 29946 47116 29948
rect 47172 29946 47196 29948
rect 47252 29946 47258 29948
rect 47012 29894 47014 29946
rect 47194 29894 47196 29946
rect 46950 29892 46956 29894
rect 47012 29892 47036 29894
rect 47092 29892 47116 29894
rect 47172 29892 47196 29894
rect 47252 29892 47258 29894
rect 46950 29883 47258 29892
rect 51950 29948 52258 29957
rect 51950 29946 51956 29948
rect 52012 29946 52036 29948
rect 52092 29946 52116 29948
rect 52172 29946 52196 29948
rect 52252 29946 52258 29948
rect 52012 29894 52014 29946
rect 52194 29894 52196 29946
rect 51950 29892 51956 29894
rect 52012 29892 52036 29894
rect 52092 29892 52116 29894
rect 52172 29892 52196 29894
rect 52252 29892 52258 29894
rect 51950 29883 52258 29892
rect 56950 29948 57258 29957
rect 56950 29946 56956 29948
rect 57012 29946 57036 29948
rect 57092 29946 57116 29948
rect 57172 29946 57196 29948
rect 57252 29946 57258 29948
rect 57012 29894 57014 29946
rect 57194 29894 57196 29946
rect 56950 29892 56956 29894
rect 57012 29892 57036 29894
rect 57092 29892 57116 29894
rect 57172 29892 57196 29894
rect 57252 29892 57258 29894
rect 56950 29883 57258 29892
rect 58532 29640 58584 29646
rect 58532 29582 58584 29588
rect 58544 29481 58572 29582
rect 58530 29472 58586 29481
rect 2610 29404 2918 29413
rect 2610 29402 2616 29404
rect 2672 29402 2696 29404
rect 2752 29402 2776 29404
rect 2832 29402 2856 29404
rect 2912 29402 2918 29404
rect 2672 29350 2674 29402
rect 2854 29350 2856 29402
rect 2610 29348 2616 29350
rect 2672 29348 2696 29350
rect 2752 29348 2776 29350
rect 2832 29348 2856 29350
rect 2912 29348 2918 29350
rect 2610 29339 2918 29348
rect 7610 29404 7918 29413
rect 7610 29402 7616 29404
rect 7672 29402 7696 29404
rect 7752 29402 7776 29404
rect 7832 29402 7856 29404
rect 7912 29402 7918 29404
rect 7672 29350 7674 29402
rect 7854 29350 7856 29402
rect 7610 29348 7616 29350
rect 7672 29348 7696 29350
rect 7752 29348 7776 29350
rect 7832 29348 7856 29350
rect 7912 29348 7918 29350
rect 7610 29339 7918 29348
rect 12610 29404 12918 29413
rect 12610 29402 12616 29404
rect 12672 29402 12696 29404
rect 12752 29402 12776 29404
rect 12832 29402 12856 29404
rect 12912 29402 12918 29404
rect 12672 29350 12674 29402
rect 12854 29350 12856 29402
rect 12610 29348 12616 29350
rect 12672 29348 12696 29350
rect 12752 29348 12776 29350
rect 12832 29348 12856 29350
rect 12912 29348 12918 29350
rect 12610 29339 12918 29348
rect 17610 29404 17918 29413
rect 17610 29402 17616 29404
rect 17672 29402 17696 29404
rect 17752 29402 17776 29404
rect 17832 29402 17856 29404
rect 17912 29402 17918 29404
rect 17672 29350 17674 29402
rect 17854 29350 17856 29402
rect 17610 29348 17616 29350
rect 17672 29348 17696 29350
rect 17752 29348 17776 29350
rect 17832 29348 17856 29350
rect 17912 29348 17918 29350
rect 17610 29339 17918 29348
rect 22610 29404 22918 29413
rect 22610 29402 22616 29404
rect 22672 29402 22696 29404
rect 22752 29402 22776 29404
rect 22832 29402 22856 29404
rect 22912 29402 22918 29404
rect 22672 29350 22674 29402
rect 22854 29350 22856 29402
rect 22610 29348 22616 29350
rect 22672 29348 22696 29350
rect 22752 29348 22776 29350
rect 22832 29348 22856 29350
rect 22912 29348 22918 29350
rect 22610 29339 22918 29348
rect 27610 29404 27918 29413
rect 27610 29402 27616 29404
rect 27672 29402 27696 29404
rect 27752 29402 27776 29404
rect 27832 29402 27856 29404
rect 27912 29402 27918 29404
rect 27672 29350 27674 29402
rect 27854 29350 27856 29402
rect 27610 29348 27616 29350
rect 27672 29348 27696 29350
rect 27752 29348 27776 29350
rect 27832 29348 27856 29350
rect 27912 29348 27918 29350
rect 27610 29339 27918 29348
rect 32610 29404 32918 29413
rect 32610 29402 32616 29404
rect 32672 29402 32696 29404
rect 32752 29402 32776 29404
rect 32832 29402 32856 29404
rect 32912 29402 32918 29404
rect 32672 29350 32674 29402
rect 32854 29350 32856 29402
rect 32610 29348 32616 29350
rect 32672 29348 32696 29350
rect 32752 29348 32776 29350
rect 32832 29348 32856 29350
rect 32912 29348 32918 29350
rect 32610 29339 32918 29348
rect 37610 29404 37918 29413
rect 37610 29402 37616 29404
rect 37672 29402 37696 29404
rect 37752 29402 37776 29404
rect 37832 29402 37856 29404
rect 37912 29402 37918 29404
rect 37672 29350 37674 29402
rect 37854 29350 37856 29402
rect 37610 29348 37616 29350
rect 37672 29348 37696 29350
rect 37752 29348 37776 29350
rect 37832 29348 37856 29350
rect 37912 29348 37918 29350
rect 37610 29339 37918 29348
rect 42610 29404 42918 29413
rect 42610 29402 42616 29404
rect 42672 29402 42696 29404
rect 42752 29402 42776 29404
rect 42832 29402 42856 29404
rect 42912 29402 42918 29404
rect 42672 29350 42674 29402
rect 42854 29350 42856 29402
rect 42610 29348 42616 29350
rect 42672 29348 42696 29350
rect 42752 29348 42776 29350
rect 42832 29348 42856 29350
rect 42912 29348 42918 29350
rect 42610 29339 42918 29348
rect 47610 29404 47918 29413
rect 47610 29402 47616 29404
rect 47672 29402 47696 29404
rect 47752 29402 47776 29404
rect 47832 29402 47856 29404
rect 47912 29402 47918 29404
rect 47672 29350 47674 29402
rect 47854 29350 47856 29402
rect 47610 29348 47616 29350
rect 47672 29348 47696 29350
rect 47752 29348 47776 29350
rect 47832 29348 47856 29350
rect 47912 29348 47918 29350
rect 47610 29339 47918 29348
rect 52610 29404 52918 29413
rect 52610 29402 52616 29404
rect 52672 29402 52696 29404
rect 52752 29402 52776 29404
rect 52832 29402 52856 29404
rect 52912 29402 52918 29404
rect 52672 29350 52674 29402
rect 52854 29350 52856 29402
rect 52610 29348 52616 29350
rect 52672 29348 52696 29350
rect 52752 29348 52776 29350
rect 52832 29348 52856 29350
rect 52912 29348 52918 29350
rect 52610 29339 52918 29348
rect 57610 29404 57918 29413
rect 58530 29407 58586 29416
rect 57610 29402 57616 29404
rect 57672 29402 57696 29404
rect 57752 29402 57776 29404
rect 57832 29402 57856 29404
rect 57912 29402 57918 29404
rect 57672 29350 57674 29402
rect 57854 29350 57856 29402
rect 57610 29348 57616 29350
rect 57672 29348 57696 29350
rect 57752 29348 57776 29350
rect 57832 29348 57856 29350
rect 57912 29348 57918 29350
rect 57610 29339 57918 29348
rect 58532 29028 58584 29034
rect 58532 28970 58584 28976
rect 1950 28860 2258 28869
rect 1950 28858 1956 28860
rect 2012 28858 2036 28860
rect 2092 28858 2116 28860
rect 2172 28858 2196 28860
rect 2252 28858 2258 28860
rect 2012 28806 2014 28858
rect 2194 28806 2196 28858
rect 1950 28804 1956 28806
rect 2012 28804 2036 28806
rect 2092 28804 2116 28806
rect 2172 28804 2196 28806
rect 2252 28804 2258 28806
rect 1950 28795 2258 28804
rect 6950 28860 7258 28869
rect 6950 28858 6956 28860
rect 7012 28858 7036 28860
rect 7092 28858 7116 28860
rect 7172 28858 7196 28860
rect 7252 28858 7258 28860
rect 7012 28806 7014 28858
rect 7194 28806 7196 28858
rect 6950 28804 6956 28806
rect 7012 28804 7036 28806
rect 7092 28804 7116 28806
rect 7172 28804 7196 28806
rect 7252 28804 7258 28806
rect 6950 28795 7258 28804
rect 11950 28860 12258 28869
rect 11950 28858 11956 28860
rect 12012 28858 12036 28860
rect 12092 28858 12116 28860
rect 12172 28858 12196 28860
rect 12252 28858 12258 28860
rect 12012 28806 12014 28858
rect 12194 28806 12196 28858
rect 11950 28804 11956 28806
rect 12012 28804 12036 28806
rect 12092 28804 12116 28806
rect 12172 28804 12196 28806
rect 12252 28804 12258 28806
rect 11950 28795 12258 28804
rect 16950 28860 17258 28869
rect 16950 28858 16956 28860
rect 17012 28858 17036 28860
rect 17092 28858 17116 28860
rect 17172 28858 17196 28860
rect 17252 28858 17258 28860
rect 17012 28806 17014 28858
rect 17194 28806 17196 28858
rect 16950 28804 16956 28806
rect 17012 28804 17036 28806
rect 17092 28804 17116 28806
rect 17172 28804 17196 28806
rect 17252 28804 17258 28806
rect 16950 28795 17258 28804
rect 21950 28860 22258 28869
rect 21950 28858 21956 28860
rect 22012 28858 22036 28860
rect 22092 28858 22116 28860
rect 22172 28858 22196 28860
rect 22252 28858 22258 28860
rect 22012 28806 22014 28858
rect 22194 28806 22196 28858
rect 21950 28804 21956 28806
rect 22012 28804 22036 28806
rect 22092 28804 22116 28806
rect 22172 28804 22196 28806
rect 22252 28804 22258 28806
rect 21950 28795 22258 28804
rect 26950 28860 27258 28869
rect 26950 28858 26956 28860
rect 27012 28858 27036 28860
rect 27092 28858 27116 28860
rect 27172 28858 27196 28860
rect 27252 28858 27258 28860
rect 27012 28806 27014 28858
rect 27194 28806 27196 28858
rect 26950 28804 26956 28806
rect 27012 28804 27036 28806
rect 27092 28804 27116 28806
rect 27172 28804 27196 28806
rect 27252 28804 27258 28806
rect 26950 28795 27258 28804
rect 31950 28860 32258 28869
rect 31950 28858 31956 28860
rect 32012 28858 32036 28860
rect 32092 28858 32116 28860
rect 32172 28858 32196 28860
rect 32252 28858 32258 28860
rect 32012 28806 32014 28858
rect 32194 28806 32196 28858
rect 31950 28804 31956 28806
rect 32012 28804 32036 28806
rect 32092 28804 32116 28806
rect 32172 28804 32196 28806
rect 32252 28804 32258 28806
rect 31950 28795 32258 28804
rect 36950 28860 37258 28869
rect 36950 28858 36956 28860
rect 37012 28858 37036 28860
rect 37092 28858 37116 28860
rect 37172 28858 37196 28860
rect 37252 28858 37258 28860
rect 37012 28806 37014 28858
rect 37194 28806 37196 28858
rect 36950 28804 36956 28806
rect 37012 28804 37036 28806
rect 37092 28804 37116 28806
rect 37172 28804 37196 28806
rect 37252 28804 37258 28806
rect 36950 28795 37258 28804
rect 41950 28860 42258 28869
rect 41950 28858 41956 28860
rect 42012 28858 42036 28860
rect 42092 28858 42116 28860
rect 42172 28858 42196 28860
rect 42252 28858 42258 28860
rect 42012 28806 42014 28858
rect 42194 28806 42196 28858
rect 41950 28804 41956 28806
rect 42012 28804 42036 28806
rect 42092 28804 42116 28806
rect 42172 28804 42196 28806
rect 42252 28804 42258 28806
rect 41950 28795 42258 28804
rect 46950 28860 47258 28869
rect 46950 28858 46956 28860
rect 47012 28858 47036 28860
rect 47092 28858 47116 28860
rect 47172 28858 47196 28860
rect 47252 28858 47258 28860
rect 47012 28806 47014 28858
rect 47194 28806 47196 28858
rect 46950 28804 46956 28806
rect 47012 28804 47036 28806
rect 47092 28804 47116 28806
rect 47172 28804 47196 28806
rect 47252 28804 47258 28806
rect 46950 28795 47258 28804
rect 51950 28860 52258 28869
rect 51950 28858 51956 28860
rect 52012 28858 52036 28860
rect 52092 28858 52116 28860
rect 52172 28858 52196 28860
rect 52252 28858 52258 28860
rect 52012 28806 52014 28858
rect 52194 28806 52196 28858
rect 51950 28804 51956 28806
rect 52012 28804 52036 28806
rect 52092 28804 52116 28806
rect 52172 28804 52196 28806
rect 52252 28804 52258 28806
rect 51950 28795 52258 28804
rect 56950 28860 57258 28869
rect 56950 28858 56956 28860
rect 57012 28858 57036 28860
rect 57092 28858 57116 28860
rect 57172 28858 57196 28860
rect 57252 28858 57258 28860
rect 57012 28806 57014 28858
rect 57194 28806 57196 28858
rect 56950 28804 56956 28806
rect 57012 28804 57036 28806
rect 57092 28804 57116 28806
rect 57172 28804 57196 28806
rect 57252 28804 57258 28806
rect 56950 28795 57258 28804
rect 58544 28665 58572 28970
rect 58530 28656 58586 28665
rect 58530 28591 58586 28600
rect 2610 28316 2918 28325
rect 2610 28314 2616 28316
rect 2672 28314 2696 28316
rect 2752 28314 2776 28316
rect 2832 28314 2856 28316
rect 2912 28314 2918 28316
rect 2672 28262 2674 28314
rect 2854 28262 2856 28314
rect 2610 28260 2616 28262
rect 2672 28260 2696 28262
rect 2752 28260 2776 28262
rect 2832 28260 2856 28262
rect 2912 28260 2918 28262
rect 2610 28251 2918 28260
rect 7610 28316 7918 28325
rect 7610 28314 7616 28316
rect 7672 28314 7696 28316
rect 7752 28314 7776 28316
rect 7832 28314 7856 28316
rect 7912 28314 7918 28316
rect 7672 28262 7674 28314
rect 7854 28262 7856 28314
rect 7610 28260 7616 28262
rect 7672 28260 7696 28262
rect 7752 28260 7776 28262
rect 7832 28260 7856 28262
rect 7912 28260 7918 28262
rect 7610 28251 7918 28260
rect 12610 28316 12918 28325
rect 12610 28314 12616 28316
rect 12672 28314 12696 28316
rect 12752 28314 12776 28316
rect 12832 28314 12856 28316
rect 12912 28314 12918 28316
rect 12672 28262 12674 28314
rect 12854 28262 12856 28314
rect 12610 28260 12616 28262
rect 12672 28260 12696 28262
rect 12752 28260 12776 28262
rect 12832 28260 12856 28262
rect 12912 28260 12918 28262
rect 12610 28251 12918 28260
rect 17610 28316 17918 28325
rect 17610 28314 17616 28316
rect 17672 28314 17696 28316
rect 17752 28314 17776 28316
rect 17832 28314 17856 28316
rect 17912 28314 17918 28316
rect 17672 28262 17674 28314
rect 17854 28262 17856 28314
rect 17610 28260 17616 28262
rect 17672 28260 17696 28262
rect 17752 28260 17776 28262
rect 17832 28260 17856 28262
rect 17912 28260 17918 28262
rect 17610 28251 17918 28260
rect 22610 28316 22918 28325
rect 22610 28314 22616 28316
rect 22672 28314 22696 28316
rect 22752 28314 22776 28316
rect 22832 28314 22856 28316
rect 22912 28314 22918 28316
rect 22672 28262 22674 28314
rect 22854 28262 22856 28314
rect 22610 28260 22616 28262
rect 22672 28260 22696 28262
rect 22752 28260 22776 28262
rect 22832 28260 22856 28262
rect 22912 28260 22918 28262
rect 22610 28251 22918 28260
rect 27610 28316 27918 28325
rect 27610 28314 27616 28316
rect 27672 28314 27696 28316
rect 27752 28314 27776 28316
rect 27832 28314 27856 28316
rect 27912 28314 27918 28316
rect 27672 28262 27674 28314
rect 27854 28262 27856 28314
rect 27610 28260 27616 28262
rect 27672 28260 27696 28262
rect 27752 28260 27776 28262
rect 27832 28260 27856 28262
rect 27912 28260 27918 28262
rect 27610 28251 27918 28260
rect 32610 28316 32918 28325
rect 32610 28314 32616 28316
rect 32672 28314 32696 28316
rect 32752 28314 32776 28316
rect 32832 28314 32856 28316
rect 32912 28314 32918 28316
rect 32672 28262 32674 28314
rect 32854 28262 32856 28314
rect 32610 28260 32616 28262
rect 32672 28260 32696 28262
rect 32752 28260 32776 28262
rect 32832 28260 32856 28262
rect 32912 28260 32918 28262
rect 32610 28251 32918 28260
rect 37610 28316 37918 28325
rect 37610 28314 37616 28316
rect 37672 28314 37696 28316
rect 37752 28314 37776 28316
rect 37832 28314 37856 28316
rect 37912 28314 37918 28316
rect 37672 28262 37674 28314
rect 37854 28262 37856 28314
rect 37610 28260 37616 28262
rect 37672 28260 37696 28262
rect 37752 28260 37776 28262
rect 37832 28260 37856 28262
rect 37912 28260 37918 28262
rect 37610 28251 37918 28260
rect 42610 28316 42918 28325
rect 42610 28314 42616 28316
rect 42672 28314 42696 28316
rect 42752 28314 42776 28316
rect 42832 28314 42856 28316
rect 42912 28314 42918 28316
rect 42672 28262 42674 28314
rect 42854 28262 42856 28314
rect 42610 28260 42616 28262
rect 42672 28260 42696 28262
rect 42752 28260 42776 28262
rect 42832 28260 42856 28262
rect 42912 28260 42918 28262
rect 42610 28251 42918 28260
rect 47610 28316 47918 28325
rect 47610 28314 47616 28316
rect 47672 28314 47696 28316
rect 47752 28314 47776 28316
rect 47832 28314 47856 28316
rect 47912 28314 47918 28316
rect 47672 28262 47674 28314
rect 47854 28262 47856 28314
rect 47610 28260 47616 28262
rect 47672 28260 47696 28262
rect 47752 28260 47776 28262
rect 47832 28260 47856 28262
rect 47912 28260 47918 28262
rect 47610 28251 47918 28260
rect 52610 28316 52918 28325
rect 52610 28314 52616 28316
rect 52672 28314 52696 28316
rect 52752 28314 52776 28316
rect 52832 28314 52856 28316
rect 52912 28314 52918 28316
rect 52672 28262 52674 28314
rect 52854 28262 52856 28314
rect 52610 28260 52616 28262
rect 52672 28260 52696 28262
rect 52752 28260 52776 28262
rect 52832 28260 52856 28262
rect 52912 28260 52918 28262
rect 52610 28251 52918 28260
rect 57610 28316 57918 28325
rect 57610 28314 57616 28316
rect 57672 28314 57696 28316
rect 57752 28314 57776 28316
rect 57832 28314 57856 28316
rect 57912 28314 57918 28316
rect 57672 28262 57674 28314
rect 57854 28262 57856 28314
rect 57610 28260 57616 28262
rect 57672 28260 57696 28262
rect 57752 28260 57776 28262
rect 57832 28260 57856 28262
rect 57912 28260 57918 28262
rect 57610 28251 57918 28260
rect 58532 27872 58584 27878
rect 58530 27840 58532 27849
rect 58584 27840 58586 27849
rect 1950 27772 2258 27781
rect 1950 27770 1956 27772
rect 2012 27770 2036 27772
rect 2092 27770 2116 27772
rect 2172 27770 2196 27772
rect 2252 27770 2258 27772
rect 2012 27718 2014 27770
rect 2194 27718 2196 27770
rect 1950 27716 1956 27718
rect 2012 27716 2036 27718
rect 2092 27716 2116 27718
rect 2172 27716 2196 27718
rect 2252 27716 2258 27718
rect 1950 27707 2258 27716
rect 6950 27772 7258 27781
rect 6950 27770 6956 27772
rect 7012 27770 7036 27772
rect 7092 27770 7116 27772
rect 7172 27770 7196 27772
rect 7252 27770 7258 27772
rect 7012 27718 7014 27770
rect 7194 27718 7196 27770
rect 6950 27716 6956 27718
rect 7012 27716 7036 27718
rect 7092 27716 7116 27718
rect 7172 27716 7196 27718
rect 7252 27716 7258 27718
rect 6950 27707 7258 27716
rect 11950 27772 12258 27781
rect 11950 27770 11956 27772
rect 12012 27770 12036 27772
rect 12092 27770 12116 27772
rect 12172 27770 12196 27772
rect 12252 27770 12258 27772
rect 12012 27718 12014 27770
rect 12194 27718 12196 27770
rect 11950 27716 11956 27718
rect 12012 27716 12036 27718
rect 12092 27716 12116 27718
rect 12172 27716 12196 27718
rect 12252 27716 12258 27718
rect 11950 27707 12258 27716
rect 16950 27772 17258 27781
rect 16950 27770 16956 27772
rect 17012 27770 17036 27772
rect 17092 27770 17116 27772
rect 17172 27770 17196 27772
rect 17252 27770 17258 27772
rect 17012 27718 17014 27770
rect 17194 27718 17196 27770
rect 16950 27716 16956 27718
rect 17012 27716 17036 27718
rect 17092 27716 17116 27718
rect 17172 27716 17196 27718
rect 17252 27716 17258 27718
rect 16950 27707 17258 27716
rect 21950 27772 22258 27781
rect 21950 27770 21956 27772
rect 22012 27770 22036 27772
rect 22092 27770 22116 27772
rect 22172 27770 22196 27772
rect 22252 27770 22258 27772
rect 22012 27718 22014 27770
rect 22194 27718 22196 27770
rect 21950 27716 21956 27718
rect 22012 27716 22036 27718
rect 22092 27716 22116 27718
rect 22172 27716 22196 27718
rect 22252 27716 22258 27718
rect 21950 27707 22258 27716
rect 26950 27772 27258 27781
rect 26950 27770 26956 27772
rect 27012 27770 27036 27772
rect 27092 27770 27116 27772
rect 27172 27770 27196 27772
rect 27252 27770 27258 27772
rect 27012 27718 27014 27770
rect 27194 27718 27196 27770
rect 26950 27716 26956 27718
rect 27012 27716 27036 27718
rect 27092 27716 27116 27718
rect 27172 27716 27196 27718
rect 27252 27716 27258 27718
rect 26950 27707 27258 27716
rect 31950 27772 32258 27781
rect 31950 27770 31956 27772
rect 32012 27770 32036 27772
rect 32092 27770 32116 27772
rect 32172 27770 32196 27772
rect 32252 27770 32258 27772
rect 32012 27718 32014 27770
rect 32194 27718 32196 27770
rect 31950 27716 31956 27718
rect 32012 27716 32036 27718
rect 32092 27716 32116 27718
rect 32172 27716 32196 27718
rect 32252 27716 32258 27718
rect 31950 27707 32258 27716
rect 36950 27772 37258 27781
rect 36950 27770 36956 27772
rect 37012 27770 37036 27772
rect 37092 27770 37116 27772
rect 37172 27770 37196 27772
rect 37252 27770 37258 27772
rect 37012 27718 37014 27770
rect 37194 27718 37196 27770
rect 36950 27716 36956 27718
rect 37012 27716 37036 27718
rect 37092 27716 37116 27718
rect 37172 27716 37196 27718
rect 37252 27716 37258 27718
rect 36950 27707 37258 27716
rect 41950 27772 42258 27781
rect 41950 27770 41956 27772
rect 42012 27770 42036 27772
rect 42092 27770 42116 27772
rect 42172 27770 42196 27772
rect 42252 27770 42258 27772
rect 42012 27718 42014 27770
rect 42194 27718 42196 27770
rect 41950 27716 41956 27718
rect 42012 27716 42036 27718
rect 42092 27716 42116 27718
rect 42172 27716 42196 27718
rect 42252 27716 42258 27718
rect 41950 27707 42258 27716
rect 46950 27772 47258 27781
rect 46950 27770 46956 27772
rect 47012 27770 47036 27772
rect 47092 27770 47116 27772
rect 47172 27770 47196 27772
rect 47252 27770 47258 27772
rect 47012 27718 47014 27770
rect 47194 27718 47196 27770
rect 46950 27716 46956 27718
rect 47012 27716 47036 27718
rect 47092 27716 47116 27718
rect 47172 27716 47196 27718
rect 47252 27716 47258 27718
rect 46950 27707 47258 27716
rect 51950 27772 52258 27781
rect 51950 27770 51956 27772
rect 52012 27770 52036 27772
rect 52092 27770 52116 27772
rect 52172 27770 52196 27772
rect 52252 27770 52258 27772
rect 52012 27718 52014 27770
rect 52194 27718 52196 27770
rect 51950 27716 51956 27718
rect 52012 27716 52036 27718
rect 52092 27716 52116 27718
rect 52172 27716 52196 27718
rect 52252 27716 52258 27718
rect 51950 27707 52258 27716
rect 56950 27772 57258 27781
rect 58530 27775 58586 27784
rect 56950 27770 56956 27772
rect 57012 27770 57036 27772
rect 57092 27770 57116 27772
rect 57172 27770 57196 27772
rect 57252 27770 57258 27772
rect 57012 27718 57014 27770
rect 57194 27718 57196 27770
rect 56950 27716 56956 27718
rect 57012 27716 57036 27718
rect 57092 27716 57116 27718
rect 57172 27716 57196 27718
rect 57252 27716 57258 27718
rect 56950 27707 57258 27716
rect 58532 27464 58584 27470
rect 58532 27406 58584 27412
rect 2610 27228 2918 27237
rect 2610 27226 2616 27228
rect 2672 27226 2696 27228
rect 2752 27226 2776 27228
rect 2832 27226 2856 27228
rect 2912 27226 2918 27228
rect 2672 27174 2674 27226
rect 2854 27174 2856 27226
rect 2610 27172 2616 27174
rect 2672 27172 2696 27174
rect 2752 27172 2776 27174
rect 2832 27172 2856 27174
rect 2912 27172 2918 27174
rect 2610 27163 2918 27172
rect 7610 27228 7918 27237
rect 7610 27226 7616 27228
rect 7672 27226 7696 27228
rect 7752 27226 7776 27228
rect 7832 27226 7856 27228
rect 7912 27226 7918 27228
rect 7672 27174 7674 27226
rect 7854 27174 7856 27226
rect 7610 27172 7616 27174
rect 7672 27172 7696 27174
rect 7752 27172 7776 27174
rect 7832 27172 7856 27174
rect 7912 27172 7918 27174
rect 7610 27163 7918 27172
rect 12610 27228 12918 27237
rect 12610 27226 12616 27228
rect 12672 27226 12696 27228
rect 12752 27226 12776 27228
rect 12832 27226 12856 27228
rect 12912 27226 12918 27228
rect 12672 27174 12674 27226
rect 12854 27174 12856 27226
rect 12610 27172 12616 27174
rect 12672 27172 12696 27174
rect 12752 27172 12776 27174
rect 12832 27172 12856 27174
rect 12912 27172 12918 27174
rect 12610 27163 12918 27172
rect 17610 27228 17918 27237
rect 17610 27226 17616 27228
rect 17672 27226 17696 27228
rect 17752 27226 17776 27228
rect 17832 27226 17856 27228
rect 17912 27226 17918 27228
rect 17672 27174 17674 27226
rect 17854 27174 17856 27226
rect 17610 27172 17616 27174
rect 17672 27172 17696 27174
rect 17752 27172 17776 27174
rect 17832 27172 17856 27174
rect 17912 27172 17918 27174
rect 17610 27163 17918 27172
rect 22610 27228 22918 27237
rect 22610 27226 22616 27228
rect 22672 27226 22696 27228
rect 22752 27226 22776 27228
rect 22832 27226 22856 27228
rect 22912 27226 22918 27228
rect 22672 27174 22674 27226
rect 22854 27174 22856 27226
rect 22610 27172 22616 27174
rect 22672 27172 22696 27174
rect 22752 27172 22776 27174
rect 22832 27172 22856 27174
rect 22912 27172 22918 27174
rect 22610 27163 22918 27172
rect 27610 27228 27918 27237
rect 27610 27226 27616 27228
rect 27672 27226 27696 27228
rect 27752 27226 27776 27228
rect 27832 27226 27856 27228
rect 27912 27226 27918 27228
rect 27672 27174 27674 27226
rect 27854 27174 27856 27226
rect 27610 27172 27616 27174
rect 27672 27172 27696 27174
rect 27752 27172 27776 27174
rect 27832 27172 27856 27174
rect 27912 27172 27918 27174
rect 27610 27163 27918 27172
rect 32610 27228 32918 27237
rect 32610 27226 32616 27228
rect 32672 27226 32696 27228
rect 32752 27226 32776 27228
rect 32832 27226 32856 27228
rect 32912 27226 32918 27228
rect 32672 27174 32674 27226
rect 32854 27174 32856 27226
rect 32610 27172 32616 27174
rect 32672 27172 32696 27174
rect 32752 27172 32776 27174
rect 32832 27172 32856 27174
rect 32912 27172 32918 27174
rect 32610 27163 32918 27172
rect 37610 27228 37918 27237
rect 37610 27226 37616 27228
rect 37672 27226 37696 27228
rect 37752 27226 37776 27228
rect 37832 27226 37856 27228
rect 37912 27226 37918 27228
rect 37672 27174 37674 27226
rect 37854 27174 37856 27226
rect 37610 27172 37616 27174
rect 37672 27172 37696 27174
rect 37752 27172 37776 27174
rect 37832 27172 37856 27174
rect 37912 27172 37918 27174
rect 37610 27163 37918 27172
rect 42610 27228 42918 27237
rect 42610 27226 42616 27228
rect 42672 27226 42696 27228
rect 42752 27226 42776 27228
rect 42832 27226 42856 27228
rect 42912 27226 42918 27228
rect 42672 27174 42674 27226
rect 42854 27174 42856 27226
rect 42610 27172 42616 27174
rect 42672 27172 42696 27174
rect 42752 27172 42776 27174
rect 42832 27172 42856 27174
rect 42912 27172 42918 27174
rect 42610 27163 42918 27172
rect 47610 27228 47918 27237
rect 47610 27226 47616 27228
rect 47672 27226 47696 27228
rect 47752 27226 47776 27228
rect 47832 27226 47856 27228
rect 47912 27226 47918 27228
rect 47672 27174 47674 27226
rect 47854 27174 47856 27226
rect 47610 27172 47616 27174
rect 47672 27172 47696 27174
rect 47752 27172 47776 27174
rect 47832 27172 47856 27174
rect 47912 27172 47918 27174
rect 47610 27163 47918 27172
rect 52610 27228 52918 27237
rect 52610 27226 52616 27228
rect 52672 27226 52696 27228
rect 52752 27226 52776 27228
rect 52832 27226 52856 27228
rect 52912 27226 52918 27228
rect 52672 27174 52674 27226
rect 52854 27174 52856 27226
rect 52610 27172 52616 27174
rect 52672 27172 52696 27174
rect 52752 27172 52776 27174
rect 52832 27172 52856 27174
rect 52912 27172 52918 27174
rect 52610 27163 52918 27172
rect 57610 27228 57918 27237
rect 57610 27226 57616 27228
rect 57672 27226 57696 27228
rect 57752 27226 57776 27228
rect 57832 27226 57856 27228
rect 57912 27226 57918 27228
rect 57672 27174 57674 27226
rect 57854 27174 57856 27226
rect 57610 27172 57616 27174
rect 57672 27172 57696 27174
rect 57752 27172 57776 27174
rect 57832 27172 57856 27174
rect 57912 27172 57918 27174
rect 57610 27163 57918 27172
rect 58544 27033 58572 27406
rect 58530 27024 58586 27033
rect 58530 26959 58586 26968
rect 1950 26684 2258 26693
rect 1950 26682 1956 26684
rect 2012 26682 2036 26684
rect 2092 26682 2116 26684
rect 2172 26682 2196 26684
rect 2252 26682 2258 26684
rect 2012 26630 2014 26682
rect 2194 26630 2196 26682
rect 1950 26628 1956 26630
rect 2012 26628 2036 26630
rect 2092 26628 2116 26630
rect 2172 26628 2196 26630
rect 2252 26628 2258 26630
rect 1950 26619 2258 26628
rect 6950 26684 7258 26693
rect 6950 26682 6956 26684
rect 7012 26682 7036 26684
rect 7092 26682 7116 26684
rect 7172 26682 7196 26684
rect 7252 26682 7258 26684
rect 7012 26630 7014 26682
rect 7194 26630 7196 26682
rect 6950 26628 6956 26630
rect 7012 26628 7036 26630
rect 7092 26628 7116 26630
rect 7172 26628 7196 26630
rect 7252 26628 7258 26630
rect 6950 26619 7258 26628
rect 11950 26684 12258 26693
rect 11950 26682 11956 26684
rect 12012 26682 12036 26684
rect 12092 26682 12116 26684
rect 12172 26682 12196 26684
rect 12252 26682 12258 26684
rect 12012 26630 12014 26682
rect 12194 26630 12196 26682
rect 11950 26628 11956 26630
rect 12012 26628 12036 26630
rect 12092 26628 12116 26630
rect 12172 26628 12196 26630
rect 12252 26628 12258 26630
rect 11950 26619 12258 26628
rect 16950 26684 17258 26693
rect 16950 26682 16956 26684
rect 17012 26682 17036 26684
rect 17092 26682 17116 26684
rect 17172 26682 17196 26684
rect 17252 26682 17258 26684
rect 17012 26630 17014 26682
rect 17194 26630 17196 26682
rect 16950 26628 16956 26630
rect 17012 26628 17036 26630
rect 17092 26628 17116 26630
rect 17172 26628 17196 26630
rect 17252 26628 17258 26630
rect 16950 26619 17258 26628
rect 21950 26684 22258 26693
rect 21950 26682 21956 26684
rect 22012 26682 22036 26684
rect 22092 26682 22116 26684
rect 22172 26682 22196 26684
rect 22252 26682 22258 26684
rect 22012 26630 22014 26682
rect 22194 26630 22196 26682
rect 21950 26628 21956 26630
rect 22012 26628 22036 26630
rect 22092 26628 22116 26630
rect 22172 26628 22196 26630
rect 22252 26628 22258 26630
rect 21950 26619 22258 26628
rect 26950 26684 27258 26693
rect 26950 26682 26956 26684
rect 27012 26682 27036 26684
rect 27092 26682 27116 26684
rect 27172 26682 27196 26684
rect 27252 26682 27258 26684
rect 27012 26630 27014 26682
rect 27194 26630 27196 26682
rect 26950 26628 26956 26630
rect 27012 26628 27036 26630
rect 27092 26628 27116 26630
rect 27172 26628 27196 26630
rect 27252 26628 27258 26630
rect 26950 26619 27258 26628
rect 31950 26684 32258 26693
rect 31950 26682 31956 26684
rect 32012 26682 32036 26684
rect 32092 26682 32116 26684
rect 32172 26682 32196 26684
rect 32252 26682 32258 26684
rect 32012 26630 32014 26682
rect 32194 26630 32196 26682
rect 31950 26628 31956 26630
rect 32012 26628 32036 26630
rect 32092 26628 32116 26630
rect 32172 26628 32196 26630
rect 32252 26628 32258 26630
rect 31950 26619 32258 26628
rect 36950 26684 37258 26693
rect 36950 26682 36956 26684
rect 37012 26682 37036 26684
rect 37092 26682 37116 26684
rect 37172 26682 37196 26684
rect 37252 26682 37258 26684
rect 37012 26630 37014 26682
rect 37194 26630 37196 26682
rect 36950 26628 36956 26630
rect 37012 26628 37036 26630
rect 37092 26628 37116 26630
rect 37172 26628 37196 26630
rect 37252 26628 37258 26630
rect 36950 26619 37258 26628
rect 41950 26684 42258 26693
rect 41950 26682 41956 26684
rect 42012 26682 42036 26684
rect 42092 26682 42116 26684
rect 42172 26682 42196 26684
rect 42252 26682 42258 26684
rect 42012 26630 42014 26682
rect 42194 26630 42196 26682
rect 41950 26628 41956 26630
rect 42012 26628 42036 26630
rect 42092 26628 42116 26630
rect 42172 26628 42196 26630
rect 42252 26628 42258 26630
rect 41950 26619 42258 26628
rect 46950 26684 47258 26693
rect 46950 26682 46956 26684
rect 47012 26682 47036 26684
rect 47092 26682 47116 26684
rect 47172 26682 47196 26684
rect 47252 26682 47258 26684
rect 47012 26630 47014 26682
rect 47194 26630 47196 26682
rect 46950 26628 46956 26630
rect 47012 26628 47036 26630
rect 47092 26628 47116 26630
rect 47172 26628 47196 26630
rect 47252 26628 47258 26630
rect 46950 26619 47258 26628
rect 51950 26684 52258 26693
rect 51950 26682 51956 26684
rect 52012 26682 52036 26684
rect 52092 26682 52116 26684
rect 52172 26682 52196 26684
rect 52252 26682 52258 26684
rect 52012 26630 52014 26682
rect 52194 26630 52196 26682
rect 51950 26628 51956 26630
rect 52012 26628 52036 26630
rect 52092 26628 52116 26630
rect 52172 26628 52196 26630
rect 52252 26628 52258 26630
rect 51950 26619 52258 26628
rect 56950 26684 57258 26693
rect 56950 26682 56956 26684
rect 57012 26682 57036 26684
rect 57092 26682 57116 26684
rect 57172 26682 57196 26684
rect 57252 26682 57258 26684
rect 57012 26630 57014 26682
rect 57194 26630 57196 26682
rect 56950 26628 56956 26630
rect 57012 26628 57036 26630
rect 57092 26628 57116 26630
rect 57172 26628 57196 26630
rect 57252 26628 57258 26630
rect 56950 26619 57258 26628
rect 58348 26376 58400 26382
rect 58348 26318 58400 26324
rect 58360 26217 58388 26318
rect 58346 26208 58402 26217
rect 2610 26140 2918 26149
rect 2610 26138 2616 26140
rect 2672 26138 2696 26140
rect 2752 26138 2776 26140
rect 2832 26138 2856 26140
rect 2912 26138 2918 26140
rect 2672 26086 2674 26138
rect 2854 26086 2856 26138
rect 2610 26084 2616 26086
rect 2672 26084 2696 26086
rect 2752 26084 2776 26086
rect 2832 26084 2856 26086
rect 2912 26084 2918 26086
rect 2610 26075 2918 26084
rect 7610 26140 7918 26149
rect 7610 26138 7616 26140
rect 7672 26138 7696 26140
rect 7752 26138 7776 26140
rect 7832 26138 7856 26140
rect 7912 26138 7918 26140
rect 7672 26086 7674 26138
rect 7854 26086 7856 26138
rect 7610 26084 7616 26086
rect 7672 26084 7696 26086
rect 7752 26084 7776 26086
rect 7832 26084 7856 26086
rect 7912 26084 7918 26086
rect 7610 26075 7918 26084
rect 12610 26140 12918 26149
rect 12610 26138 12616 26140
rect 12672 26138 12696 26140
rect 12752 26138 12776 26140
rect 12832 26138 12856 26140
rect 12912 26138 12918 26140
rect 12672 26086 12674 26138
rect 12854 26086 12856 26138
rect 12610 26084 12616 26086
rect 12672 26084 12696 26086
rect 12752 26084 12776 26086
rect 12832 26084 12856 26086
rect 12912 26084 12918 26086
rect 12610 26075 12918 26084
rect 17610 26140 17918 26149
rect 17610 26138 17616 26140
rect 17672 26138 17696 26140
rect 17752 26138 17776 26140
rect 17832 26138 17856 26140
rect 17912 26138 17918 26140
rect 17672 26086 17674 26138
rect 17854 26086 17856 26138
rect 17610 26084 17616 26086
rect 17672 26084 17696 26086
rect 17752 26084 17776 26086
rect 17832 26084 17856 26086
rect 17912 26084 17918 26086
rect 17610 26075 17918 26084
rect 22610 26140 22918 26149
rect 22610 26138 22616 26140
rect 22672 26138 22696 26140
rect 22752 26138 22776 26140
rect 22832 26138 22856 26140
rect 22912 26138 22918 26140
rect 22672 26086 22674 26138
rect 22854 26086 22856 26138
rect 22610 26084 22616 26086
rect 22672 26084 22696 26086
rect 22752 26084 22776 26086
rect 22832 26084 22856 26086
rect 22912 26084 22918 26086
rect 22610 26075 22918 26084
rect 27610 26140 27918 26149
rect 27610 26138 27616 26140
rect 27672 26138 27696 26140
rect 27752 26138 27776 26140
rect 27832 26138 27856 26140
rect 27912 26138 27918 26140
rect 27672 26086 27674 26138
rect 27854 26086 27856 26138
rect 27610 26084 27616 26086
rect 27672 26084 27696 26086
rect 27752 26084 27776 26086
rect 27832 26084 27856 26086
rect 27912 26084 27918 26086
rect 27610 26075 27918 26084
rect 32610 26140 32918 26149
rect 32610 26138 32616 26140
rect 32672 26138 32696 26140
rect 32752 26138 32776 26140
rect 32832 26138 32856 26140
rect 32912 26138 32918 26140
rect 32672 26086 32674 26138
rect 32854 26086 32856 26138
rect 32610 26084 32616 26086
rect 32672 26084 32696 26086
rect 32752 26084 32776 26086
rect 32832 26084 32856 26086
rect 32912 26084 32918 26086
rect 32610 26075 32918 26084
rect 37610 26140 37918 26149
rect 37610 26138 37616 26140
rect 37672 26138 37696 26140
rect 37752 26138 37776 26140
rect 37832 26138 37856 26140
rect 37912 26138 37918 26140
rect 37672 26086 37674 26138
rect 37854 26086 37856 26138
rect 37610 26084 37616 26086
rect 37672 26084 37696 26086
rect 37752 26084 37776 26086
rect 37832 26084 37856 26086
rect 37912 26084 37918 26086
rect 37610 26075 37918 26084
rect 42610 26140 42918 26149
rect 42610 26138 42616 26140
rect 42672 26138 42696 26140
rect 42752 26138 42776 26140
rect 42832 26138 42856 26140
rect 42912 26138 42918 26140
rect 42672 26086 42674 26138
rect 42854 26086 42856 26138
rect 42610 26084 42616 26086
rect 42672 26084 42696 26086
rect 42752 26084 42776 26086
rect 42832 26084 42856 26086
rect 42912 26084 42918 26086
rect 42610 26075 42918 26084
rect 47610 26140 47918 26149
rect 47610 26138 47616 26140
rect 47672 26138 47696 26140
rect 47752 26138 47776 26140
rect 47832 26138 47856 26140
rect 47912 26138 47918 26140
rect 47672 26086 47674 26138
rect 47854 26086 47856 26138
rect 47610 26084 47616 26086
rect 47672 26084 47696 26086
rect 47752 26084 47776 26086
rect 47832 26084 47856 26086
rect 47912 26084 47918 26086
rect 47610 26075 47918 26084
rect 52610 26140 52918 26149
rect 52610 26138 52616 26140
rect 52672 26138 52696 26140
rect 52752 26138 52776 26140
rect 52832 26138 52856 26140
rect 52912 26138 52918 26140
rect 52672 26086 52674 26138
rect 52854 26086 52856 26138
rect 52610 26084 52616 26086
rect 52672 26084 52696 26086
rect 52752 26084 52776 26086
rect 52832 26084 52856 26086
rect 52912 26084 52918 26086
rect 52610 26075 52918 26084
rect 57610 26140 57918 26149
rect 58346 26143 58402 26152
rect 57610 26138 57616 26140
rect 57672 26138 57696 26140
rect 57752 26138 57776 26140
rect 57832 26138 57856 26140
rect 57912 26138 57918 26140
rect 57672 26086 57674 26138
rect 57854 26086 57856 26138
rect 57610 26084 57616 26086
rect 57672 26084 57696 26086
rect 57752 26084 57776 26086
rect 57832 26084 57856 26086
rect 57912 26084 57918 26086
rect 57610 26075 57918 26084
rect 58532 25696 58584 25702
rect 58532 25638 58584 25644
rect 1950 25596 2258 25605
rect 1950 25594 1956 25596
rect 2012 25594 2036 25596
rect 2092 25594 2116 25596
rect 2172 25594 2196 25596
rect 2252 25594 2258 25596
rect 2012 25542 2014 25594
rect 2194 25542 2196 25594
rect 1950 25540 1956 25542
rect 2012 25540 2036 25542
rect 2092 25540 2116 25542
rect 2172 25540 2196 25542
rect 2252 25540 2258 25542
rect 1950 25531 2258 25540
rect 6950 25596 7258 25605
rect 6950 25594 6956 25596
rect 7012 25594 7036 25596
rect 7092 25594 7116 25596
rect 7172 25594 7196 25596
rect 7252 25594 7258 25596
rect 7012 25542 7014 25594
rect 7194 25542 7196 25594
rect 6950 25540 6956 25542
rect 7012 25540 7036 25542
rect 7092 25540 7116 25542
rect 7172 25540 7196 25542
rect 7252 25540 7258 25542
rect 6950 25531 7258 25540
rect 11950 25596 12258 25605
rect 11950 25594 11956 25596
rect 12012 25594 12036 25596
rect 12092 25594 12116 25596
rect 12172 25594 12196 25596
rect 12252 25594 12258 25596
rect 12012 25542 12014 25594
rect 12194 25542 12196 25594
rect 11950 25540 11956 25542
rect 12012 25540 12036 25542
rect 12092 25540 12116 25542
rect 12172 25540 12196 25542
rect 12252 25540 12258 25542
rect 11950 25531 12258 25540
rect 16950 25596 17258 25605
rect 16950 25594 16956 25596
rect 17012 25594 17036 25596
rect 17092 25594 17116 25596
rect 17172 25594 17196 25596
rect 17252 25594 17258 25596
rect 17012 25542 17014 25594
rect 17194 25542 17196 25594
rect 16950 25540 16956 25542
rect 17012 25540 17036 25542
rect 17092 25540 17116 25542
rect 17172 25540 17196 25542
rect 17252 25540 17258 25542
rect 16950 25531 17258 25540
rect 21950 25596 22258 25605
rect 21950 25594 21956 25596
rect 22012 25594 22036 25596
rect 22092 25594 22116 25596
rect 22172 25594 22196 25596
rect 22252 25594 22258 25596
rect 22012 25542 22014 25594
rect 22194 25542 22196 25594
rect 21950 25540 21956 25542
rect 22012 25540 22036 25542
rect 22092 25540 22116 25542
rect 22172 25540 22196 25542
rect 22252 25540 22258 25542
rect 21950 25531 22258 25540
rect 26950 25596 27258 25605
rect 26950 25594 26956 25596
rect 27012 25594 27036 25596
rect 27092 25594 27116 25596
rect 27172 25594 27196 25596
rect 27252 25594 27258 25596
rect 27012 25542 27014 25594
rect 27194 25542 27196 25594
rect 26950 25540 26956 25542
rect 27012 25540 27036 25542
rect 27092 25540 27116 25542
rect 27172 25540 27196 25542
rect 27252 25540 27258 25542
rect 26950 25531 27258 25540
rect 31950 25596 32258 25605
rect 31950 25594 31956 25596
rect 32012 25594 32036 25596
rect 32092 25594 32116 25596
rect 32172 25594 32196 25596
rect 32252 25594 32258 25596
rect 32012 25542 32014 25594
rect 32194 25542 32196 25594
rect 31950 25540 31956 25542
rect 32012 25540 32036 25542
rect 32092 25540 32116 25542
rect 32172 25540 32196 25542
rect 32252 25540 32258 25542
rect 31950 25531 32258 25540
rect 36950 25596 37258 25605
rect 36950 25594 36956 25596
rect 37012 25594 37036 25596
rect 37092 25594 37116 25596
rect 37172 25594 37196 25596
rect 37252 25594 37258 25596
rect 37012 25542 37014 25594
rect 37194 25542 37196 25594
rect 36950 25540 36956 25542
rect 37012 25540 37036 25542
rect 37092 25540 37116 25542
rect 37172 25540 37196 25542
rect 37252 25540 37258 25542
rect 36950 25531 37258 25540
rect 41950 25596 42258 25605
rect 41950 25594 41956 25596
rect 42012 25594 42036 25596
rect 42092 25594 42116 25596
rect 42172 25594 42196 25596
rect 42252 25594 42258 25596
rect 42012 25542 42014 25594
rect 42194 25542 42196 25594
rect 41950 25540 41956 25542
rect 42012 25540 42036 25542
rect 42092 25540 42116 25542
rect 42172 25540 42196 25542
rect 42252 25540 42258 25542
rect 41950 25531 42258 25540
rect 46950 25596 47258 25605
rect 46950 25594 46956 25596
rect 47012 25594 47036 25596
rect 47092 25594 47116 25596
rect 47172 25594 47196 25596
rect 47252 25594 47258 25596
rect 47012 25542 47014 25594
rect 47194 25542 47196 25594
rect 46950 25540 46956 25542
rect 47012 25540 47036 25542
rect 47092 25540 47116 25542
rect 47172 25540 47196 25542
rect 47252 25540 47258 25542
rect 46950 25531 47258 25540
rect 51950 25596 52258 25605
rect 51950 25594 51956 25596
rect 52012 25594 52036 25596
rect 52092 25594 52116 25596
rect 52172 25594 52196 25596
rect 52252 25594 52258 25596
rect 52012 25542 52014 25594
rect 52194 25542 52196 25594
rect 51950 25540 51956 25542
rect 52012 25540 52036 25542
rect 52092 25540 52116 25542
rect 52172 25540 52196 25542
rect 52252 25540 52258 25542
rect 51950 25531 52258 25540
rect 56950 25596 57258 25605
rect 56950 25594 56956 25596
rect 57012 25594 57036 25596
rect 57092 25594 57116 25596
rect 57172 25594 57196 25596
rect 57252 25594 57258 25596
rect 57012 25542 57014 25594
rect 57194 25542 57196 25594
rect 56950 25540 56956 25542
rect 57012 25540 57036 25542
rect 57092 25540 57116 25542
rect 57172 25540 57196 25542
rect 57252 25540 57258 25542
rect 56950 25531 57258 25540
rect 58544 25401 58572 25638
rect 58530 25392 58586 25401
rect 58530 25327 58586 25336
rect 2610 25052 2918 25061
rect 2610 25050 2616 25052
rect 2672 25050 2696 25052
rect 2752 25050 2776 25052
rect 2832 25050 2856 25052
rect 2912 25050 2918 25052
rect 2672 24998 2674 25050
rect 2854 24998 2856 25050
rect 2610 24996 2616 24998
rect 2672 24996 2696 24998
rect 2752 24996 2776 24998
rect 2832 24996 2856 24998
rect 2912 24996 2918 24998
rect 2610 24987 2918 24996
rect 7610 25052 7918 25061
rect 7610 25050 7616 25052
rect 7672 25050 7696 25052
rect 7752 25050 7776 25052
rect 7832 25050 7856 25052
rect 7912 25050 7918 25052
rect 7672 24998 7674 25050
rect 7854 24998 7856 25050
rect 7610 24996 7616 24998
rect 7672 24996 7696 24998
rect 7752 24996 7776 24998
rect 7832 24996 7856 24998
rect 7912 24996 7918 24998
rect 7610 24987 7918 24996
rect 12610 25052 12918 25061
rect 12610 25050 12616 25052
rect 12672 25050 12696 25052
rect 12752 25050 12776 25052
rect 12832 25050 12856 25052
rect 12912 25050 12918 25052
rect 12672 24998 12674 25050
rect 12854 24998 12856 25050
rect 12610 24996 12616 24998
rect 12672 24996 12696 24998
rect 12752 24996 12776 24998
rect 12832 24996 12856 24998
rect 12912 24996 12918 24998
rect 12610 24987 12918 24996
rect 17610 25052 17918 25061
rect 17610 25050 17616 25052
rect 17672 25050 17696 25052
rect 17752 25050 17776 25052
rect 17832 25050 17856 25052
rect 17912 25050 17918 25052
rect 17672 24998 17674 25050
rect 17854 24998 17856 25050
rect 17610 24996 17616 24998
rect 17672 24996 17696 24998
rect 17752 24996 17776 24998
rect 17832 24996 17856 24998
rect 17912 24996 17918 24998
rect 17610 24987 17918 24996
rect 22610 25052 22918 25061
rect 22610 25050 22616 25052
rect 22672 25050 22696 25052
rect 22752 25050 22776 25052
rect 22832 25050 22856 25052
rect 22912 25050 22918 25052
rect 22672 24998 22674 25050
rect 22854 24998 22856 25050
rect 22610 24996 22616 24998
rect 22672 24996 22696 24998
rect 22752 24996 22776 24998
rect 22832 24996 22856 24998
rect 22912 24996 22918 24998
rect 22610 24987 22918 24996
rect 27610 25052 27918 25061
rect 27610 25050 27616 25052
rect 27672 25050 27696 25052
rect 27752 25050 27776 25052
rect 27832 25050 27856 25052
rect 27912 25050 27918 25052
rect 27672 24998 27674 25050
rect 27854 24998 27856 25050
rect 27610 24996 27616 24998
rect 27672 24996 27696 24998
rect 27752 24996 27776 24998
rect 27832 24996 27856 24998
rect 27912 24996 27918 24998
rect 27610 24987 27918 24996
rect 32610 25052 32918 25061
rect 32610 25050 32616 25052
rect 32672 25050 32696 25052
rect 32752 25050 32776 25052
rect 32832 25050 32856 25052
rect 32912 25050 32918 25052
rect 32672 24998 32674 25050
rect 32854 24998 32856 25050
rect 32610 24996 32616 24998
rect 32672 24996 32696 24998
rect 32752 24996 32776 24998
rect 32832 24996 32856 24998
rect 32912 24996 32918 24998
rect 32610 24987 32918 24996
rect 37610 25052 37918 25061
rect 37610 25050 37616 25052
rect 37672 25050 37696 25052
rect 37752 25050 37776 25052
rect 37832 25050 37856 25052
rect 37912 25050 37918 25052
rect 37672 24998 37674 25050
rect 37854 24998 37856 25050
rect 37610 24996 37616 24998
rect 37672 24996 37696 24998
rect 37752 24996 37776 24998
rect 37832 24996 37856 24998
rect 37912 24996 37918 24998
rect 37610 24987 37918 24996
rect 42610 25052 42918 25061
rect 42610 25050 42616 25052
rect 42672 25050 42696 25052
rect 42752 25050 42776 25052
rect 42832 25050 42856 25052
rect 42912 25050 42918 25052
rect 42672 24998 42674 25050
rect 42854 24998 42856 25050
rect 42610 24996 42616 24998
rect 42672 24996 42696 24998
rect 42752 24996 42776 24998
rect 42832 24996 42856 24998
rect 42912 24996 42918 24998
rect 42610 24987 42918 24996
rect 47610 25052 47918 25061
rect 47610 25050 47616 25052
rect 47672 25050 47696 25052
rect 47752 25050 47776 25052
rect 47832 25050 47856 25052
rect 47912 25050 47918 25052
rect 47672 24998 47674 25050
rect 47854 24998 47856 25050
rect 47610 24996 47616 24998
rect 47672 24996 47696 24998
rect 47752 24996 47776 24998
rect 47832 24996 47856 24998
rect 47912 24996 47918 24998
rect 47610 24987 47918 24996
rect 52610 25052 52918 25061
rect 52610 25050 52616 25052
rect 52672 25050 52696 25052
rect 52752 25050 52776 25052
rect 52832 25050 52856 25052
rect 52912 25050 52918 25052
rect 52672 24998 52674 25050
rect 52854 24998 52856 25050
rect 52610 24996 52616 24998
rect 52672 24996 52696 24998
rect 52752 24996 52776 24998
rect 52832 24996 52856 24998
rect 52912 24996 52918 24998
rect 52610 24987 52918 24996
rect 57610 25052 57918 25061
rect 57610 25050 57616 25052
rect 57672 25050 57696 25052
rect 57752 25050 57776 25052
rect 57832 25050 57856 25052
rect 57912 25050 57918 25052
rect 57672 24998 57674 25050
rect 57854 24998 57856 25050
rect 57610 24996 57616 24998
rect 57672 24996 57696 24998
rect 57752 24996 57776 24998
rect 57832 24996 57856 24998
rect 57912 24996 57918 24998
rect 57610 24987 57918 24996
rect 58532 24608 58584 24614
rect 58530 24576 58532 24585
rect 58584 24576 58586 24585
rect 1950 24508 2258 24517
rect 1950 24506 1956 24508
rect 2012 24506 2036 24508
rect 2092 24506 2116 24508
rect 2172 24506 2196 24508
rect 2252 24506 2258 24508
rect 2012 24454 2014 24506
rect 2194 24454 2196 24506
rect 1950 24452 1956 24454
rect 2012 24452 2036 24454
rect 2092 24452 2116 24454
rect 2172 24452 2196 24454
rect 2252 24452 2258 24454
rect 1950 24443 2258 24452
rect 6950 24508 7258 24517
rect 6950 24506 6956 24508
rect 7012 24506 7036 24508
rect 7092 24506 7116 24508
rect 7172 24506 7196 24508
rect 7252 24506 7258 24508
rect 7012 24454 7014 24506
rect 7194 24454 7196 24506
rect 6950 24452 6956 24454
rect 7012 24452 7036 24454
rect 7092 24452 7116 24454
rect 7172 24452 7196 24454
rect 7252 24452 7258 24454
rect 6950 24443 7258 24452
rect 11950 24508 12258 24517
rect 11950 24506 11956 24508
rect 12012 24506 12036 24508
rect 12092 24506 12116 24508
rect 12172 24506 12196 24508
rect 12252 24506 12258 24508
rect 12012 24454 12014 24506
rect 12194 24454 12196 24506
rect 11950 24452 11956 24454
rect 12012 24452 12036 24454
rect 12092 24452 12116 24454
rect 12172 24452 12196 24454
rect 12252 24452 12258 24454
rect 11950 24443 12258 24452
rect 16950 24508 17258 24517
rect 16950 24506 16956 24508
rect 17012 24506 17036 24508
rect 17092 24506 17116 24508
rect 17172 24506 17196 24508
rect 17252 24506 17258 24508
rect 17012 24454 17014 24506
rect 17194 24454 17196 24506
rect 16950 24452 16956 24454
rect 17012 24452 17036 24454
rect 17092 24452 17116 24454
rect 17172 24452 17196 24454
rect 17252 24452 17258 24454
rect 16950 24443 17258 24452
rect 21950 24508 22258 24517
rect 21950 24506 21956 24508
rect 22012 24506 22036 24508
rect 22092 24506 22116 24508
rect 22172 24506 22196 24508
rect 22252 24506 22258 24508
rect 22012 24454 22014 24506
rect 22194 24454 22196 24506
rect 21950 24452 21956 24454
rect 22012 24452 22036 24454
rect 22092 24452 22116 24454
rect 22172 24452 22196 24454
rect 22252 24452 22258 24454
rect 21950 24443 22258 24452
rect 26950 24508 27258 24517
rect 26950 24506 26956 24508
rect 27012 24506 27036 24508
rect 27092 24506 27116 24508
rect 27172 24506 27196 24508
rect 27252 24506 27258 24508
rect 27012 24454 27014 24506
rect 27194 24454 27196 24506
rect 26950 24452 26956 24454
rect 27012 24452 27036 24454
rect 27092 24452 27116 24454
rect 27172 24452 27196 24454
rect 27252 24452 27258 24454
rect 26950 24443 27258 24452
rect 31950 24508 32258 24517
rect 31950 24506 31956 24508
rect 32012 24506 32036 24508
rect 32092 24506 32116 24508
rect 32172 24506 32196 24508
rect 32252 24506 32258 24508
rect 32012 24454 32014 24506
rect 32194 24454 32196 24506
rect 31950 24452 31956 24454
rect 32012 24452 32036 24454
rect 32092 24452 32116 24454
rect 32172 24452 32196 24454
rect 32252 24452 32258 24454
rect 31950 24443 32258 24452
rect 36950 24508 37258 24517
rect 36950 24506 36956 24508
rect 37012 24506 37036 24508
rect 37092 24506 37116 24508
rect 37172 24506 37196 24508
rect 37252 24506 37258 24508
rect 37012 24454 37014 24506
rect 37194 24454 37196 24506
rect 36950 24452 36956 24454
rect 37012 24452 37036 24454
rect 37092 24452 37116 24454
rect 37172 24452 37196 24454
rect 37252 24452 37258 24454
rect 36950 24443 37258 24452
rect 41950 24508 42258 24517
rect 41950 24506 41956 24508
rect 42012 24506 42036 24508
rect 42092 24506 42116 24508
rect 42172 24506 42196 24508
rect 42252 24506 42258 24508
rect 42012 24454 42014 24506
rect 42194 24454 42196 24506
rect 41950 24452 41956 24454
rect 42012 24452 42036 24454
rect 42092 24452 42116 24454
rect 42172 24452 42196 24454
rect 42252 24452 42258 24454
rect 41950 24443 42258 24452
rect 46950 24508 47258 24517
rect 46950 24506 46956 24508
rect 47012 24506 47036 24508
rect 47092 24506 47116 24508
rect 47172 24506 47196 24508
rect 47252 24506 47258 24508
rect 47012 24454 47014 24506
rect 47194 24454 47196 24506
rect 46950 24452 46956 24454
rect 47012 24452 47036 24454
rect 47092 24452 47116 24454
rect 47172 24452 47196 24454
rect 47252 24452 47258 24454
rect 46950 24443 47258 24452
rect 51950 24508 52258 24517
rect 51950 24506 51956 24508
rect 52012 24506 52036 24508
rect 52092 24506 52116 24508
rect 52172 24506 52196 24508
rect 52252 24506 52258 24508
rect 52012 24454 52014 24506
rect 52194 24454 52196 24506
rect 51950 24452 51956 24454
rect 52012 24452 52036 24454
rect 52092 24452 52116 24454
rect 52172 24452 52196 24454
rect 52252 24452 52258 24454
rect 51950 24443 52258 24452
rect 56950 24508 57258 24517
rect 58530 24511 58586 24520
rect 56950 24506 56956 24508
rect 57012 24506 57036 24508
rect 57092 24506 57116 24508
rect 57172 24506 57196 24508
rect 57252 24506 57258 24508
rect 57012 24454 57014 24506
rect 57194 24454 57196 24506
rect 56950 24452 56956 24454
rect 57012 24452 57036 24454
rect 57092 24452 57116 24454
rect 57172 24452 57196 24454
rect 57252 24452 57258 24454
rect 56950 24443 57258 24452
rect 58532 24200 58584 24206
rect 58532 24142 58584 24148
rect 2610 23964 2918 23973
rect 2610 23962 2616 23964
rect 2672 23962 2696 23964
rect 2752 23962 2776 23964
rect 2832 23962 2856 23964
rect 2912 23962 2918 23964
rect 2672 23910 2674 23962
rect 2854 23910 2856 23962
rect 2610 23908 2616 23910
rect 2672 23908 2696 23910
rect 2752 23908 2776 23910
rect 2832 23908 2856 23910
rect 2912 23908 2918 23910
rect 2610 23899 2918 23908
rect 7610 23964 7918 23973
rect 7610 23962 7616 23964
rect 7672 23962 7696 23964
rect 7752 23962 7776 23964
rect 7832 23962 7856 23964
rect 7912 23962 7918 23964
rect 7672 23910 7674 23962
rect 7854 23910 7856 23962
rect 7610 23908 7616 23910
rect 7672 23908 7696 23910
rect 7752 23908 7776 23910
rect 7832 23908 7856 23910
rect 7912 23908 7918 23910
rect 7610 23899 7918 23908
rect 12610 23964 12918 23973
rect 12610 23962 12616 23964
rect 12672 23962 12696 23964
rect 12752 23962 12776 23964
rect 12832 23962 12856 23964
rect 12912 23962 12918 23964
rect 12672 23910 12674 23962
rect 12854 23910 12856 23962
rect 12610 23908 12616 23910
rect 12672 23908 12696 23910
rect 12752 23908 12776 23910
rect 12832 23908 12856 23910
rect 12912 23908 12918 23910
rect 12610 23899 12918 23908
rect 17610 23964 17918 23973
rect 17610 23962 17616 23964
rect 17672 23962 17696 23964
rect 17752 23962 17776 23964
rect 17832 23962 17856 23964
rect 17912 23962 17918 23964
rect 17672 23910 17674 23962
rect 17854 23910 17856 23962
rect 17610 23908 17616 23910
rect 17672 23908 17696 23910
rect 17752 23908 17776 23910
rect 17832 23908 17856 23910
rect 17912 23908 17918 23910
rect 17610 23899 17918 23908
rect 22610 23964 22918 23973
rect 22610 23962 22616 23964
rect 22672 23962 22696 23964
rect 22752 23962 22776 23964
rect 22832 23962 22856 23964
rect 22912 23962 22918 23964
rect 22672 23910 22674 23962
rect 22854 23910 22856 23962
rect 22610 23908 22616 23910
rect 22672 23908 22696 23910
rect 22752 23908 22776 23910
rect 22832 23908 22856 23910
rect 22912 23908 22918 23910
rect 22610 23899 22918 23908
rect 27610 23964 27918 23973
rect 27610 23962 27616 23964
rect 27672 23962 27696 23964
rect 27752 23962 27776 23964
rect 27832 23962 27856 23964
rect 27912 23962 27918 23964
rect 27672 23910 27674 23962
rect 27854 23910 27856 23962
rect 27610 23908 27616 23910
rect 27672 23908 27696 23910
rect 27752 23908 27776 23910
rect 27832 23908 27856 23910
rect 27912 23908 27918 23910
rect 27610 23899 27918 23908
rect 32610 23964 32918 23973
rect 32610 23962 32616 23964
rect 32672 23962 32696 23964
rect 32752 23962 32776 23964
rect 32832 23962 32856 23964
rect 32912 23962 32918 23964
rect 32672 23910 32674 23962
rect 32854 23910 32856 23962
rect 32610 23908 32616 23910
rect 32672 23908 32696 23910
rect 32752 23908 32776 23910
rect 32832 23908 32856 23910
rect 32912 23908 32918 23910
rect 32610 23899 32918 23908
rect 37610 23964 37918 23973
rect 37610 23962 37616 23964
rect 37672 23962 37696 23964
rect 37752 23962 37776 23964
rect 37832 23962 37856 23964
rect 37912 23962 37918 23964
rect 37672 23910 37674 23962
rect 37854 23910 37856 23962
rect 37610 23908 37616 23910
rect 37672 23908 37696 23910
rect 37752 23908 37776 23910
rect 37832 23908 37856 23910
rect 37912 23908 37918 23910
rect 37610 23899 37918 23908
rect 42610 23964 42918 23973
rect 42610 23962 42616 23964
rect 42672 23962 42696 23964
rect 42752 23962 42776 23964
rect 42832 23962 42856 23964
rect 42912 23962 42918 23964
rect 42672 23910 42674 23962
rect 42854 23910 42856 23962
rect 42610 23908 42616 23910
rect 42672 23908 42696 23910
rect 42752 23908 42776 23910
rect 42832 23908 42856 23910
rect 42912 23908 42918 23910
rect 42610 23899 42918 23908
rect 47610 23964 47918 23973
rect 47610 23962 47616 23964
rect 47672 23962 47696 23964
rect 47752 23962 47776 23964
rect 47832 23962 47856 23964
rect 47912 23962 47918 23964
rect 47672 23910 47674 23962
rect 47854 23910 47856 23962
rect 47610 23908 47616 23910
rect 47672 23908 47696 23910
rect 47752 23908 47776 23910
rect 47832 23908 47856 23910
rect 47912 23908 47918 23910
rect 47610 23899 47918 23908
rect 52610 23964 52918 23973
rect 52610 23962 52616 23964
rect 52672 23962 52696 23964
rect 52752 23962 52776 23964
rect 52832 23962 52856 23964
rect 52912 23962 52918 23964
rect 52672 23910 52674 23962
rect 52854 23910 52856 23962
rect 52610 23908 52616 23910
rect 52672 23908 52696 23910
rect 52752 23908 52776 23910
rect 52832 23908 52856 23910
rect 52912 23908 52918 23910
rect 52610 23899 52918 23908
rect 57610 23964 57918 23973
rect 57610 23962 57616 23964
rect 57672 23962 57696 23964
rect 57752 23962 57776 23964
rect 57832 23962 57856 23964
rect 57912 23962 57918 23964
rect 57672 23910 57674 23962
rect 57854 23910 57856 23962
rect 57610 23908 57616 23910
rect 57672 23908 57696 23910
rect 57752 23908 57776 23910
rect 57832 23908 57856 23910
rect 57912 23908 57918 23910
rect 57610 23899 57918 23908
rect 58544 23769 58572 24142
rect 58530 23760 58586 23769
rect 58530 23695 58586 23704
rect 1950 23420 2258 23429
rect 1950 23418 1956 23420
rect 2012 23418 2036 23420
rect 2092 23418 2116 23420
rect 2172 23418 2196 23420
rect 2252 23418 2258 23420
rect 2012 23366 2014 23418
rect 2194 23366 2196 23418
rect 1950 23364 1956 23366
rect 2012 23364 2036 23366
rect 2092 23364 2116 23366
rect 2172 23364 2196 23366
rect 2252 23364 2258 23366
rect 1950 23355 2258 23364
rect 6950 23420 7258 23429
rect 6950 23418 6956 23420
rect 7012 23418 7036 23420
rect 7092 23418 7116 23420
rect 7172 23418 7196 23420
rect 7252 23418 7258 23420
rect 7012 23366 7014 23418
rect 7194 23366 7196 23418
rect 6950 23364 6956 23366
rect 7012 23364 7036 23366
rect 7092 23364 7116 23366
rect 7172 23364 7196 23366
rect 7252 23364 7258 23366
rect 6950 23355 7258 23364
rect 11950 23420 12258 23429
rect 11950 23418 11956 23420
rect 12012 23418 12036 23420
rect 12092 23418 12116 23420
rect 12172 23418 12196 23420
rect 12252 23418 12258 23420
rect 12012 23366 12014 23418
rect 12194 23366 12196 23418
rect 11950 23364 11956 23366
rect 12012 23364 12036 23366
rect 12092 23364 12116 23366
rect 12172 23364 12196 23366
rect 12252 23364 12258 23366
rect 11950 23355 12258 23364
rect 16950 23420 17258 23429
rect 16950 23418 16956 23420
rect 17012 23418 17036 23420
rect 17092 23418 17116 23420
rect 17172 23418 17196 23420
rect 17252 23418 17258 23420
rect 17012 23366 17014 23418
rect 17194 23366 17196 23418
rect 16950 23364 16956 23366
rect 17012 23364 17036 23366
rect 17092 23364 17116 23366
rect 17172 23364 17196 23366
rect 17252 23364 17258 23366
rect 16950 23355 17258 23364
rect 21950 23420 22258 23429
rect 21950 23418 21956 23420
rect 22012 23418 22036 23420
rect 22092 23418 22116 23420
rect 22172 23418 22196 23420
rect 22252 23418 22258 23420
rect 22012 23366 22014 23418
rect 22194 23366 22196 23418
rect 21950 23364 21956 23366
rect 22012 23364 22036 23366
rect 22092 23364 22116 23366
rect 22172 23364 22196 23366
rect 22252 23364 22258 23366
rect 21950 23355 22258 23364
rect 26950 23420 27258 23429
rect 26950 23418 26956 23420
rect 27012 23418 27036 23420
rect 27092 23418 27116 23420
rect 27172 23418 27196 23420
rect 27252 23418 27258 23420
rect 27012 23366 27014 23418
rect 27194 23366 27196 23418
rect 26950 23364 26956 23366
rect 27012 23364 27036 23366
rect 27092 23364 27116 23366
rect 27172 23364 27196 23366
rect 27252 23364 27258 23366
rect 26950 23355 27258 23364
rect 31950 23420 32258 23429
rect 31950 23418 31956 23420
rect 32012 23418 32036 23420
rect 32092 23418 32116 23420
rect 32172 23418 32196 23420
rect 32252 23418 32258 23420
rect 32012 23366 32014 23418
rect 32194 23366 32196 23418
rect 31950 23364 31956 23366
rect 32012 23364 32036 23366
rect 32092 23364 32116 23366
rect 32172 23364 32196 23366
rect 32252 23364 32258 23366
rect 31950 23355 32258 23364
rect 36950 23420 37258 23429
rect 36950 23418 36956 23420
rect 37012 23418 37036 23420
rect 37092 23418 37116 23420
rect 37172 23418 37196 23420
rect 37252 23418 37258 23420
rect 37012 23366 37014 23418
rect 37194 23366 37196 23418
rect 36950 23364 36956 23366
rect 37012 23364 37036 23366
rect 37092 23364 37116 23366
rect 37172 23364 37196 23366
rect 37252 23364 37258 23366
rect 36950 23355 37258 23364
rect 41950 23420 42258 23429
rect 41950 23418 41956 23420
rect 42012 23418 42036 23420
rect 42092 23418 42116 23420
rect 42172 23418 42196 23420
rect 42252 23418 42258 23420
rect 42012 23366 42014 23418
rect 42194 23366 42196 23418
rect 41950 23364 41956 23366
rect 42012 23364 42036 23366
rect 42092 23364 42116 23366
rect 42172 23364 42196 23366
rect 42252 23364 42258 23366
rect 41950 23355 42258 23364
rect 46950 23420 47258 23429
rect 46950 23418 46956 23420
rect 47012 23418 47036 23420
rect 47092 23418 47116 23420
rect 47172 23418 47196 23420
rect 47252 23418 47258 23420
rect 47012 23366 47014 23418
rect 47194 23366 47196 23418
rect 46950 23364 46956 23366
rect 47012 23364 47036 23366
rect 47092 23364 47116 23366
rect 47172 23364 47196 23366
rect 47252 23364 47258 23366
rect 46950 23355 47258 23364
rect 51950 23420 52258 23429
rect 51950 23418 51956 23420
rect 52012 23418 52036 23420
rect 52092 23418 52116 23420
rect 52172 23418 52196 23420
rect 52252 23418 52258 23420
rect 52012 23366 52014 23418
rect 52194 23366 52196 23418
rect 51950 23364 51956 23366
rect 52012 23364 52036 23366
rect 52092 23364 52116 23366
rect 52172 23364 52196 23366
rect 52252 23364 52258 23366
rect 51950 23355 52258 23364
rect 56950 23420 57258 23429
rect 56950 23418 56956 23420
rect 57012 23418 57036 23420
rect 57092 23418 57116 23420
rect 57172 23418 57196 23420
rect 57252 23418 57258 23420
rect 57012 23366 57014 23418
rect 57194 23366 57196 23418
rect 56950 23364 56956 23366
rect 57012 23364 57036 23366
rect 57092 23364 57116 23366
rect 57172 23364 57196 23366
rect 57252 23364 57258 23366
rect 56950 23355 57258 23364
rect 58532 23112 58584 23118
rect 58532 23054 58584 23060
rect 58544 22953 58572 23054
rect 58530 22944 58586 22953
rect 2610 22876 2918 22885
rect 2610 22874 2616 22876
rect 2672 22874 2696 22876
rect 2752 22874 2776 22876
rect 2832 22874 2856 22876
rect 2912 22874 2918 22876
rect 2672 22822 2674 22874
rect 2854 22822 2856 22874
rect 2610 22820 2616 22822
rect 2672 22820 2696 22822
rect 2752 22820 2776 22822
rect 2832 22820 2856 22822
rect 2912 22820 2918 22822
rect 2610 22811 2918 22820
rect 7610 22876 7918 22885
rect 7610 22874 7616 22876
rect 7672 22874 7696 22876
rect 7752 22874 7776 22876
rect 7832 22874 7856 22876
rect 7912 22874 7918 22876
rect 7672 22822 7674 22874
rect 7854 22822 7856 22874
rect 7610 22820 7616 22822
rect 7672 22820 7696 22822
rect 7752 22820 7776 22822
rect 7832 22820 7856 22822
rect 7912 22820 7918 22822
rect 7610 22811 7918 22820
rect 12610 22876 12918 22885
rect 12610 22874 12616 22876
rect 12672 22874 12696 22876
rect 12752 22874 12776 22876
rect 12832 22874 12856 22876
rect 12912 22874 12918 22876
rect 12672 22822 12674 22874
rect 12854 22822 12856 22874
rect 12610 22820 12616 22822
rect 12672 22820 12696 22822
rect 12752 22820 12776 22822
rect 12832 22820 12856 22822
rect 12912 22820 12918 22822
rect 12610 22811 12918 22820
rect 17610 22876 17918 22885
rect 17610 22874 17616 22876
rect 17672 22874 17696 22876
rect 17752 22874 17776 22876
rect 17832 22874 17856 22876
rect 17912 22874 17918 22876
rect 17672 22822 17674 22874
rect 17854 22822 17856 22874
rect 17610 22820 17616 22822
rect 17672 22820 17696 22822
rect 17752 22820 17776 22822
rect 17832 22820 17856 22822
rect 17912 22820 17918 22822
rect 17610 22811 17918 22820
rect 22610 22876 22918 22885
rect 22610 22874 22616 22876
rect 22672 22874 22696 22876
rect 22752 22874 22776 22876
rect 22832 22874 22856 22876
rect 22912 22874 22918 22876
rect 22672 22822 22674 22874
rect 22854 22822 22856 22874
rect 22610 22820 22616 22822
rect 22672 22820 22696 22822
rect 22752 22820 22776 22822
rect 22832 22820 22856 22822
rect 22912 22820 22918 22822
rect 22610 22811 22918 22820
rect 27610 22876 27918 22885
rect 27610 22874 27616 22876
rect 27672 22874 27696 22876
rect 27752 22874 27776 22876
rect 27832 22874 27856 22876
rect 27912 22874 27918 22876
rect 27672 22822 27674 22874
rect 27854 22822 27856 22874
rect 27610 22820 27616 22822
rect 27672 22820 27696 22822
rect 27752 22820 27776 22822
rect 27832 22820 27856 22822
rect 27912 22820 27918 22822
rect 27610 22811 27918 22820
rect 32610 22876 32918 22885
rect 32610 22874 32616 22876
rect 32672 22874 32696 22876
rect 32752 22874 32776 22876
rect 32832 22874 32856 22876
rect 32912 22874 32918 22876
rect 32672 22822 32674 22874
rect 32854 22822 32856 22874
rect 32610 22820 32616 22822
rect 32672 22820 32696 22822
rect 32752 22820 32776 22822
rect 32832 22820 32856 22822
rect 32912 22820 32918 22822
rect 32610 22811 32918 22820
rect 37610 22876 37918 22885
rect 37610 22874 37616 22876
rect 37672 22874 37696 22876
rect 37752 22874 37776 22876
rect 37832 22874 37856 22876
rect 37912 22874 37918 22876
rect 37672 22822 37674 22874
rect 37854 22822 37856 22874
rect 37610 22820 37616 22822
rect 37672 22820 37696 22822
rect 37752 22820 37776 22822
rect 37832 22820 37856 22822
rect 37912 22820 37918 22822
rect 37610 22811 37918 22820
rect 42610 22876 42918 22885
rect 42610 22874 42616 22876
rect 42672 22874 42696 22876
rect 42752 22874 42776 22876
rect 42832 22874 42856 22876
rect 42912 22874 42918 22876
rect 42672 22822 42674 22874
rect 42854 22822 42856 22874
rect 42610 22820 42616 22822
rect 42672 22820 42696 22822
rect 42752 22820 42776 22822
rect 42832 22820 42856 22822
rect 42912 22820 42918 22822
rect 42610 22811 42918 22820
rect 47610 22876 47918 22885
rect 47610 22874 47616 22876
rect 47672 22874 47696 22876
rect 47752 22874 47776 22876
rect 47832 22874 47856 22876
rect 47912 22874 47918 22876
rect 47672 22822 47674 22874
rect 47854 22822 47856 22874
rect 47610 22820 47616 22822
rect 47672 22820 47696 22822
rect 47752 22820 47776 22822
rect 47832 22820 47856 22822
rect 47912 22820 47918 22822
rect 47610 22811 47918 22820
rect 52610 22876 52918 22885
rect 52610 22874 52616 22876
rect 52672 22874 52696 22876
rect 52752 22874 52776 22876
rect 52832 22874 52856 22876
rect 52912 22874 52918 22876
rect 52672 22822 52674 22874
rect 52854 22822 52856 22874
rect 52610 22820 52616 22822
rect 52672 22820 52696 22822
rect 52752 22820 52776 22822
rect 52832 22820 52856 22822
rect 52912 22820 52918 22822
rect 52610 22811 52918 22820
rect 57610 22876 57918 22885
rect 58530 22879 58586 22888
rect 57610 22874 57616 22876
rect 57672 22874 57696 22876
rect 57752 22874 57776 22876
rect 57832 22874 57856 22876
rect 57912 22874 57918 22876
rect 57672 22822 57674 22874
rect 57854 22822 57856 22874
rect 57610 22820 57616 22822
rect 57672 22820 57696 22822
rect 57752 22820 57776 22822
rect 57832 22820 57856 22822
rect 57912 22820 57918 22822
rect 57610 22811 57918 22820
rect 58532 22432 58584 22438
rect 58532 22374 58584 22380
rect 1950 22332 2258 22341
rect 1950 22330 1956 22332
rect 2012 22330 2036 22332
rect 2092 22330 2116 22332
rect 2172 22330 2196 22332
rect 2252 22330 2258 22332
rect 2012 22278 2014 22330
rect 2194 22278 2196 22330
rect 1950 22276 1956 22278
rect 2012 22276 2036 22278
rect 2092 22276 2116 22278
rect 2172 22276 2196 22278
rect 2252 22276 2258 22278
rect 1950 22267 2258 22276
rect 6950 22332 7258 22341
rect 6950 22330 6956 22332
rect 7012 22330 7036 22332
rect 7092 22330 7116 22332
rect 7172 22330 7196 22332
rect 7252 22330 7258 22332
rect 7012 22278 7014 22330
rect 7194 22278 7196 22330
rect 6950 22276 6956 22278
rect 7012 22276 7036 22278
rect 7092 22276 7116 22278
rect 7172 22276 7196 22278
rect 7252 22276 7258 22278
rect 6950 22267 7258 22276
rect 11950 22332 12258 22341
rect 11950 22330 11956 22332
rect 12012 22330 12036 22332
rect 12092 22330 12116 22332
rect 12172 22330 12196 22332
rect 12252 22330 12258 22332
rect 12012 22278 12014 22330
rect 12194 22278 12196 22330
rect 11950 22276 11956 22278
rect 12012 22276 12036 22278
rect 12092 22276 12116 22278
rect 12172 22276 12196 22278
rect 12252 22276 12258 22278
rect 11950 22267 12258 22276
rect 16950 22332 17258 22341
rect 16950 22330 16956 22332
rect 17012 22330 17036 22332
rect 17092 22330 17116 22332
rect 17172 22330 17196 22332
rect 17252 22330 17258 22332
rect 17012 22278 17014 22330
rect 17194 22278 17196 22330
rect 16950 22276 16956 22278
rect 17012 22276 17036 22278
rect 17092 22276 17116 22278
rect 17172 22276 17196 22278
rect 17252 22276 17258 22278
rect 16950 22267 17258 22276
rect 21950 22332 22258 22341
rect 21950 22330 21956 22332
rect 22012 22330 22036 22332
rect 22092 22330 22116 22332
rect 22172 22330 22196 22332
rect 22252 22330 22258 22332
rect 22012 22278 22014 22330
rect 22194 22278 22196 22330
rect 21950 22276 21956 22278
rect 22012 22276 22036 22278
rect 22092 22276 22116 22278
rect 22172 22276 22196 22278
rect 22252 22276 22258 22278
rect 21950 22267 22258 22276
rect 26950 22332 27258 22341
rect 26950 22330 26956 22332
rect 27012 22330 27036 22332
rect 27092 22330 27116 22332
rect 27172 22330 27196 22332
rect 27252 22330 27258 22332
rect 27012 22278 27014 22330
rect 27194 22278 27196 22330
rect 26950 22276 26956 22278
rect 27012 22276 27036 22278
rect 27092 22276 27116 22278
rect 27172 22276 27196 22278
rect 27252 22276 27258 22278
rect 26950 22267 27258 22276
rect 31950 22332 32258 22341
rect 31950 22330 31956 22332
rect 32012 22330 32036 22332
rect 32092 22330 32116 22332
rect 32172 22330 32196 22332
rect 32252 22330 32258 22332
rect 32012 22278 32014 22330
rect 32194 22278 32196 22330
rect 31950 22276 31956 22278
rect 32012 22276 32036 22278
rect 32092 22276 32116 22278
rect 32172 22276 32196 22278
rect 32252 22276 32258 22278
rect 31950 22267 32258 22276
rect 36950 22332 37258 22341
rect 36950 22330 36956 22332
rect 37012 22330 37036 22332
rect 37092 22330 37116 22332
rect 37172 22330 37196 22332
rect 37252 22330 37258 22332
rect 37012 22278 37014 22330
rect 37194 22278 37196 22330
rect 36950 22276 36956 22278
rect 37012 22276 37036 22278
rect 37092 22276 37116 22278
rect 37172 22276 37196 22278
rect 37252 22276 37258 22278
rect 36950 22267 37258 22276
rect 41950 22332 42258 22341
rect 41950 22330 41956 22332
rect 42012 22330 42036 22332
rect 42092 22330 42116 22332
rect 42172 22330 42196 22332
rect 42252 22330 42258 22332
rect 42012 22278 42014 22330
rect 42194 22278 42196 22330
rect 41950 22276 41956 22278
rect 42012 22276 42036 22278
rect 42092 22276 42116 22278
rect 42172 22276 42196 22278
rect 42252 22276 42258 22278
rect 41950 22267 42258 22276
rect 46950 22332 47258 22341
rect 46950 22330 46956 22332
rect 47012 22330 47036 22332
rect 47092 22330 47116 22332
rect 47172 22330 47196 22332
rect 47252 22330 47258 22332
rect 47012 22278 47014 22330
rect 47194 22278 47196 22330
rect 46950 22276 46956 22278
rect 47012 22276 47036 22278
rect 47092 22276 47116 22278
rect 47172 22276 47196 22278
rect 47252 22276 47258 22278
rect 46950 22267 47258 22276
rect 51950 22332 52258 22341
rect 51950 22330 51956 22332
rect 52012 22330 52036 22332
rect 52092 22330 52116 22332
rect 52172 22330 52196 22332
rect 52252 22330 52258 22332
rect 52012 22278 52014 22330
rect 52194 22278 52196 22330
rect 51950 22276 51956 22278
rect 52012 22276 52036 22278
rect 52092 22276 52116 22278
rect 52172 22276 52196 22278
rect 52252 22276 52258 22278
rect 51950 22267 52258 22276
rect 56950 22332 57258 22341
rect 56950 22330 56956 22332
rect 57012 22330 57036 22332
rect 57092 22330 57116 22332
rect 57172 22330 57196 22332
rect 57252 22330 57258 22332
rect 57012 22278 57014 22330
rect 57194 22278 57196 22330
rect 56950 22276 56956 22278
rect 57012 22276 57036 22278
rect 57092 22276 57116 22278
rect 57172 22276 57196 22278
rect 57252 22276 57258 22278
rect 56950 22267 57258 22276
rect 58544 22137 58572 22374
rect 58530 22128 58586 22137
rect 58530 22063 58586 22072
rect 2610 21788 2918 21797
rect 2610 21786 2616 21788
rect 2672 21786 2696 21788
rect 2752 21786 2776 21788
rect 2832 21786 2856 21788
rect 2912 21786 2918 21788
rect 2672 21734 2674 21786
rect 2854 21734 2856 21786
rect 2610 21732 2616 21734
rect 2672 21732 2696 21734
rect 2752 21732 2776 21734
rect 2832 21732 2856 21734
rect 2912 21732 2918 21734
rect 2610 21723 2918 21732
rect 7610 21788 7918 21797
rect 7610 21786 7616 21788
rect 7672 21786 7696 21788
rect 7752 21786 7776 21788
rect 7832 21786 7856 21788
rect 7912 21786 7918 21788
rect 7672 21734 7674 21786
rect 7854 21734 7856 21786
rect 7610 21732 7616 21734
rect 7672 21732 7696 21734
rect 7752 21732 7776 21734
rect 7832 21732 7856 21734
rect 7912 21732 7918 21734
rect 7610 21723 7918 21732
rect 12610 21788 12918 21797
rect 12610 21786 12616 21788
rect 12672 21786 12696 21788
rect 12752 21786 12776 21788
rect 12832 21786 12856 21788
rect 12912 21786 12918 21788
rect 12672 21734 12674 21786
rect 12854 21734 12856 21786
rect 12610 21732 12616 21734
rect 12672 21732 12696 21734
rect 12752 21732 12776 21734
rect 12832 21732 12856 21734
rect 12912 21732 12918 21734
rect 12610 21723 12918 21732
rect 17610 21788 17918 21797
rect 17610 21786 17616 21788
rect 17672 21786 17696 21788
rect 17752 21786 17776 21788
rect 17832 21786 17856 21788
rect 17912 21786 17918 21788
rect 17672 21734 17674 21786
rect 17854 21734 17856 21786
rect 17610 21732 17616 21734
rect 17672 21732 17696 21734
rect 17752 21732 17776 21734
rect 17832 21732 17856 21734
rect 17912 21732 17918 21734
rect 17610 21723 17918 21732
rect 22610 21788 22918 21797
rect 22610 21786 22616 21788
rect 22672 21786 22696 21788
rect 22752 21786 22776 21788
rect 22832 21786 22856 21788
rect 22912 21786 22918 21788
rect 22672 21734 22674 21786
rect 22854 21734 22856 21786
rect 22610 21732 22616 21734
rect 22672 21732 22696 21734
rect 22752 21732 22776 21734
rect 22832 21732 22856 21734
rect 22912 21732 22918 21734
rect 22610 21723 22918 21732
rect 27610 21788 27918 21797
rect 27610 21786 27616 21788
rect 27672 21786 27696 21788
rect 27752 21786 27776 21788
rect 27832 21786 27856 21788
rect 27912 21786 27918 21788
rect 27672 21734 27674 21786
rect 27854 21734 27856 21786
rect 27610 21732 27616 21734
rect 27672 21732 27696 21734
rect 27752 21732 27776 21734
rect 27832 21732 27856 21734
rect 27912 21732 27918 21734
rect 27610 21723 27918 21732
rect 32610 21788 32918 21797
rect 32610 21786 32616 21788
rect 32672 21786 32696 21788
rect 32752 21786 32776 21788
rect 32832 21786 32856 21788
rect 32912 21786 32918 21788
rect 32672 21734 32674 21786
rect 32854 21734 32856 21786
rect 32610 21732 32616 21734
rect 32672 21732 32696 21734
rect 32752 21732 32776 21734
rect 32832 21732 32856 21734
rect 32912 21732 32918 21734
rect 32610 21723 32918 21732
rect 37610 21788 37918 21797
rect 37610 21786 37616 21788
rect 37672 21786 37696 21788
rect 37752 21786 37776 21788
rect 37832 21786 37856 21788
rect 37912 21786 37918 21788
rect 37672 21734 37674 21786
rect 37854 21734 37856 21786
rect 37610 21732 37616 21734
rect 37672 21732 37696 21734
rect 37752 21732 37776 21734
rect 37832 21732 37856 21734
rect 37912 21732 37918 21734
rect 37610 21723 37918 21732
rect 42610 21788 42918 21797
rect 42610 21786 42616 21788
rect 42672 21786 42696 21788
rect 42752 21786 42776 21788
rect 42832 21786 42856 21788
rect 42912 21786 42918 21788
rect 42672 21734 42674 21786
rect 42854 21734 42856 21786
rect 42610 21732 42616 21734
rect 42672 21732 42696 21734
rect 42752 21732 42776 21734
rect 42832 21732 42856 21734
rect 42912 21732 42918 21734
rect 42610 21723 42918 21732
rect 47610 21788 47918 21797
rect 47610 21786 47616 21788
rect 47672 21786 47696 21788
rect 47752 21786 47776 21788
rect 47832 21786 47856 21788
rect 47912 21786 47918 21788
rect 47672 21734 47674 21786
rect 47854 21734 47856 21786
rect 47610 21732 47616 21734
rect 47672 21732 47696 21734
rect 47752 21732 47776 21734
rect 47832 21732 47856 21734
rect 47912 21732 47918 21734
rect 47610 21723 47918 21732
rect 52610 21788 52918 21797
rect 52610 21786 52616 21788
rect 52672 21786 52696 21788
rect 52752 21786 52776 21788
rect 52832 21786 52856 21788
rect 52912 21786 52918 21788
rect 52672 21734 52674 21786
rect 52854 21734 52856 21786
rect 52610 21732 52616 21734
rect 52672 21732 52696 21734
rect 52752 21732 52776 21734
rect 52832 21732 52856 21734
rect 52912 21732 52918 21734
rect 52610 21723 52918 21732
rect 57610 21788 57918 21797
rect 57610 21786 57616 21788
rect 57672 21786 57696 21788
rect 57752 21786 57776 21788
rect 57832 21786 57856 21788
rect 57912 21786 57918 21788
rect 57672 21734 57674 21786
rect 57854 21734 57856 21786
rect 57610 21732 57616 21734
rect 57672 21732 57696 21734
rect 57752 21732 57776 21734
rect 57832 21732 57856 21734
rect 57912 21732 57918 21734
rect 57610 21723 57918 21732
rect 58532 21344 58584 21350
rect 58530 21312 58532 21321
rect 58584 21312 58586 21321
rect 1950 21244 2258 21253
rect 1950 21242 1956 21244
rect 2012 21242 2036 21244
rect 2092 21242 2116 21244
rect 2172 21242 2196 21244
rect 2252 21242 2258 21244
rect 2012 21190 2014 21242
rect 2194 21190 2196 21242
rect 1950 21188 1956 21190
rect 2012 21188 2036 21190
rect 2092 21188 2116 21190
rect 2172 21188 2196 21190
rect 2252 21188 2258 21190
rect 1950 21179 2258 21188
rect 6950 21244 7258 21253
rect 6950 21242 6956 21244
rect 7012 21242 7036 21244
rect 7092 21242 7116 21244
rect 7172 21242 7196 21244
rect 7252 21242 7258 21244
rect 7012 21190 7014 21242
rect 7194 21190 7196 21242
rect 6950 21188 6956 21190
rect 7012 21188 7036 21190
rect 7092 21188 7116 21190
rect 7172 21188 7196 21190
rect 7252 21188 7258 21190
rect 6950 21179 7258 21188
rect 11950 21244 12258 21253
rect 11950 21242 11956 21244
rect 12012 21242 12036 21244
rect 12092 21242 12116 21244
rect 12172 21242 12196 21244
rect 12252 21242 12258 21244
rect 12012 21190 12014 21242
rect 12194 21190 12196 21242
rect 11950 21188 11956 21190
rect 12012 21188 12036 21190
rect 12092 21188 12116 21190
rect 12172 21188 12196 21190
rect 12252 21188 12258 21190
rect 11950 21179 12258 21188
rect 16950 21244 17258 21253
rect 16950 21242 16956 21244
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17252 21242 17258 21244
rect 17012 21190 17014 21242
rect 17194 21190 17196 21242
rect 16950 21188 16956 21190
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 17252 21188 17258 21190
rect 16950 21179 17258 21188
rect 21950 21244 22258 21253
rect 21950 21242 21956 21244
rect 22012 21242 22036 21244
rect 22092 21242 22116 21244
rect 22172 21242 22196 21244
rect 22252 21242 22258 21244
rect 22012 21190 22014 21242
rect 22194 21190 22196 21242
rect 21950 21188 21956 21190
rect 22012 21188 22036 21190
rect 22092 21188 22116 21190
rect 22172 21188 22196 21190
rect 22252 21188 22258 21190
rect 21950 21179 22258 21188
rect 26950 21244 27258 21253
rect 26950 21242 26956 21244
rect 27012 21242 27036 21244
rect 27092 21242 27116 21244
rect 27172 21242 27196 21244
rect 27252 21242 27258 21244
rect 27012 21190 27014 21242
rect 27194 21190 27196 21242
rect 26950 21188 26956 21190
rect 27012 21188 27036 21190
rect 27092 21188 27116 21190
rect 27172 21188 27196 21190
rect 27252 21188 27258 21190
rect 26950 21179 27258 21188
rect 31950 21244 32258 21253
rect 31950 21242 31956 21244
rect 32012 21242 32036 21244
rect 32092 21242 32116 21244
rect 32172 21242 32196 21244
rect 32252 21242 32258 21244
rect 32012 21190 32014 21242
rect 32194 21190 32196 21242
rect 31950 21188 31956 21190
rect 32012 21188 32036 21190
rect 32092 21188 32116 21190
rect 32172 21188 32196 21190
rect 32252 21188 32258 21190
rect 31950 21179 32258 21188
rect 36950 21244 37258 21253
rect 36950 21242 36956 21244
rect 37012 21242 37036 21244
rect 37092 21242 37116 21244
rect 37172 21242 37196 21244
rect 37252 21242 37258 21244
rect 37012 21190 37014 21242
rect 37194 21190 37196 21242
rect 36950 21188 36956 21190
rect 37012 21188 37036 21190
rect 37092 21188 37116 21190
rect 37172 21188 37196 21190
rect 37252 21188 37258 21190
rect 36950 21179 37258 21188
rect 41950 21244 42258 21253
rect 41950 21242 41956 21244
rect 42012 21242 42036 21244
rect 42092 21242 42116 21244
rect 42172 21242 42196 21244
rect 42252 21242 42258 21244
rect 42012 21190 42014 21242
rect 42194 21190 42196 21242
rect 41950 21188 41956 21190
rect 42012 21188 42036 21190
rect 42092 21188 42116 21190
rect 42172 21188 42196 21190
rect 42252 21188 42258 21190
rect 41950 21179 42258 21188
rect 46950 21244 47258 21253
rect 46950 21242 46956 21244
rect 47012 21242 47036 21244
rect 47092 21242 47116 21244
rect 47172 21242 47196 21244
rect 47252 21242 47258 21244
rect 47012 21190 47014 21242
rect 47194 21190 47196 21242
rect 46950 21188 46956 21190
rect 47012 21188 47036 21190
rect 47092 21188 47116 21190
rect 47172 21188 47196 21190
rect 47252 21188 47258 21190
rect 46950 21179 47258 21188
rect 51950 21244 52258 21253
rect 51950 21242 51956 21244
rect 52012 21242 52036 21244
rect 52092 21242 52116 21244
rect 52172 21242 52196 21244
rect 52252 21242 52258 21244
rect 52012 21190 52014 21242
rect 52194 21190 52196 21242
rect 51950 21188 51956 21190
rect 52012 21188 52036 21190
rect 52092 21188 52116 21190
rect 52172 21188 52196 21190
rect 52252 21188 52258 21190
rect 51950 21179 52258 21188
rect 56950 21244 57258 21253
rect 58530 21247 58586 21256
rect 56950 21242 56956 21244
rect 57012 21242 57036 21244
rect 57092 21242 57116 21244
rect 57172 21242 57196 21244
rect 57252 21242 57258 21244
rect 57012 21190 57014 21242
rect 57194 21190 57196 21242
rect 56950 21188 56956 21190
rect 57012 21188 57036 21190
rect 57092 21188 57116 21190
rect 57172 21188 57196 21190
rect 57252 21188 57258 21190
rect 56950 21179 57258 21188
rect 58532 20936 58584 20942
rect 58532 20878 58584 20884
rect 2610 20700 2918 20709
rect 2610 20698 2616 20700
rect 2672 20698 2696 20700
rect 2752 20698 2776 20700
rect 2832 20698 2856 20700
rect 2912 20698 2918 20700
rect 2672 20646 2674 20698
rect 2854 20646 2856 20698
rect 2610 20644 2616 20646
rect 2672 20644 2696 20646
rect 2752 20644 2776 20646
rect 2832 20644 2856 20646
rect 2912 20644 2918 20646
rect 2610 20635 2918 20644
rect 7610 20700 7918 20709
rect 7610 20698 7616 20700
rect 7672 20698 7696 20700
rect 7752 20698 7776 20700
rect 7832 20698 7856 20700
rect 7912 20698 7918 20700
rect 7672 20646 7674 20698
rect 7854 20646 7856 20698
rect 7610 20644 7616 20646
rect 7672 20644 7696 20646
rect 7752 20644 7776 20646
rect 7832 20644 7856 20646
rect 7912 20644 7918 20646
rect 7610 20635 7918 20644
rect 12610 20700 12918 20709
rect 12610 20698 12616 20700
rect 12672 20698 12696 20700
rect 12752 20698 12776 20700
rect 12832 20698 12856 20700
rect 12912 20698 12918 20700
rect 12672 20646 12674 20698
rect 12854 20646 12856 20698
rect 12610 20644 12616 20646
rect 12672 20644 12696 20646
rect 12752 20644 12776 20646
rect 12832 20644 12856 20646
rect 12912 20644 12918 20646
rect 12610 20635 12918 20644
rect 17610 20700 17918 20709
rect 17610 20698 17616 20700
rect 17672 20698 17696 20700
rect 17752 20698 17776 20700
rect 17832 20698 17856 20700
rect 17912 20698 17918 20700
rect 17672 20646 17674 20698
rect 17854 20646 17856 20698
rect 17610 20644 17616 20646
rect 17672 20644 17696 20646
rect 17752 20644 17776 20646
rect 17832 20644 17856 20646
rect 17912 20644 17918 20646
rect 17610 20635 17918 20644
rect 22610 20700 22918 20709
rect 22610 20698 22616 20700
rect 22672 20698 22696 20700
rect 22752 20698 22776 20700
rect 22832 20698 22856 20700
rect 22912 20698 22918 20700
rect 22672 20646 22674 20698
rect 22854 20646 22856 20698
rect 22610 20644 22616 20646
rect 22672 20644 22696 20646
rect 22752 20644 22776 20646
rect 22832 20644 22856 20646
rect 22912 20644 22918 20646
rect 22610 20635 22918 20644
rect 27610 20700 27918 20709
rect 27610 20698 27616 20700
rect 27672 20698 27696 20700
rect 27752 20698 27776 20700
rect 27832 20698 27856 20700
rect 27912 20698 27918 20700
rect 27672 20646 27674 20698
rect 27854 20646 27856 20698
rect 27610 20644 27616 20646
rect 27672 20644 27696 20646
rect 27752 20644 27776 20646
rect 27832 20644 27856 20646
rect 27912 20644 27918 20646
rect 27610 20635 27918 20644
rect 32610 20700 32918 20709
rect 32610 20698 32616 20700
rect 32672 20698 32696 20700
rect 32752 20698 32776 20700
rect 32832 20698 32856 20700
rect 32912 20698 32918 20700
rect 32672 20646 32674 20698
rect 32854 20646 32856 20698
rect 32610 20644 32616 20646
rect 32672 20644 32696 20646
rect 32752 20644 32776 20646
rect 32832 20644 32856 20646
rect 32912 20644 32918 20646
rect 32610 20635 32918 20644
rect 37610 20700 37918 20709
rect 37610 20698 37616 20700
rect 37672 20698 37696 20700
rect 37752 20698 37776 20700
rect 37832 20698 37856 20700
rect 37912 20698 37918 20700
rect 37672 20646 37674 20698
rect 37854 20646 37856 20698
rect 37610 20644 37616 20646
rect 37672 20644 37696 20646
rect 37752 20644 37776 20646
rect 37832 20644 37856 20646
rect 37912 20644 37918 20646
rect 37610 20635 37918 20644
rect 42610 20700 42918 20709
rect 42610 20698 42616 20700
rect 42672 20698 42696 20700
rect 42752 20698 42776 20700
rect 42832 20698 42856 20700
rect 42912 20698 42918 20700
rect 42672 20646 42674 20698
rect 42854 20646 42856 20698
rect 42610 20644 42616 20646
rect 42672 20644 42696 20646
rect 42752 20644 42776 20646
rect 42832 20644 42856 20646
rect 42912 20644 42918 20646
rect 42610 20635 42918 20644
rect 47610 20700 47918 20709
rect 47610 20698 47616 20700
rect 47672 20698 47696 20700
rect 47752 20698 47776 20700
rect 47832 20698 47856 20700
rect 47912 20698 47918 20700
rect 47672 20646 47674 20698
rect 47854 20646 47856 20698
rect 47610 20644 47616 20646
rect 47672 20644 47696 20646
rect 47752 20644 47776 20646
rect 47832 20644 47856 20646
rect 47912 20644 47918 20646
rect 47610 20635 47918 20644
rect 52610 20700 52918 20709
rect 52610 20698 52616 20700
rect 52672 20698 52696 20700
rect 52752 20698 52776 20700
rect 52832 20698 52856 20700
rect 52912 20698 52918 20700
rect 52672 20646 52674 20698
rect 52854 20646 52856 20698
rect 52610 20644 52616 20646
rect 52672 20644 52696 20646
rect 52752 20644 52776 20646
rect 52832 20644 52856 20646
rect 52912 20644 52918 20646
rect 52610 20635 52918 20644
rect 57610 20700 57918 20709
rect 57610 20698 57616 20700
rect 57672 20698 57696 20700
rect 57752 20698 57776 20700
rect 57832 20698 57856 20700
rect 57912 20698 57918 20700
rect 57672 20646 57674 20698
rect 57854 20646 57856 20698
rect 57610 20644 57616 20646
rect 57672 20644 57696 20646
rect 57752 20644 57776 20646
rect 57832 20644 57856 20646
rect 57912 20644 57918 20646
rect 57610 20635 57918 20644
rect 58544 20505 58572 20878
rect 58530 20496 58586 20505
rect 58530 20431 58586 20440
rect 1950 20156 2258 20165
rect 1950 20154 1956 20156
rect 2012 20154 2036 20156
rect 2092 20154 2116 20156
rect 2172 20154 2196 20156
rect 2252 20154 2258 20156
rect 2012 20102 2014 20154
rect 2194 20102 2196 20154
rect 1950 20100 1956 20102
rect 2012 20100 2036 20102
rect 2092 20100 2116 20102
rect 2172 20100 2196 20102
rect 2252 20100 2258 20102
rect 1950 20091 2258 20100
rect 6950 20156 7258 20165
rect 6950 20154 6956 20156
rect 7012 20154 7036 20156
rect 7092 20154 7116 20156
rect 7172 20154 7196 20156
rect 7252 20154 7258 20156
rect 7012 20102 7014 20154
rect 7194 20102 7196 20154
rect 6950 20100 6956 20102
rect 7012 20100 7036 20102
rect 7092 20100 7116 20102
rect 7172 20100 7196 20102
rect 7252 20100 7258 20102
rect 6950 20091 7258 20100
rect 11950 20156 12258 20165
rect 11950 20154 11956 20156
rect 12012 20154 12036 20156
rect 12092 20154 12116 20156
rect 12172 20154 12196 20156
rect 12252 20154 12258 20156
rect 12012 20102 12014 20154
rect 12194 20102 12196 20154
rect 11950 20100 11956 20102
rect 12012 20100 12036 20102
rect 12092 20100 12116 20102
rect 12172 20100 12196 20102
rect 12252 20100 12258 20102
rect 11950 20091 12258 20100
rect 16950 20156 17258 20165
rect 16950 20154 16956 20156
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17252 20154 17258 20156
rect 17012 20102 17014 20154
rect 17194 20102 17196 20154
rect 16950 20100 16956 20102
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 17252 20100 17258 20102
rect 16950 20091 17258 20100
rect 21950 20156 22258 20165
rect 21950 20154 21956 20156
rect 22012 20154 22036 20156
rect 22092 20154 22116 20156
rect 22172 20154 22196 20156
rect 22252 20154 22258 20156
rect 22012 20102 22014 20154
rect 22194 20102 22196 20154
rect 21950 20100 21956 20102
rect 22012 20100 22036 20102
rect 22092 20100 22116 20102
rect 22172 20100 22196 20102
rect 22252 20100 22258 20102
rect 21950 20091 22258 20100
rect 26950 20156 27258 20165
rect 26950 20154 26956 20156
rect 27012 20154 27036 20156
rect 27092 20154 27116 20156
rect 27172 20154 27196 20156
rect 27252 20154 27258 20156
rect 27012 20102 27014 20154
rect 27194 20102 27196 20154
rect 26950 20100 26956 20102
rect 27012 20100 27036 20102
rect 27092 20100 27116 20102
rect 27172 20100 27196 20102
rect 27252 20100 27258 20102
rect 26950 20091 27258 20100
rect 31950 20156 32258 20165
rect 31950 20154 31956 20156
rect 32012 20154 32036 20156
rect 32092 20154 32116 20156
rect 32172 20154 32196 20156
rect 32252 20154 32258 20156
rect 32012 20102 32014 20154
rect 32194 20102 32196 20154
rect 31950 20100 31956 20102
rect 32012 20100 32036 20102
rect 32092 20100 32116 20102
rect 32172 20100 32196 20102
rect 32252 20100 32258 20102
rect 31950 20091 32258 20100
rect 36950 20156 37258 20165
rect 36950 20154 36956 20156
rect 37012 20154 37036 20156
rect 37092 20154 37116 20156
rect 37172 20154 37196 20156
rect 37252 20154 37258 20156
rect 37012 20102 37014 20154
rect 37194 20102 37196 20154
rect 36950 20100 36956 20102
rect 37012 20100 37036 20102
rect 37092 20100 37116 20102
rect 37172 20100 37196 20102
rect 37252 20100 37258 20102
rect 36950 20091 37258 20100
rect 41950 20156 42258 20165
rect 41950 20154 41956 20156
rect 42012 20154 42036 20156
rect 42092 20154 42116 20156
rect 42172 20154 42196 20156
rect 42252 20154 42258 20156
rect 42012 20102 42014 20154
rect 42194 20102 42196 20154
rect 41950 20100 41956 20102
rect 42012 20100 42036 20102
rect 42092 20100 42116 20102
rect 42172 20100 42196 20102
rect 42252 20100 42258 20102
rect 41950 20091 42258 20100
rect 46950 20156 47258 20165
rect 46950 20154 46956 20156
rect 47012 20154 47036 20156
rect 47092 20154 47116 20156
rect 47172 20154 47196 20156
rect 47252 20154 47258 20156
rect 47012 20102 47014 20154
rect 47194 20102 47196 20154
rect 46950 20100 46956 20102
rect 47012 20100 47036 20102
rect 47092 20100 47116 20102
rect 47172 20100 47196 20102
rect 47252 20100 47258 20102
rect 46950 20091 47258 20100
rect 51950 20156 52258 20165
rect 51950 20154 51956 20156
rect 52012 20154 52036 20156
rect 52092 20154 52116 20156
rect 52172 20154 52196 20156
rect 52252 20154 52258 20156
rect 52012 20102 52014 20154
rect 52194 20102 52196 20154
rect 51950 20100 51956 20102
rect 52012 20100 52036 20102
rect 52092 20100 52116 20102
rect 52172 20100 52196 20102
rect 52252 20100 52258 20102
rect 51950 20091 52258 20100
rect 56950 20156 57258 20165
rect 56950 20154 56956 20156
rect 57012 20154 57036 20156
rect 57092 20154 57116 20156
rect 57172 20154 57196 20156
rect 57252 20154 57258 20156
rect 57012 20102 57014 20154
rect 57194 20102 57196 20154
rect 56950 20100 56956 20102
rect 57012 20100 57036 20102
rect 57092 20100 57116 20102
rect 57172 20100 57196 20102
rect 57252 20100 57258 20102
rect 56950 20091 57258 20100
rect 58532 19848 58584 19854
rect 58532 19790 58584 19796
rect 58544 19689 58572 19790
rect 58530 19680 58586 19689
rect 2610 19612 2918 19621
rect 2610 19610 2616 19612
rect 2672 19610 2696 19612
rect 2752 19610 2776 19612
rect 2832 19610 2856 19612
rect 2912 19610 2918 19612
rect 2672 19558 2674 19610
rect 2854 19558 2856 19610
rect 2610 19556 2616 19558
rect 2672 19556 2696 19558
rect 2752 19556 2776 19558
rect 2832 19556 2856 19558
rect 2912 19556 2918 19558
rect 2610 19547 2918 19556
rect 7610 19612 7918 19621
rect 7610 19610 7616 19612
rect 7672 19610 7696 19612
rect 7752 19610 7776 19612
rect 7832 19610 7856 19612
rect 7912 19610 7918 19612
rect 7672 19558 7674 19610
rect 7854 19558 7856 19610
rect 7610 19556 7616 19558
rect 7672 19556 7696 19558
rect 7752 19556 7776 19558
rect 7832 19556 7856 19558
rect 7912 19556 7918 19558
rect 7610 19547 7918 19556
rect 12610 19612 12918 19621
rect 12610 19610 12616 19612
rect 12672 19610 12696 19612
rect 12752 19610 12776 19612
rect 12832 19610 12856 19612
rect 12912 19610 12918 19612
rect 12672 19558 12674 19610
rect 12854 19558 12856 19610
rect 12610 19556 12616 19558
rect 12672 19556 12696 19558
rect 12752 19556 12776 19558
rect 12832 19556 12856 19558
rect 12912 19556 12918 19558
rect 12610 19547 12918 19556
rect 17610 19612 17918 19621
rect 17610 19610 17616 19612
rect 17672 19610 17696 19612
rect 17752 19610 17776 19612
rect 17832 19610 17856 19612
rect 17912 19610 17918 19612
rect 17672 19558 17674 19610
rect 17854 19558 17856 19610
rect 17610 19556 17616 19558
rect 17672 19556 17696 19558
rect 17752 19556 17776 19558
rect 17832 19556 17856 19558
rect 17912 19556 17918 19558
rect 17610 19547 17918 19556
rect 22610 19612 22918 19621
rect 22610 19610 22616 19612
rect 22672 19610 22696 19612
rect 22752 19610 22776 19612
rect 22832 19610 22856 19612
rect 22912 19610 22918 19612
rect 22672 19558 22674 19610
rect 22854 19558 22856 19610
rect 22610 19556 22616 19558
rect 22672 19556 22696 19558
rect 22752 19556 22776 19558
rect 22832 19556 22856 19558
rect 22912 19556 22918 19558
rect 22610 19547 22918 19556
rect 27610 19612 27918 19621
rect 27610 19610 27616 19612
rect 27672 19610 27696 19612
rect 27752 19610 27776 19612
rect 27832 19610 27856 19612
rect 27912 19610 27918 19612
rect 27672 19558 27674 19610
rect 27854 19558 27856 19610
rect 27610 19556 27616 19558
rect 27672 19556 27696 19558
rect 27752 19556 27776 19558
rect 27832 19556 27856 19558
rect 27912 19556 27918 19558
rect 27610 19547 27918 19556
rect 32610 19612 32918 19621
rect 32610 19610 32616 19612
rect 32672 19610 32696 19612
rect 32752 19610 32776 19612
rect 32832 19610 32856 19612
rect 32912 19610 32918 19612
rect 32672 19558 32674 19610
rect 32854 19558 32856 19610
rect 32610 19556 32616 19558
rect 32672 19556 32696 19558
rect 32752 19556 32776 19558
rect 32832 19556 32856 19558
rect 32912 19556 32918 19558
rect 32610 19547 32918 19556
rect 37610 19612 37918 19621
rect 37610 19610 37616 19612
rect 37672 19610 37696 19612
rect 37752 19610 37776 19612
rect 37832 19610 37856 19612
rect 37912 19610 37918 19612
rect 37672 19558 37674 19610
rect 37854 19558 37856 19610
rect 37610 19556 37616 19558
rect 37672 19556 37696 19558
rect 37752 19556 37776 19558
rect 37832 19556 37856 19558
rect 37912 19556 37918 19558
rect 37610 19547 37918 19556
rect 42610 19612 42918 19621
rect 42610 19610 42616 19612
rect 42672 19610 42696 19612
rect 42752 19610 42776 19612
rect 42832 19610 42856 19612
rect 42912 19610 42918 19612
rect 42672 19558 42674 19610
rect 42854 19558 42856 19610
rect 42610 19556 42616 19558
rect 42672 19556 42696 19558
rect 42752 19556 42776 19558
rect 42832 19556 42856 19558
rect 42912 19556 42918 19558
rect 42610 19547 42918 19556
rect 47610 19612 47918 19621
rect 47610 19610 47616 19612
rect 47672 19610 47696 19612
rect 47752 19610 47776 19612
rect 47832 19610 47856 19612
rect 47912 19610 47918 19612
rect 47672 19558 47674 19610
rect 47854 19558 47856 19610
rect 47610 19556 47616 19558
rect 47672 19556 47696 19558
rect 47752 19556 47776 19558
rect 47832 19556 47856 19558
rect 47912 19556 47918 19558
rect 47610 19547 47918 19556
rect 52610 19612 52918 19621
rect 52610 19610 52616 19612
rect 52672 19610 52696 19612
rect 52752 19610 52776 19612
rect 52832 19610 52856 19612
rect 52912 19610 52918 19612
rect 52672 19558 52674 19610
rect 52854 19558 52856 19610
rect 52610 19556 52616 19558
rect 52672 19556 52696 19558
rect 52752 19556 52776 19558
rect 52832 19556 52856 19558
rect 52912 19556 52918 19558
rect 52610 19547 52918 19556
rect 57610 19612 57918 19621
rect 58530 19615 58586 19624
rect 57610 19610 57616 19612
rect 57672 19610 57696 19612
rect 57752 19610 57776 19612
rect 57832 19610 57856 19612
rect 57912 19610 57918 19612
rect 57672 19558 57674 19610
rect 57854 19558 57856 19610
rect 57610 19556 57616 19558
rect 57672 19556 57696 19558
rect 57752 19556 57776 19558
rect 57832 19556 57856 19558
rect 57912 19556 57918 19558
rect 57610 19547 57918 19556
rect 58532 19168 58584 19174
rect 58532 19110 58584 19116
rect 1950 19068 2258 19077
rect 1950 19066 1956 19068
rect 2012 19066 2036 19068
rect 2092 19066 2116 19068
rect 2172 19066 2196 19068
rect 2252 19066 2258 19068
rect 2012 19014 2014 19066
rect 2194 19014 2196 19066
rect 1950 19012 1956 19014
rect 2012 19012 2036 19014
rect 2092 19012 2116 19014
rect 2172 19012 2196 19014
rect 2252 19012 2258 19014
rect 1950 19003 2258 19012
rect 6950 19068 7258 19077
rect 6950 19066 6956 19068
rect 7012 19066 7036 19068
rect 7092 19066 7116 19068
rect 7172 19066 7196 19068
rect 7252 19066 7258 19068
rect 7012 19014 7014 19066
rect 7194 19014 7196 19066
rect 6950 19012 6956 19014
rect 7012 19012 7036 19014
rect 7092 19012 7116 19014
rect 7172 19012 7196 19014
rect 7252 19012 7258 19014
rect 6950 19003 7258 19012
rect 11950 19068 12258 19077
rect 11950 19066 11956 19068
rect 12012 19066 12036 19068
rect 12092 19066 12116 19068
rect 12172 19066 12196 19068
rect 12252 19066 12258 19068
rect 12012 19014 12014 19066
rect 12194 19014 12196 19066
rect 11950 19012 11956 19014
rect 12012 19012 12036 19014
rect 12092 19012 12116 19014
rect 12172 19012 12196 19014
rect 12252 19012 12258 19014
rect 11950 19003 12258 19012
rect 16950 19068 17258 19077
rect 16950 19066 16956 19068
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17252 19066 17258 19068
rect 17012 19014 17014 19066
rect 17194 19014 17196 19066
rect 16950 19012 16956 19014
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 17252 19012 17258 19014
rect 16950 19003 17258 19012
rect 21950 19068 22258 19077
rect 21950 19066 21956 19068
rect 22012 19066 22036 19068
rect 22092 19066 22116 19068
rect 22172 19066 22196 19068
rect 22252 19066 22258 19068
rect 22012 19014 22014 19066
rect 22194 19014 22196 19066
rect 21950 19012 21956 19014
rect 22012 19012 22036 19014
rect 22092 19012 22116 19014
rect 22172 19012 22196 19014
rect 22252 19012 22258 19014
rect 21950 19003 22258 19012
rect 26950 19068 27258 19077
rect 26950 19066 26956 19068
rect 27012 19066 27036 19068
rect 27092 19066 27116 19068
rect 27172 19066 27196 19068
rect 27252 19066 27258 19068
rect 27012 19014 27014 19066
rect 27194 19014 27196 19066
rect 26950 19012 26956 19014
rect 27012 19012 27036 19014
rect 27092 19012 27116 19014
rect 27172 19012 27196 19014
rect 27252 19012 27258 19014
rect 26950 19003 27258 19012
rect 31950 19068 32258 19077
rect 31950 19066 31956 19068
rect 32012 19066 32036 19068
rect 32092 19066 32116 19068
rect 32172 19066 32196 19068
rect 32252 19066 32258 19068
rect 32012 19014 32014 19066
rect 32194 19014 32196 19066
rect 31950 19012 31956 19014
rect 32012 19012 32036 19014
rect 32092 19012 32116 19014
rect 32172 19012 32196 19014
rect 32252 19012 32258 19014
rect 31950 19003 32258 19012
rect 36950 19068 37258 19077
rect 36950 19066 36956 19068
rect 37012 19066 37036 19068
rect 37092 19066 37116 19068
rect 37172 19066 37196 19068
rect 37252 19066 37258 19068
rect 37012 19014 37014 19066
rect 37194 19014 37196 19066
rect 36950 19012 36956 19014
rect 37012 19012 37036 19014
rect 37092 19012 37116 19014
rect 37172 19012 37196 19014
rect 37252 19012 37258 19014
rect 36950 19003 37258 19012
rect 41950 19068 42258 19077
rect 41950 19066 41956 19068
rect 42012 19066 42036 19068
rect 42092 19066 42116 19068
rect 42172 19066 42196 19068
rect 42252 19066 42258 19068
rect 42012 19014 42014 19066
rect 42194 19014 42196 19066
rect 41950 19012 41956 19014
rect 42012 19012 42036 19014
rect 42092 19012 42116 19014
rect 42172 19012 42196 19014
rect 42252 19012 42258 19014
rect 41950 19003 42258 19012
rect 46950 19068 47258 19077
rect 46950 19066 46956 19068
rect 47012 19066 47036 19068
rect 47092 19066 47116 19068
rect 47172 19066 47196 19068
rect 47252 19066 47258 19068
rect 47012 19014 47014 19066
rect 47194 19014 47196 19066
rect 46950 19012 46956 19014
rect 47012 19012 47036 19014
rect 47092 19012 47116 19014
rect 47172 19012 47196 19014
rect 47252 19012 47258 19014
rect 46950 19003 47258 19012
rect 51950 19068 52258 19077
rect 51950 19066 51956 19068
rect 52012 19066 52036 19068
rect 52092 19066 52116 19068
rect 52172 19066 52196 19068
rect 52252 19066 52258 19068
rect 52012 19014 52014 19066
rect 52194 19014 52196 19066
rect 51950 19012 51956 19014
rect 52012 19012 52036 19014
rect 52092 19012 52116 19014
rect 52172 19012 52196 19014
rect 52252 19012 52258 19014
rect 51950 19003 52258 19012
rect 56950 19068 57258 19077
rect 56950 19066 56956 19068
rect 57012 19066 57036 19068
rect 57092 19066 57116 19068
rect 57172 19066 57196 19068
rect 57252 19066 57258 19068
rect 57012 19014 57014 19066
rect 57194 19014 57196 19066
rect 56950 19012 56956 19014
rect 57012 19012 57036 19014
rect 57092 19012 57116 19014
rect 57172 19012 57196 19014
rect 57252 19012 57258 19014
rect 56950 19003 57258 19012
rect 58544 18873 58572 19110
rect 58530 18864 58586 18873
rect 58530 18799 58586 18808
rect 2610 18524 2918 18533
rect 2610 18522 2616 18524
rect 2672 18522 2696 18524
rect 2752 18522 2776 18524
rect 2832 18522 2856 18524
rect 2912 18522 2918 18524
rect 2672 18470 2674 18522
rect 2854 18470 2856 18522
rect 2610 18468 2616 18470
rect 2672 18468 2696 18470
rect 2752 18468 2776 18470
rect 2832 18468 2856 18470
rect 2912 18468 2918 18470
rect 2610 18459 2918 18468
rect 7610 18524 7918 18533
rect 7610 18522 7616 18524
rect 7672 18522 7696 18524
rect 7752 18522 7776 18524
rect 7832 18522 7856 18524
rect 7912 18522 7918 18524
rect 7672 18470 7674 18522
rect 7854 18470 7856 18522
rect 7610 18468 7616 18470
rect 7672 18468 7696 18470
rect 7752 18468 7776 18470
rect 7832 18468 7856 18470
rect 7912 18468 7918 18470
rect 7610 18459 7918 18468
rect 12610 18524 12918 18533
rect 12610 18522 12616 18524
rect 12672 18522 12696 18524
rect 12752 18522 12776 18524
rect 12832 18522 12856 18524
rect 12912 18522 12918 18524
rect 12672 18470 12674 18522
rect 12854 18470 12856 18522
rect 12610 18468 12616 18470
rect 12672 18468 12696 18470
rect 12752 18468 12776 18470
rect 12832 18468 12856 18470
rect 12912 18468 12918 18470
rect 12610 18459 12918 18468
rect 17610 18524 17918 18533
rect 17610 18522 17616 18524
rect 17672 18522 17696 18524
rect 17752 18522 17776 18524
rect 17832 18522 17856 18524
rect 17912 18522 17918 18524
rect 17672 18470 17674 18522
rect 17854 18470 17856 18522
rect 17610 18468 17616 18470
rect 17672 18468 17696 18470
rect 17752 18468 17776 18470
rect 17832 18468 17856 18470
rect 17912 18468 17918 18470
rect 17610 18459 17918 18468
rect 22610 18524 22918 18533
rect 22610 18522 22616 18524
rect 22672 18522 22696 18524
rect 22752 18522 22776 18524
rect 22832 18522 22856 18524
rect 22912 18522 22918 18524
rect 22672 18470 22674 18522
rect 22854 18470 22856 18522
rect 22610 18468 22616 18470
rect 22672 18468 22696 18470
rect 22752 18468 22776 18470
rect 22832 18468 22856 18470
rect 22912 18468 22918 18470
rect 22610 18459 22918 18468
rect 27610 18524 27918 18533
rect 27610 18522 27616 18524
rect 27672 18522 27696 18524
rect 27752 18522 27776 18524
rect 27832 18522 27856 18524
rect 27912 18522 27918 18524
rect 27672 18470 27674 18522
rect 27854 18470 27856 18522
rect 27610 18468 27616 18470
rect 27672 18468 27696 18470
rect 27752 18468 27776 18470
rect 27832 18468 27856 18470
rect 27912 18468 27918 18470
rect 27610 18459 27918 18468
rect 32610 18524 32918 18533
rect 32610 18522 32616 18524
rect 32672 18522 32696 18524
rect 32752 18522 32776 18524
rect 32832 18522 32856 18524
rect 32912 18522 32918 18524
rect 32672 18470 32674 18522
rect 32854 18470 32856 18522
rect 32610 18468 32616 18470
rect 32672 18468 32696 18470
rect 32752 18468 32776 18470
rect 32832 18468 32856 18470
rect 32912 18468 32918 18470
rect 32610 18459 32918 18468
rect 37610 18524 37918 18533
rect 37610 18522 37616 18524
rect 37672 18522 37696 18524
rect 37752 18522 37776 18524
rect 37832 18522 37856 18524
rect 37912 18522 37918 18524
rect 37672 18470 37674 18522
rect 37854 18470 37856 18522
rect 37610 18468 37616 18470
rect 37672 18468 37696 18470
rect 37752 18468 37776 18470
rect 37832 18468 37856 18470
rect 37912 18468 37918 18470
rect 37610 18459 37918 18468
rect 42610 18524 42918 18533
rect 42610 18522 42616 18524
rect 42672 18522 42696 18524
rect 42752 18522 42776 18524
rect 42832 18522 42856 18524
rect 42912 18522 42918 18524
rect 42672 18470 42674 18522
rect 42854 18470 42856 18522
rect 42610 18468 42616 18470
rect 42672 18468 42696 18470
rect 42752 18468 42776 18470
rect 42832 18468 42856 18470
rect 42912 18468 42918 18470
rect 42610 18459 42918 18468
rect 47610 18524 47918 18533
rect 47610 18522 47616 18524
rect 47672 18522 47696 18524
rect 47752 18522 47776 18524
rect 47832 18522 47856 18524
rect 47912 18522 47918 18524
rect 47672 18470 47674 18522
rect 47854 18470 47856 18522
rect 47610 18468 47616 18470
rect 47672 18468 47696 18470
rect 47752 18468 47776 18470
rect 47832 18468 47856 18470
rect 47912 18468 47918 18470
rect 47610 18459 47918 18468
rect 52610 18524 52918 18533
rect 52610 18522 52616 18524
rect 52672 18522 52696 18524
rect 52752 18522 52776 18524
rect 52832 18522 52856 18524
rect 52912 18522 52918 18524
rect 52672 18470 52674 18522
rect 52854 18470 52856 18522
rect 52610 18468 52616 18470
rect 52672 18468 52696 18470
rect 52752 18468 52776 18470
rect 52832 18468 52856 18470
rect 52912 18468 52918 18470
rect 52610 18459 52918 18468
rect 57610 18524 57918 18533
rect 57610 18522 57616 18524
rect 57672 18522 57696 18524
rect 57752 18522 57776 18524
rect 57832 18522 57856 18524
rect 57912 18522 57918 18524
rect 57672 18470 57674 18522
rect 57854 18470 57856 18522
rect 57610 18468 57616 18470
rect 57672 18468 57696 18470
rect 57752 18468 57776 18470
rect 57832 18468 57856 18470
rect 57912 18468 57918 18470
rect 57610 18459 57918 18468
rect 58532 18080 58584 18086
rect 58530 18048 58532 18057
rect 58584 18048 58586 18057
rect 1950 17980 2258 17989
rect 1950 17978 1956 17980
rect 2012 17978 2036 17980
rect 2092 17978 2116 17980
rect 2172 17978 2196 17980
rect 2252 17978 2258 17980
rect 2012 17926 2014 17978
rect 2194 17926 2196 17978
rect 1950 17924 1956 17926
rect 2012 17924 2036 17926
rect 2092 17924 2116 17926
rect 2172 17924 2196 17926
rect 2252 17924 2258 17926
rect 1950 17915 2258 17924
rect 6950 17980 7258 17989
rect 6950 17978 6956 17980
rect 7012 17978 7036 17980
rect 7092 17978 7116 17980
rect 7172 17978 7196 17980
rect 7252 17978 7258 17980
rect 7012 17926 7014 17978
rect 7194 17926 7196 17978
rect 6950 17924 6956 17926
rect 7012 17924 7036 17926
rect 7092 17924 7116 17926
rect 7172 17924 7196 17926
rect 7252 17924 7258 17926
rect 6950 17915 7258 17924
rect 11950 17980 12258 17989
rect 11950 17978 11956 17980
rect 12012 17978 12036 17980
rect 12092 17978 12116 17980
rect 12172 17978 12196 17980
rect 12252 17978 12258 17980
rect 12012 17926 12014 17978
rect 12194 17926 12196 17978
rect 11950 17924 11956 17926
rect 12012 17924 12036 17926
rect 12092 17924 12116 17926
rect 12172 17924 12196 17926
rect 12252 17924 12258 17926
rect 11950 17915 12258 17924
rect 16950 17980 17258 17989
rect 16950 17978 16956 17980
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17252 17978 17258 17980
rect 17012 17926 17014 17978
rect 17194 17926 17196 17978
rect 16950 17924 16956 17926
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 17252 17924 17258 17926
rect 16950 17915 17258 17924
rect 21950 17980 22258 17989
rect 21950 17978 21956 17980
rect 22012 17978 22036 17980
rect 22092 17978 22116 17980
rect 22172 17978 22196 17980
rect 22252 17978 22258 17980
rect 22012 17926 22014 17978
rect 22194 17926 22196 17978
rect 21950 17924 21956 17926
rect 22012 17924 22036 17926
rect 22092 17924 22116 17926
rect 22172 17924 22196 17926
rect 22252 17924 22258 17926
rect 21950 17915 22258 17924
rect 26950 17980 27258 17989
rect 26950 17978 26956 17980
rect 27012 17978 27036 17980
rect 27092 17978 27116 17980
rect 27172 17978 27196 17980
rect 27252 17978 27258 17980
rect 27012 17926 27014 17978
rect 27194 17926 27196 17978
rect 26950 17924 26956 17926
rect 27012 17924 27036 17926
rect 27092 17924 27116 17926
rect 27172 17924 27196 17926
rect 27252 17924 27258 17926
rect 26950 17915 27258 17924
rect 31950 17980 32258 17989
rect 31950 17978 31956 17980
rect 32012 17978 32036 17980
rect 32092 17978 32116 17980
rect 32172 17978 32196 17980
rect 32252 17978 32258 17980
rect 32012 17926 32014 17978
rect 32194 17926 32196 17978
rect 31950 17924 31956 17926
rect 32012 17924 32036 17926
rect 32092 17924 32116 17926
rect 32172 17924 32196 17926
rect 32252 17924 32258 17926
rect 31950 17915 32258 17924
rect 36950 17980 37258 17989
rect 36950 17978 36956 17980
rect 37012 17978 37036 17980
rect 37092 17978 37116 17980
rect 37172 17978 37196 17980
rect 37252 17978 37258 17980
rect 37012 17926 37014 17978
rect 37194 17926 37196 17978
rect 36950 17924 36956 17926
rect 37012 17924 37036 17926
rect 37092 17924 37116 17926
rect 37172 17924 37196 17926
rect 37252 17924 37258 17926
rect 36950 17915 37258 17924
rect 41950 17980 42258 17989
rect 41950 17978 41956 17980
rect 42012 17978 42036 17980
rect 42092 17978 42116 17980
rect 42172 17978 42196 17980
rect 42252 17978 42258 17980
rect 42012 17926 42014 17978
rect 42194 17926 42196 17978
rect 41950 17924 41956 17926
rect 42012 17924 42036 17926
rect 42092 17924 42116 17926
rect 42172 17924 42196 17926
rect 42252 17924 42258 17926
rect 41950 17915 42258 17924
rect 46950 17980 47258 17989
rect 46950 17978 46956 17980
rect 47012 17978 47036 17980
rect 47092 17978 47116 17980
rect 47172 17978 47196 17980
rect 47252 17978 47258 17980
rect 47012 17926 47014 17978
rect 47194 17926 47196 17978
rect 46950 17924 46956 17926
rect 47012 17924 47036 17926
rect 47092 17924 47116 17926
rect 47172 17924 47196 17926
rect 47252 17924 47258 17926
rect 46950 17915 47258 17924
rect 51950 17980 52258 17989
rect 51950 17978 51956 17980
rect 52012 17978 52036 17980
rect 52092 17978 52116 17980
rect 52172 17978 52196 17980
rect 52252 17978 52258 17980
rect 52012 17926 52014 17978
rect 52194 17926 52196 17978
rect 51950 17924 51956 17926
rect 52012 17924 52036 17926
rect 52092 17924 52116 17926
rect 52172 17924 52196 17926
rect 52252 17924 52258 17926
rect 51950 17915 52258 17924
rect 56950 17980 57258 17989
rect 58530 17983 58586 17992
rect 56950 17978 56956 17980
rect 57012 17978 57036 17980
rect 57092 17978 57116 17980
rect 57172 17978 57196 17980
rect 57252 17978 57258 17980
rect 57012 17926 57014 17978
rect 57194 17926 57196 17978
rect 56950 17924 56956 17926
rect 57012 17924 57036 17926
rect 57092 17924 57116 17926
rect 57172 17924 57196 17926
rect 57252 17924 57258 17926
rect 56950 17915 57258 17924
rect 58532 17672 58584 17678
rect 58532 17614 58584 17620
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7610 17371 7918 17380
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 17610 17436 17918 17445
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 22610 17436 22918 17445
rect 22610 17434 22616 17436
rect 22672 17434 22696 17436
rect 22752 17434 22776 17436
rect 22832 17434 22856 17436
rect 22912 17434 22918 17436
rect 22672 17382 22674 17434
rect 22854 17382 22856 17434
rect 22610 17380 22616 17382
rect 22672 17380 22696 17382
rect 22752 17380 22776 17382
rect 22832 17380 22856 17382
rect 22912 17380 22918 17382
rect 22610 17371 22918 17380
rect 27610 17436 27918 17445
rect 27610 17434 27616 17436
rect 27672 17434 27696 17436
rect 27752 17434 27776 17436
rect 27832 17434 27856 17436
rect 27912 17434 27918 17436
rect 27672 17382 27674 17434
rect 27854 17382 27856 17434
rect 27610 17380 27616 17382
rect 27672 17380 27696 17382
rect 27752 17380 27776 17382
rect 27832 17380 27856 17382
rect 27912 17380 27918 17382
rect 27610 17371 27918 17380
rect 32610 17436 32918 17445
rect 32610 17434 32616 17436
rect 32672 17434 32696 17436
rect 32752 17434 32776 17436
rect 32832 17434 32856 17436
rect 32912 17434 32918 17436
rect 32672 17382 32674 17434
rect 32854 17382 32856 17434
rect 32610 17380 32616 17382
rect 32672 17380 32696 17382
rect 32752 17380 32776 17382
rect 32832 17380 32856 17382
rect 32912 17380 32918 17382
rect 32610 17371 32918 17380
rect 37610 17436 37918 17445
rect 37610 17434 37616 17436
rect 37672 17434 37696 17436
rect 37752 17434 37776 17436
rect 37832 17434 37856 17436
rect 37912 17434 37918 17436
rect 37672 17382 37674 17434
rect 37854 17382 37856 17434
rect 37610 17380 37616 17382
rect 37672 17380 37696 17382
rect 37752 17380 37776 17382
rect 37832 17380 37856 17382
rect 37912 17380 37918 17382
rect 37610 17371 37918 17380
rect 42610 17436 42918 17445
rect 42610 17434 42616 17436
rect 42672 17434 42696 17436
rect 42752 17434 42776 17436
rect 42832 17434 42856 17436
rect 42912 17434 42918 17436
rect 42672 17382 42674 17434
rect 42854 17382 42856 17434
rect 42610 17380 42616 17382
rect 42672 17380 42696 17382
rect 42752 17380 42776 17382
rect 42832 17380 42856 17382
rect 42912 17380 42918 17382
rect 42610 17371 42918 17380
rect 47610 17436 47918 17445
rect 47610 17434 47616 17436
rect 47672 17434 47696 17436
rect 47752 17434 47776 17436
rect 47832 17434 47856 17436
rect 47912 17434 47918 17436
rect 47672 17382 47674 17434
rect 47854 17382 47856 17434
rect 47610 17380 47616 17382
rect 47672 17380 47696 17382
rect 47752 17380 47776 17382
rect 47832 17380 47856 17382
rect 47912 17380 47918 17382
rect 47610 17371 47918 17380
rect 52610 17436 52918 17445
rect 52610 17434 52616 17436
rect 52672 17434 52696 17436
rect 52752 17434 52776 17436
rect 52832 17434 52856 17436
rect 52912 17434 52918 17436
rect 52672 17382 52674 17434
rect 52854 17382 52856 17434
rect 52610 17380 52616 17382
rect 52672 17380 52696 17382
rect 52752 17380 52776 17382
rect 52832 17380 52856 17382
rect 52912 17380 52918 17382
rect 52610 17371 52918 17380
rect 57610 17436 57918 17445
rect 57610 17434 57616 17436
rect 57672 17434 57696 17436
rect 57752 17434 57776 17436
rect 57832 17434 57856 17436
rect 57912 17434 57918 17436
rect 57672 17382 57674 17434
rect 57854 17382 57856 17434
rect 57610 17380 57616 17382
rect 57672 17380 57696 17382
rect 57752 17380 57776 17382
rect 57832 17380 57856 17382
rect 57912 17380 57918 17382
rect 57610 17371 57918 17380
rect 58544 17241 58572 17614
rect 58530 17232 58586 17241
rect 58530 17167 58586 17176
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 11950 16892 12258 16901
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 21950 16892 22258 16901
rect 21950 16890 21956 16892
rect 22012 16890 22036 16892
rect 22092 16890 22116 16892
rect 22172 16890 22196 16892
rect 22252 16890 22258 16892
rect 22012 16838 22014 16890
rect 22194 16838 22196 16890
rect 21950 16836 21956 16838
rect 22012 16836 22036 16838
rect 22092 16836 22116 16838
rect 22172 16836 22196 16838
rect 22252 16836 22258 16838
rect 21950 16827 22258 16836
rect 26950 16892 27258 16901
rect 26950 16890 26956 16892
rect 27012 16890 27036 16892
rect 27092 16890 27116 16892
rect 27172 16890 27196 16892
rect 27252 16890 27258 16892
rect 27012 16838 27014 16890
rect 27194 16838 27196 16890
rect 26950 16836 26956 16838
rect 27012 16836 27036 16838
rect 27092 16836 27116 16838
rect 27172 16836 27196 16838
rect 27252 16836 27258 16838
rect 26950 16827 27258 16836
rect 31950 16892 32258 16901
rect 31950 16890 31956 16892
rect 32012 16890 32036 16892
rect 32092 16890 32116 16892
rect 32172 16890 32196 16892
rect 32252 16890 32258 16892
rect 32012 16838 32014 16890
rect 32194 16838 32196 16890
rect 31950 16836 31956 16838
rect 32012 16836 32036 16838
rect 32092 16836 32116 16838
rect 32172 16836 32196 16838
rect 32252 16836 32258 16838
rect 31950 16827 32258 16836
rect 36950 16892 37258 16901
rect 36950 16890 36956 16892
rect 37012 16890 37036 16892
rect 37092 16890 37116 16892
rect 37172 16890 37196 16892
rect 37252 16890 37258 16892
rect 37012 16838 37014 16890
rect 37194 16838 37196 16890
rect 36950 16836 36956 16838
rect 37012 16836 37036 16838
rect 37092 16836 37116 16838
rect 37172 16836 37196 16838
rect 37252 16836 37258 16838
rect 36950 16827 37258 16836
rect 41950 16892 42258 16901
rect 41950 16890 41956 16892
rect 42012 16890 42036 16892
rect 42092 16890 42116 16892
rect 42172 16890 42196 16892
rect 42252 16890 42258 16892
rect 42012 16838 42014 16890
rect 42194 16838 42196 16890
rect 41950 16836 41956 16838
rect 42012 16836 42036 16838
rect 42092 16836 42116 16838
rect 42172 16836 42196 16838
rect 42252 16836 42258 16838
rect 41950 16827 42258 16836
rect 46950 16892 47258 16901
rect 46950 16890 46956 16892
rect 47012 16890 47036 16892
rect 47092 16890 47116 16892
rect 47172 16890 47196 16892
rect 47252 16890 47258 16892
rect 47012 16838 47014 16890
rect 47194 16838 47196 16890
rect 46950 16836 46956 16838
rect 47012 16836 47036 16838
rect 47092 16836 47116 16838
rect 47172 16836 47196 16838
rect 47252 16836 47258 16838
rect 46950 16827 47258 16836
rect 51950 16892 52258 16901
rect 51950 16890 51956 16892
rect 52012 16890 52036 16892
rect 52092 16890 52116 16892
rect 52172 16890 52196 16892
rect 52252 16890 52258 16892
rect 52012 16838 52014 16890
rect 52194 16838 52196 16890
rect 51950 16836 51956 16838
rect 52012 16836 52036 16838
rect 52092 16836 52116 16838
rect 52172 16836 52196 16838
rect 52252 16836 52258 16838
rect 51950 16827 52258 16836
rect 56950 16892 57258 16901
rect 56950 16890 56956 16892
rect 57012 16890 57036 16892
rect 57092 16890 57116 16892
rect 57172 16890 57196 16892
rect 57252 16890 57258 16892
rect 57012 16838 57014 16890
rect 57194 16838 57196 16890
rect 56950 16836 56956 16838
rect 57012 16836 57036 16838
rect 57092 16836 57116 16838
rect 57172 16836 57196 16838
rect 57252 16836 57258 16838
rect 56950 16827 57258 16836
rect 57980 16652 58032 16658
rect 57980 16594 58032 16600
rect 57886 16552 57942 16561
rect 57992 16538 58020 16594
rect 57942 16510 58020 16538
rect 57886 16487 57942 16496
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 7610 16348 7918 16357
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7610 16283 7918 16292
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 17610 16348 17918 16357
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 22610 16348 22918 16357
rect 22610 16346 22616 16348
rect 22672 16346 22696 16348
rect 22752 16346 22776 16348
rect 22832 16346 22856 16348
rect 22912 16346 22918 16348
rect 22672 16294 22674 16346
rect 22854 16294 22856 16346
rect 22610 16292 22616 16294
rect 22672 16292 22696 16294
rect 22752 16292 22776 16294
rect 22832 16292 22856 16294
rect 22912 16292 22918 16294
rect 22610 16283 22918 16292
rect 27610 16348 27918 16357
rect 27610 16346 27616 16348
rect 27672 16346 27696 16348
rect 27752 16346 27776 16348
rect 27832 16346 27856 16348
rect 27912 16346 27918 16348
rect 27672 16294 27674 16346
rect 27854 16294 27856 16346
rect 27610 16292 27616 16294
rect 27672 16292 27696 16294
rect 27752 16292 27776 16294
rect 27832 16292 27856 16294
rect 27912 16292 27918 16294
rect 27610 16283 27918 16292
rect 32610 16348 32918 16357
rect 32610 16346 32616 16348
rect 32672 16346 32696 16348
rect 32752 16346 32776 16348
rect 32832 16346 32856 16348
rect 32912 16346 32918 16348
rect 32672 16294 32674 16346
rect 32854 16294 32856 16346
rect 32610 16292 32616 16294
rect 32672 16292 32696 16294
rect 32752 16292 32776 16294
rect 32832 16292 32856 16294
rect 32912 16292 32918 16294
rect 32610 16283 32918 16292
rect 37610 16348 37918 16357
rect 37610 16346 37616 16348
rect 37672 16346 37696 16348
rect 37752 16346 37776 16348
rect 37832 16346 37856 16348
rect 37912 16346 37918 16348
rect 37672 16294 37674 16346
rect 37854 16294 37856 16346
rect 37610 16292 37616 16294
rect 37672 16292 37696 16294
rect 37752 16292 37776 16294
rect 37832 16292 37856 16294
rect 37912 16292 37918 16294
rect 37610 16283 37918 16292
rect 42610 16348 42918 16357
rect 42610 16346 42616 16348
rect 42672 16346 42696 16348
rect 42752 16346 42776 16348
rect 42832 16346 42856 16348
rect 42912 16346 42918 16348
rect 42672 16294 42674 16346
rect 42854 16294 42856 16346
rect 42610 16292 42616 16294
rect 42672 16292 42696 16294
rect 42752 16292 42776 16294
rect 42832 16292 42856 16294
rect 42912 16292 42918 16294
rect 42610 16283 42918 16292
rect 47610 16348 47918 16357
rect 47610 16346 47616 16348
rect 47672 16346 47696 16348
rect 47752 16346 47776 16348
rect 47832 16346 47856 16348
rect 47912 16346 47918 16348
rect 47672 16294 47674 16346
rect 47854 16294 47856 16346
rect 47610 16292 47616 16294
rect 47672 16292 47696 16294
rect 47752 16292 47776 16294
rect 47832 16292 47856 16294
rect 47912 16292 47918 16294
rect 47610 16283 47918 16292
rect 52610 16348 52918 16357
rect 52610 16346 52616 16348
rect 52672 16346 52696 16348
rect 52752 16346 52776 16348
rect 52832 16346 52856 16348
rect 52912 16346 52918 16348
rect 52672 16294 52674 16346
rect 52854 16294 52856 16346
rect 52610 16292 52616 16294
rect 52672 16292 52696 16294
rect 52752 16292 52776 16294
rect 52832 16292 52856 16294
rect 52912 16292 52918 16294
rect 52610 16283 52918 16292
rect 57610 16348 57918 16357
rect 57610 16346 57616 16348
rect 57672 16346 57696 16348
rect 57752 16346 57776 16348
rect 57832 16346 57856 16348
rect 57912 16346 57918 16348
rect 57672 16294 57674 16346
rect 57854 16294 57856 16346
rect 57610 16292 57616 16294
rect 57672 16292 57696 16294
rect 57752 16292 57776 16294
rect 57832 16292 57856 16294
rect 57912 16292 57918 16294
rect 57610 16283 57918 16292
rect 58532 15904 58584 15910
rect 58532 15846 58584 15852
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 21950 15804 22258 15813
rect 21950 15802 21956 15804
rect 22012 15802 22036 15804
rect 22092 15802 22116 15804
rect 22172 15802 22196 15804
rect 22252 15802 22258 15804
rect 22012 15750 22014 15802
rect 22194 15750 22196 15802
rect 21950 15748 21956 15750
rect 22012 15748 22036 15750
rect 22092 15748 22116 15750
rect 22172 15748 22196 15750
rect 22252 15748 22258 15750
rect 21950 15739 22258 15748
rect 26950 15804 27258 15813
rect 26950 15802 26956 15804
rect 27012 15802 27036 15804
rect 27092 15802 27116 15804
rect 27172 15802 27196 15804
rect 27252 15802 27258 15804
rect 27012 15750 27014 15802
rect 27194 15750 27196 15802
rect 26950 15748 26956 15750
rect 27012 15748 27036 15750
rect 27092 15748 27116 15750
rect 27172 15748 27196 15750
rect 27252 15748 27258 15750
rect 26950 15739 27258 15748
rect 31950 15804 32258 15813
rect 31950 15802 31956 15804
rect 32012 15802 32036 15804
rect 32092 15802 32116 15804
rect 32172 15802 32196 15804
rect 32252 15802 32258 15804
rect 32012 15750 32014 15802
rect 32194 15750 32196 15802
rect 31950 15748 31956 15750
rect 32012 15748 32036 15750
rect 32092 15748 32116 15750
rect 32172 15748 32196 15750
rect 32252 15748 32258 15750
rect 31950 15739 32258 15748
rect 36950 15804 37258 15813
rect 36950 15802 36956 15804
rect 37012 15802 37036 15804
rect 37092 15802 37116 15804
rect 37172 15802 37196 15804
rect 37252 15802 37258 15804
rect 37012 15750 37014 15802
rect 37194 15750 37196 15802
rect 36950 15748 36956 15750
rect 37012 15748 37036 15750
rect 37092 15748 37116 15750
rect 37172 15748 37196 15750
rect 37252 15748 37258 15750
rect 36950 15739 37258 15748
rect 41950 15804 42258 15813
rect 41950 15802 41956 15804
rect 42012 15802 42036 15804
rect 42092 15802 42116 15804
rect 42172 15802 42196 15804
rect 42252 15802 42258 15804
rect 42012 15750 42014 15802
rect 42194 15750 42196 15802
rect 41950 15748 41956 15750
rect 42012 15748 42036 15750
rect 42092 15748 42116 15750
rect 42172 15748 42196 15750
rect 42252 15748 42258 15750
rect 41950 15739 42258 15748
rect 46950 15804 47258 15813
rect 46950 15802 46956 15804
rect 47012 15802 47036 15804
rect 47092 15802 47116 15804
rect 47172 15802 47196 15804
rect 47252 15802 47258 15804
rect 47012 15750 47014 15802
rect 47194 15750 47196 15802
rect 46950 15748 46956 15750
rect 47012 15748 47036 15750
rect 47092 15748 47116 15750
rect 47172 15748 47196 15750
rect 47252 15748 47258 15750
rect 46950 15739 47258 15748
rect 51950 15804 52258 15813
rect 51950 15802 51956 15804
rect 52012 15802 52036 15804
rect 52092 15802 52116 15804
rect 52172 15802 52196 15804
rect 52252 15802 52258 15804
rect 52012 15750 52014 15802
rect 52194 15750 52196 15802
rect 51950 15748 51956 15750
rect 52012 15748 52036 15750
rect 52092 15748 52116 15750
rect 52172 15748 52196 15750
rect 52252 15748 52258 15750
rect 51950 15739 52258 15748
rect 56950 15804 57258 15813
rect 56950 15802 56956 15804
rect 57012 15802 57036 15804
rect 57092 15802 57116 15804
rect 57172 15802 57196 15804
rect 57252 15802 57258 15804
rect 57012 15750 57014 15802
rect 57194 15750 57196 15802
rect 56950 15748 56956 15750
rect 57012 15748 57036 15750
rect 57092 15748 57116 15750
rect 57172 15748 57196 15750
rect 57252 15748 57258 15750
rect 56950 15739 57258 15748
rect 58544 15609 58572 15846
rect 58530 15600 58586 15609
rect 58530 15535 58586 15544
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 17610 15260 17918 15269
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 22610 15260 22918 15269
rect 22610 15258 22616 15260
rect 22672 15258 22696 15260
rect 22752 15258 22776 15260
rect 22832 15258 22856 15260
rect 22912 15258 22918 15260
rect 22672 15206 22674 15258
rect 22854 15206 22856 15258
rect 22610 15204 22616 15206
rect 22672 15204 22696 15206
rect 22752 15204 22776 15206
rect 22832 15204 22856 15206
rect 22912 15204 22918 15206
rect 22610 15195 22918 15204
rect 27610 15260 27918 15269
rect 27610 15258 27616 15260
rect 27672 15258 27696 15260
rect 27752 15258 27776 15260
rect 27832 15258 27856 15260
rect 27912 15258 27918 15260
rect 27672 15206 27674 15258
rect 27854 15206 27856 15258
rect 27610 15204 27616 15206
rect 27672 15204 27696 15206
rect 27752 15204 27776 15206
rect 27832 15204 27856 15206
rect 27912 15204 27918 15206
rect 27610 15195 27918 15204
rect 32610 15260 32918 15269
rect 32610 15258 32616 15260
rect 32672 15258 32696 15260
rect 32752 15258 32776 15260
rect 32832 15258 32856 15260
rect 32912 15258 32918 15260
rect 32672 15206 32674 15258
rect 32854 15206 32856 15258
rect 32610 15204 32616 15206
rect 32672 15204 32696 15206
rect 32752 15204 32776 15206
rect 32832 15204 32856 15206
rect 32912 15204 32918 15206
rect 32610 15195 32918 15204
rect 37610 15260 37918 15269
rect 37610 15258 37616 15260
rect 37672 15258 37696 15260
rect 37752 15258 37776 15260
rect 37832 15258 37856 15260
rect 37912 15258 37918 15260
rect 37672 15206 37674 15258
rect 37854 15206 37856 15258
rect 37610 15204 37616 15206
rect 37672 15204 37696 15206
rect 37752 15204 37776 15206
rect 37832 15204 37856 15206
rect 37912 15204 37918 15206
rect 37610 15195 37918 15204
rect 42610 15260 42918 15269
rect 42610 15258 42616 15260
rect 42672 15258 42696 15260
rect 42752 15258 42776 15260
rect 42832 15258 42856 15260
rect 42912 15258 42918 15260
rect 42672 15206 42674 15258
rect 42854 15206 42856 15258
rect 42610 15204 42616 15206
rect 42672 15204 42696 15206
rect 42752 15204 42776 15206
rect 42832 15204 42856 15206
rect 42912 15204 42918 15206
rect 42610 15195 42918 15204
rect 47610 15260 47918 15269
rect 47610 15258 47616 15260
rect 47672 15258 47696 15260
rect 47752 15258 47776 15260
rect 47832 15258 47856 15260
rect 47912 15258 47918 15260
rect 47672 15206 47674 15258
rect 47854 15206 47856 15258
rect 47610 15204 47616 15206
rect 47672 15204 47696 15206
rect 47752 15204 47776 15206
rect 47832 15204 47856 15206
rect 47912 15204 47918 15206
rect 47610 15195 47918 15204
rect 52610 15260 52918 15269
rect 52610 15258 52616 15260
rect 52672 15258 52696 15260
rect 52752 15258 52776 15260
rect 52832 15258 52856 15260
rect 52912 15258 52918 15260
rect 52672 15206 52674 15258
rect 52854 15206 52856 15258
rect 52610 15204 52616 15206
rect 52672 15204 52696 15206
rect 52752 15204 52776 15206
rect 52832 15204 52856 15206
rect 52912 15204 52918 15206
rect 52610 15195 52918 15204
rect 57610 15260 57918 15269
rect 57610 15258 57616 15260
rect 57672 15258 57696 15260
rect 57752 15258 57776 15260
rect 57832 15258 57856 15260
rect 57912 15258 57918 15260
rect 57672 15206 57674 15258
rect 57854 15206 57856 15258
rect 57610 15204 57616 15206
rect 57672 15204 57696 15206
rect 57752 15204 57776 15206
rect 57832 15204 57856 15206
rect 57912 15204 57918 15206
rect 57610 15195 57918 15204
rect 58532 14816 58584 14822
rect 58530 14784 58532 14793
rect 58584 14784 58586 14793
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 21950 14716 22258 14725
rect 21950 14714 21956 14716
rect 22012 14714 22036 14716
rect 22092 14714 22116 14716
rect 22172 14714 22196 14716
rect 22252 14714 22258 14716
rect 22012 14662 22014 14714
rect 22194 14662 22196 14714
rect 21950 14660 21956 14662
rect 22012 14660 22036 14662
rect 22092 14660 22116 14662
rect 22172 14660 22196 14662
rect 22252 14660 22258 14662
rect 21950 14651 22258 14660
rect 26950 14716 27258 14725
rect 26950 14714 26956 14716
rect 27012 14714 27036 14716
rect 27092 14714 27116 14716
rect 27172 14714 27196 14716
rect 27252 14714 27258 14716
rect 27012 14662 27014 14714
rect 27194 14662 27196 14714
rect 26950 14660 26956 14662
rect 27012 14660 27036 14662
rect 27092 14660 27116 14662
rect 27172 14660 27196 14662
rect 27252 14660 27258 14662
rect 26950 14651 27258 14660
rect 31950 14716 32258 14725
rect 31950 14714 31956 14716
rect 32012 14714 32036 14716
rect 32092 14714 32116 14716
rect 32172 14714 32196 14716
rect 32252 14714 32258 14716
rect 32012 14662 32014 14714
rect 32194 14662 32196 14714
rect 31950 14660 31956 14662
rect 32012 14660 32036 14662
rect 32092 14660 32116 14662
rect 32172 14660 32196 14662
rect 32252 14660 32258 14662
rect 31950 14651 32258 14660
rect 36950 14716 37258 14725
rect 36950 14714 36956 14716
rect 37012 14714 37036 14716
rect 37092 14714 37116 14716
rect 37172 14714 37196 14716
rect 37252 14714 37258 14716
rect 37012 14662 37014 14714
rect 37194 14662 37196 14714
rect 36950 14660 36956 14662
rect 37012 14660 37036 14662
rect 37092 14660 37116 14662
rect 37172 14660 37196 14662
rect 37252 14660 37258 14662
rect 36950 14651 37258 14660
rect 41950 14716 42258 14725
rect 41950 14714 41956 14716
rect 42012 14714 42036 14716
rect 42092 14714 42116 14716
rect 42172 14714 42196 14716
rect 42252 14714 42258 14716
rect 42012 14662 42014 14714
rect 42194 14662 42196 14714
rect 41950 14660 41956 14662
rect 42012 14660 42036 14662
rect 42092 14660 42116 14662
rect 42172 14660 42196 14662
rect 42252 14660 42258 14662
rect 41950 14651 42258 14660
rect 46950 14716 47258 14725
rect 46950 14714 46956 14716
rect 47012 14714 47036 14716
rect 47092 14714 47116 14716
rect 47172 14714 47196 14716
rect 47252 14714 47258 14716
rect 47012 14662 47014 14714
rect 47194 14662 47196 14714
rect 46950 14660 46956 14662
rect 47012 14660 47036 14662
rect 47092 14660 47116 14662
rect 47172 14660 47196 14662
rect 47252 14660 47258 14662
rect 46950 14651 47258 14660
rect 51950 14716 52258 14725
rect 51950 14714 51956 14716
rect 52012 14714 52036 14716
rect 52092 14714 52116 14716
rect 52172 14714 52196 14716
rect 52252 14714 52258 14716
rect 52012 14662 52014 14714
rect 52194 14662 52196 14714
rect 51950 14660 51956 14662
rect 52012 14660 52036 14662
rect 52092 14660 52116 14662
rect 52172 14660 52196 14662
rect 52252 14660 52258 14662
rect 51950 14651 52258 14660
rect 56950 14716 57258 14725
rect 58530 14719 58586 14728
rect 56950 14714 56956 14716
rect 57012 14714 57036 14716
rect 57092 14714 57116 14716
rect 57172 14714 57196 14716
rect 57252 14714 57258 14716
rect 57012 14662 57014 14714
rect 57194 14662 57196 14714
rect 56950 14660 56956 14662
rect 57012 14660 57036 14662
rect 57092 14660 57116 14662
rect 57172 14660 57196 14662
rect 57252 14660 57258 14662
rect 56950 14651 57258 14660
rect 58532 14408 58584 14414
rect 58532 14350 58584 14356
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 17610 14172 17918 14181
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 22610 14172 22918 14181
rect 22610 14170 22616 14172
rect 22672 14170 22696 14172
rect 22752 14170 22776 14172
rect 22832 14170 22856 14172
rect 22912 14170 22918 14172
rect 22672 14118 22674 14170
rect 22854 14118 22856 14170
rect 22610 14116 22616 14118
rect 22672 14116 22696 14118
rect 22752 14116 22776 14118
rect 22832 14116 22856 14118
rect 22912 14116 22918 14118
rect 22610 14107 22918 14116
rect 27610 14172 27918 14181
rect 27610 14170 27616 14172
rect 27672 14170 27696 14172
rect 27752 14170 27776 14172
rect 27832 14170 27856 14172
rect 27912 14170 27918 14172
rect 27672 14118 27674 14170
rect 27854 14118 27856 14170
rect 27610 14116 27616 14118
rect 27672 14116 27696 14118
rect 27752 14116 27776 14118
rect 27832 14116 27856 14118
rect 27912 14116 27918 14118
rect 27610 14107 27918 14116
rect 32610 14172 32918 14181
rect 32610 14170 32616 14172
rect 32672 14170 32696 14172
rect 32752 14170 32776 14172
rect 32832 14170 32856 14172
rect 32912 14170 32918 14172
rect 32672 14118 32674 14170
rect 32854 14118 32856 14170
rect 32610 14116 32616 14118
rect 32672 14116 32696 14118
rect 32752 14116 32776 14118
rect 32832 14116 32856 14118
rect 32912 14116 32918 14118
rect 32610 14107 32918 14116
rect 37610 14172 37918 14181
rect 37610 14170 37616 14172
rect 37672 14170 37696 14172
rect 37752 14170 37776 14172
rect 37832 14170 37856 14172
rect 37912 14170 37918 14172
rect 37672 14118 37674 14170
rect 37854 14118 37856 14170
rect 37610 14116 37616 14118
rect 37672 14116 37696 14118
rect 37752 14116 37776 14118
rect 37832 14116 37856 14118
rect 37912 14116 37918 14118
rect 37610 14107 37918 14116
rect 42610 14172 42918 14181
rect 42610 14170 42616 14172
rect 42672 14170 42696 14172
rect 42752 14170 42776 14172
rect 42832 14170 42856 14172
rect 42912 14170 42918 14172
rect 42672 14118 42674 14170
rect 42854 14118 42856 14170
rect 42610 14116 42616 14118
rect 42672 14116 42696 14118
rect 42752 14116 42776 14118
rect 42832 14116 42856 14118
rect 42912 14116 42918 14118
rect 42610 14107 42918 14116
rect 47610 14172 47918 14181
rect 47610 14170 47616 14172
rect 47672 14170 47696 14172
rect 47752 14170 47776 14172
rect 47832 14170 47856 14172
rect 47912 14170 47918 14172
rect 47672 14118 47674 14170
rect 47854 14118 47856 14170
rect 47610 14116 47616 14118
rect 47672 14116 47696 14118
rect 47752 14116 47776 14118
rect 47832 14116 47856 14118
rect 47912 14116 47918 14118
rect 47610 14107 47918 14116
rect 52610 14172 52918 14181
rect 52610 14170 52616 14172
rect 52672 14170 52696 14172
rect 52752 14170 52776 14172
rect 52832 14170 52856 14172
rect 52912 14170 52918 14172
rect 52672 14118 52674 14170
rect 52854 14118 52856 14170
rect 52610 14116 52616 14118
rect 52672 14116 52696 14118
rect 52752 14116 52776 14118
rect 52832 14116 52856 14118
rect 52912 14116 52918 14118
rect 52610 14107 52918 14116
rect 57610 14172 57918 14181
rect 57610 14170 57616 14172
rect 57672 14170 57696 14172
rect 57752 14170 57776 14172
rect 57832 14170 57856 14172
rect 57912 14170 57918 14172
rect 57672 14118 57674 14170
rect 57854 14118 57856 14170
rect 57610 14116 57616 14118
rect 57672 14116 57696 14118
rect 57752 14116 57776 14118
rect 57832 14116 57856 14118
rect 57912 14116 57918 14118
rect 57610 14107 57918 14116
rect 58544 13977 58572 14350
rect 58530 13968 58586 13977
rect 58530 13903 58586 13912
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 21950 13628 22258 13637
rect 21950 13626 21956 13628
rect 22012 13626 22036 13628
rect 22092 13626 22116 13628
rect 22172 13626 22196 13628
rect 22252 13626 22258 13628
rect 22012 13574 22014 13626
rect 22194 13574 22196 13626
rect 21950 13572 21956 13574
rect 22012 13572 22036 13574
rect 22092 13572 22116 13574
rect 22172 13572 22196 13574
rect 22252 13572 22258 13574
rect 21950 13563 22258 13572
rect 26950 13628 27258 13637
rect 26950 13626 26956 13628
rect 27012 13626 27036 13628
rect 27092 13626 27116 13628
rect 27172 13626 27196 13628
rect 27252 13626 27258 13628
rect 27012 13574 27014 13626
rect 27194 13574 27196 13626
rect 26950 13572 26956 13574
rect 27012 13572 27036 13574
rect 27092 13572 27116 13574
rect 27172 13572 27196 13574
rect 27252 13572 27258 13574
rect 26950 13563 27258 13572
rect 31950 13628 32258 13637
rect 31950 13626 31956 13628
rect 32012 13626 32036 13628
rect 32092 13626 32116 13628
rect 32172 13626 32196 13628
rect 32252 13626 32258 13628
rect 32012 13574 32014 13626
rect 32194 13574 32196 13626
rect 31950 13572 31956 13574
rect 32012 13572 32036 13574
rect 32092 13572 32116 13574
rect 32172 13572 32196 13574
rect 32252 13572 32258 13574
rect 31950 13563 32258 13572
rect 36950 13628 37258 13637
rect 36950 13626 36956 13628
rect 37012 13626 37036 13628
rect 37092 13626 37116 13628
rect 37172 13626 37196 13628
rect 37252 13626 37258 13628
rect 37012 13574 37014 13626
rect 37194 13574 37196 13626
rect 36950 13572 36956 13574
rect 37012 13572 37036 13574
rect 37092 13572 37116 13574
rect 37172 13572 37196 13574
rect 37252 13572 37258 13574
rect 36950 13563 37258 13572
rect 41950 13628 42258 13637
rect 41950 13626 41956 13628
rect 42012 13626 42036 13628
rect 42092 13626 42116 13628
rect 42172 13626 42196 13628
rect 42252 13626 42258 13628
rect 42012 13574 42014 13626
rect 42194 13574 42196 13626
rect 41950 13572 41956 13574
rect 42012 13572 42036 13574
rect 42092 13572 42116 13574
rect 42172 13572 42196 13574
rect 42252 13572 42258 13574
rect 41950 13563 42258 13572
rect 46950 13628 47258 13637
rect 46950 13626 46956 13628
rect 47012 13626 47036 13628
rect 47092 13626 47116 13628
rect 47172 13626 47196 13628
rect 47252 13626 47258 13628
rect 47012 13574 47014 13626
rect 47194 13574 47196 13626
rect 46950 13572 46956 13574
rect 47012 13572 47036 13574
rect 47092 13572 47116 13574
rect 47172 13572 47196 13574
rect 47252 13572 47258 13574
rect 46950 13563 47258 13572
rect 51950 13628 52258 13637
rect 51950 13626 51956 13628
rect 52012 13626 52036 13628
rect 52092 13626 52116 13628
rect 52172 13626 52196 13628
rect 52252 13626 52258 13628
rect 52012 13574 52014 13626
rect 52194 13574 52196 13626
rect 51950 13572 51956 13574
rect 52012 13572 52036 13574
rect 52092 13572 52116 13574
rect 52172 13572 52196 13574
rect 52252 13572 52258 13574
rect 51950 13563 52258 13572
rect 56950 13628 57258 13637
rect 56950 13626 56956 13628
rect 57012 13626 57036 13628
rect 57092 13626 57116 13628
rect 57172 13626 57196 13628
rect 57252 13626 57258 13628
rect 57012 13574 57014 13626
rect 57194 13574 57196 13626
rect 56950 13572 56956 13574
rect 57012 13572 57036 13574
rect 57092 13572 57116 13574
rect 57172 13572 57196 13574
rect 57252 13572 57258 13574
rect 56950 13563 57258 13572
rect 58532 13320 58584 13326
rect 58532 13262 58584 13268
rect 58544 13161 58572 13262
rect 58530 13152 58586 13161
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 22610 13084 22918 13093
rect 22610 13082 22616 13084
rect 22672 13082 22696 13084
rect 22752 13082 22776 13084
rect 22832 13082 22856 13084
rect 22912 13082 22918 13084
rect 22672 13030 22674 13082
rect 22854 13030 22856 13082
rect 22610 13028 22616 13030
rect 22672 13028 22696 13030
rect 22752 13028 22776 13030
rect 22832 13028 22856 13030
rect 22912 13028 22918 13030
rect 22610 13019 22918 13028
rect 27610 13084 27918 13093
rect 27610 13082 27616 13084
rect 27672 13082 27696 13084
rect 27752 13082 27776 13084
rect 27832 13082 27856 13084
rect 27912 13082 27918 13084
rect 27672 13030 27674 13082
rect 27854 13030 27856 13082
rect 27610 13028 27616 13030
rect 27672 13028 27696 13030
rect 27752 13028 27776 13030
rect 27832 13028 27856 13030
rect 27912 13028 27918 13030
rect 27610 13019 27918 13028
rect 32610 13084 32918 13093
rect 32610 13082 32616 13084
rect 32672 13082 32696 13084
rect 32752 13082 32776 13084
rect 32832 13082 32856 13084
rect 32912 13082 32918 13084
rect 32672 13030 32674 13082
rect 32854 13030 32856 13082
rect 32610 13028 32616 13030
rect 32672 13028 32696 13030
rect 32752 13028 32776 13030
rect 32832 13028 32856 13030
rect 32912 13028 32918 13030
rect 32610 13019 32918 13028
rect 37610 13084 37918 13093
rect 37610 13082 37616 13084
rect 37672 13082 37696 13084
rect 37752 13082 37776 13084
rect 37832 13082 37856 13084
rect 37912 13082 37918 13084
rect 37672 13030 37674 13082
rect 37854 13030 37856 13082
rect 37610 13028 37616 13030
rect 37672 13028 37696 13030
rect 37752 13028 37776 13030
rect 37832 13028 37856 13030
rect 37912 13028 37918 13030
rect 37610 13019 37918 13028
rect 42610 13084 42918 13093
rect 42610 13082 42616 13084
rect 42672 13082 42696 13084
rect 42752 13082 42776 13084
rect 42832 13082 42856 13084
rect 42912 13082 42918 13084
rect 42672 13030 42674 13082
rect 42854 13030 42856 13082
rect 42610 13028 42616 13030
rect 42672 13028 42696 13030
rect 42752 13028 42776 13030
rect 42832 13028 42856 13030
rect 42912 13028 42918 13030
rect 42610 13019 42918 13028
rect 47610 13084 47918 13093
rect 47610 13082 47616 13084
rect 47672 13082 47696 13084
rect 47752 13082 47776 13084
rect 47832 13082 47856 13084
rect 47912 13082 47918 13084
rect 47672 13030 47674 13082
rect 47854 13030 47856 13082
rect 47610 13028 47616 13030
rect 47672 13028 47696 13030
rect 47752 13028 47776 13030
rect 47832 13028 47856 13030
rect 47912 13028 47918 13030
rect 47610 13019 47918 13028
rect 52610 13084 52918 13093
rect 52610 13082 52616 13084
rect 52672 13082 52696 13084
rect 52752 13082 52776 13084
rect 52832 13082 52856 13084
rect 52912 13082 52918 13084
rect 52672 13030 52674 13082
rect 52854 13030 52856 13082
rect 52610 13028 52616 13030
rect 52672 13028 52696 13030
rect 52752 13028 52776 13030
rect 52832 13028 52856 13030
rect 52912 13028 52918 13030
rect 52610 13019 52918 13028
rect 57610 13084 57918 13093
rect 58530 13087 58586 13096
rect 57610 13082 57616 13084
rect 57672 13082 57696 13084
rect 57752 13082 57776 13084
rect 57832 13082 57856 13084
rect 57912 13082 57918 13084
rect 57672 13030 57674 13082
rect 57854 13030 57856 13082
rect 57610 13028 57616 13030
rect 57672 13028 57696 13030
rect 57752 13028 57776 13030
rect 57832 13028 57856 13030
rect 57912 13028 57918 13030
rect 57610 13019 57918 13028
rect 58532 12640 58584 12646
rect 58532 12582 58584 12588
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 21950 12540 22258 12549
rect 21950 12538 21956 12540
rect 22012 12538 22036 12540
rect 22092 12538 22116 12540
rect 22172 12538 22196 12540
rect 22252 12538 22258 12540
rect 22012 12486 22014 12538
rect 22194 12486 22196 12538
rect 21950 12484 21956 12486
rect 22012 12484 22036 12486
rect 22092 12484 22116 12486
rect 22172 12484 22196 12486
rect 22252 12484 22258 12486
rect 21950 12475 22258 12484
rect 26950 12540 27258 12549
rect 26950 12538 26956 12540
rect 27012 12538 27036 12540
rect 27092 12538 27116 12540
rect 27172 12538 27196 12540
rect 27252 12538 27258 12540
rect 27012 12486 27014 12538
rect 27194 12486 27196 12538
rect 26950 12484 26956 12486
rect 27012 12484 27036 12486
rect 27092 12484 27116 12486
rect 27172 12484 27196 12486
rect 27252 12484 27258 12486
rect 26950 12475 27258 12484
rect 31950 12540 32258 12549
rect 31950 12538 31956 12540
rect 32012 12538 32036 12540
rect 32092 12538 32116 12540
rect 32172 12538 32196 12540
rect 32252 12538 32258 12540
rect 32012 12486 32014 12538
rect 32194 12486 32196 12538
rect 31950 12484 31956 12486
rect 32012 12484 32036 12486
rect 32092 12484 32116 12486
rect 32172 12484 32196 12486
rect 32252 12484 32258 12486
rect 31950 12475 32258 12484
rect 36950 12540 37258 12549
rect 36950 12538 36956 12540
rect 37012 12538 37036 12540
rect 37092 12538 37116 12540
rect 37172 12538 37196 12540
rect 37252 12538 37258 12540
rect 37012 12486 37014 12538
rect 37194 12486 37196 12538
rect 36950 12484 36956 12486
rect 37012 12484 37036 12486
rect 37092 12484 37116 12486
rect 37172 12484 37196 12486
rect 37252 12484 37258 12486
rect 36950 12475 37258 12484
rect 41950 12540 42258 12549
rect 41950 12538 41956 12540
rect 42012 12538 42036 12540
rect 42092 12538 42116 12540
rect 42172 12538 42196 12540
rect 42252 12538 42258 12540
rect 42012 12486 42014 12538
rect 42194 12486 42196 12538
rect 41950 12484 41956 12486
rect 42012 12484 42036 12486
rect 42092 12484 42116 12486
rect 42172 12484 42196 12486
rect 42252 12484 42258 12486
rect 41950 12475 42258 12484
rect 46950 12540 47258 12549
rect 46950 12538 46956 12540
rect 47012 12538 47036 12540
rect 47092 12538 47116 12540
rect 47172 12538 47196 12540
rect 47252 12538 47258 12540
rect 47012 12486 47014 12538
rect 47194 12486 47196 12538
rect 46950 12484 46956 12486
rect 47012 12484 47036 12486
rect 47092 12484 47116 12486
rect 47172 12484 47196 12486
rect 47252 12484 47258 12486
rect 46950 12475 47258 12484
rect 51950 12540 52258 12549
rect 51950 12538 51956 12540
rect 52012 12538 52036 12540
rect 52092 12538 52116 12540
rect 52172 12538 52196 12540
rect 52252 12538 52258 12540
rect 52012 12486 52014 12538
rect 52194 12486 52196 12538
rect 51950 12484 51956 12486
rect 52012 12484 52036 12486
rect 52092 12484 52116 12486
rect 52172 12484 52196 12486
rect 52252 12484 52258 12486
rect 51950 12475 52258 12484
rect 56950 12540 57258 12549
rect 56950 12538 56956 12540
rect 57012 12538 57036 12540
rect 57092 12538 57116 12540
rect 57172 12538 57196 12540
rect 57252 12538 57258 12540
rect 57012 12486 57014 12538
rect 57194 12486 57196 12538
rect 56950 12484 56956 12486
rect 57012 12484 57036 12486
rect 57092 12484 57116 12486
rect 57172 12484 57196 12486
rect 57252 12484 57258 12486
rect 56950 12475 57258 12484
rect 58544 12345 58572 12582
rect 58530 12336 58586 12345
rect 58530 12271 58586 12280
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 22610 11996 22918 12005
rect 22610 11994 22616 11996
rect 22672 11994 22696 11996
rect 22752 11994 22776 11996
rect 22832 11994 22856 11996
rect 22912 11994 22918 11996
rect 22672 11942 22674 11994
rect 22854 11942 22856 11994
rect 22610 11940 22616 11942
rect 22672 11940 22696 11942
rect 22752 11940 22776 11942
rect 22832 11940 22856 11942
rect 22912 11940 22918 11942
rect 22610 11931 22918 11940
rect 27610 11996 27918 12005
rect 27610 11994 27616 11996
rect 27672 11994 27696 11996
rect 27752 11994 27776 11996
rect 27832 11994 27856 11996
rect 27912 11994 27918 11996
rect 27672 11942 27674 11994
rect 27854 11942 27856 11994
rect 27610 11940 27616 11942
rect 27672 11940 27696 11942
rect 27752 11940 27776 11942
rect 27832 11940 27856 11942
rect 27912 11940 27918 11942
rect 27610 11931 27918 11940
rect 32610 11996 32918 12005
rect 32610 11994 32616 11996
rect 32672 11994 32696 11996
rect 32752 11994 32776 11996
rect 32832 11994 32856 11996
rect 32912 11994 32918 11996
rect 32672 11942 32674 11994
rect 32854 11942 32856 11994
rect 32610 11940 32616 11942
rect 32672 11940 32696 11942
rect 32752 11940 32776 11942
rect 32832 11940 32856 11942
rect 32912 11940 32918 11942
rect 32610 11931 32918 11940
rect 37610 11996 37918 12005
rect 37610 11994 37616 11996
rect 37672 11994 37696 11996
rect 37752 11994 37776 11996
rect 37832 11994 37856 11996
rect 37912 11994 37918 11996
rect 37672 11942 37674 11994
rect 37854 11942 37856 11994
rect 37610 11940 37616 11942
rect 37672 11940 37696 11942
rect 37752 11940 37776 11942
rect 37832 11940 37856 11942
rect 37912 11940 37918 11942
rect 37610 11931 37918 11940
rect 42610 11996 42918 12005
rect 42610 11994 42616 11996
rect 42672 11994 42696 11996
rect 42752 11994 42776 11996
rect 42832 11994 42856 11996
rect 42912 11994 42918 11996
rect 42672 11942 42674 11994
rect 42854 11942 42856 11994
rect 42610 11940 42616 11942
rect 42672 11940 42696 11942
rect 42752 11940 42776 11942
rect 42832 11940 42856 11942
rect 42912 11940 42918 11942
rect 42610 11931 42918 11940
rect 47610 11996 47918 12005
rect 47610 11994 47616 11996
rect 47672 11994 47696 11996
rect 47752 11994 47776 11996
rect 47832 11994 47856 11996
rect 47912 11994 47918 11996
rect 47672 11942 47674 11994
rect 47854 11942 47856 11994
rect 47610 11940 47616 11942
rect 47672 11940 47696 11942
rect 47752 11940 47776 11942
rect 47832 11940 47856 11942
rect 47912 11940 47918 11942
rect 47610 11931 47918 11940
rect 52610 11996 52918 12005
rect 52610 11994 52616 11996
rect 52672 11994 52696 11996
rect 52752 11994 52776 11996
rect 52832 11994 52856 11996
rect 52912 11994 52918 11996
rect 52672 11942 52674 11994
rect 52854 11942 52856 11994
rect 52610 11940 52616 11942
rect 52672 11940 52696 11942
rect 52752 11940 52776 11942
rect 52832 11940 52856 11942
rect 52912 11940 52918 11942
rect 52610 11931 52918 11940
rect 57610 11996 57918 12005
rect 57610 11994 57616 11996
rect 57672 11994 57696 11996
rect 57752 11994 57776 11996
rect 57832 11994 57856 11996
rect 57912 11994 57918 11996
rect 57672 11942 57674 11994
rect 57854 11942 57856 11994
rect 57610 11940 57616 11942
rect 57672 11940 57696 11942
rect 57752 11940 57776 11942
rect 57832 11940 57856 11942
rect 57912 11940 57918 11942
rect 57610 11931 57918 11940
rect 58532 11552 58584 11558
rect 58530 11520 58532 11529
rect 58584 11520 58586 11529
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 21950 11452 22258 11461
rect 21950 11450 21956 11452
rect 22012 11450 22036 11452
rect 22092 11450 22116 11452
rect 22172 11450 22196 11452
rect 22252 11450 22258 11452
rect 22012 11398 22014 11450
rect 22194 11398 22196 11450
rect 21950 11396 21956 11398
rect 22012 11396 22036 11398
rect 22092 11396 22116 11398
rect 22172 11396 22196 11398
rect 22252 11396 22258 11398
rect 21950 11387 22258 11396
rect 26950 11452 27258 11461
rect 26950 11450 26956 11452
rect 27012 11450 27036 11452
rect 27092 11450 27116 11452
rect 27172 11450 27196 11452
rect 27252 11450 27258 11452
rect 27012 11398 27014 11450
rect 27194 11398 27196 11450
rect 26950 11396 26956 11398
rect 27012 11396 27036 11398
rect 27092 11396 27116 11398
rect 27172 11396 27196 11398
rect 27252 11396 27258 11398
rect 26950 11387 27258 11396
rect 31950 11452 32258 11461
rect 31950 11450 31956 11452
rect 32012 11450 32036 11452
rect 32092 11450 32116 11452
rect 32172 11450 32196 11452
rect 32252 11450 32258 11452
rect 32012 11398 32014 11450
rect 32194 11398 32196 11450
rect 31950 11396 31956 11398
rect 32012 11396 32036 11398
rect 32092 11396 32116 11398
rect 32172 11396 32196 11398
rect 32252 11396 32258 11398
rect 31950 11387 32258 11396
rect 36950 11452 37258 11461
rect 36950 11450 36956 11452
rect 37012 11450 37036 11452
rect 37092 11450 37116 11452
rect 37172 11450 37196 11452
rect 37252 11450 37258 11452
rect 37012 11398 37014 11450
rect 37194 11398 37196 11450
rect 36950 11396 36956 11398
rect 37012 11396 37036 11398
rect 37092 11396 37116 11398
rect 37172 11396 37196 11398
rect 37252 11396 37258 11398
rect 36950 11387 37258 11396
rect 41950 11452 42258 11461
rect 41950 11450 41956 11452
rect 42012 11450 42036 11452
rect 42092 11450 42116 11452
rect 42172 11450 42196 11452
rect 42252 11450 42258 11452
rect 42012 11398 42014 11450
rect 42194 11398 42196 11450
rect 41950 11396 41956 11398
rect 42012 11396 42036 11398
rect 42092 11396 42116 11398
rect 42172 11396 42196 11398
rect 42252 11396 42258 11398
rect 41950 11387 42258 11396
rect 46950 11452 47258 11461
rect 46950 11450 46956 11452
rect 47012 11450 47036 11452
rect 47092 11450 47116 11452
rect 47172 11450 47196 11452
rect 47252 11450 47258 11452
rect 47012 11398 47014 11450
rect 47194 11398 47196 11450
rect 46950 11396 46956 11398
rect 47012 11396 47036 11398
rect 47092 11396 47116 11398
rect 47172 11396 47196 11398
rect 47252 11396 47258 11398
rect 46950 11387 47258 11396
rect 51950 11452 52258 11461
rect 51950 11450 51956 11452
rect 52012 11450 52036 11452
rect 52092 11450 52116 11452
rect 52172 11450 52196 11452
rect 52252 11450 52258 11452
rect 52012 11398 52014 11450
rect 52194 11398 52196 11450
rect 51950 11396 51956 11398
rect 52012 11396 52036 11398
rect 52092 11396 52116 11398
rect 52172 11396 52196 11398
rect 52252 11396 52258 11398
rect 51950 11387 52258 11396
rect 56950 11452 57258 11461
rect 58530 11455 58586 11464
rect 56950 11450 56956 11452
rect 57012 11450 57036 11452
rect 57092 11450 57116 11452
rect 57172 11450 57196 11452
rect 57252 11450 57258 11452
rect 57012 11398 57014 11450
rect 57194 11398 57196 11450
rect 56950 11396 56956 11398
rect 57012 11396 57036 11398
rect 57092 11396 57116 11398
rect 57172 11396 57196 11398
rect 57252 11396 57258 11398
rect 56950 11387 57258 11396
rect 58532 11144 58584 11150
rect 58532 11086 58584 11092
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 22610 10908 22918 10917
rect 22610 10906 22616 10908
rect 22672 10906 22696 10908
rect 22752 10906 22776 10908
rect 22832 10906 22856 10908
rect 22912 10906 22918 10908
rect 22672 10854 22674 10906
rect 22854 10854 22856 10906
rect 22610 10852 22616 10854
rect 22672 10852 22696 10854
rect 22752 10852 22776 10854
rect 22832 10852 22856 10854
rect 22912 10852 22918 10854
rect 22610 10843 22918 10852
rect 27610 10908 27918 10917
rect 27610 10906 27616 10908
rect 27672 10906 27696 10908
rect 27752 10906 27776 10908
rect 27832 10906 27856 10908
rect 27912 10906 27918 10908
rect 27672 10854 27674 10906
rect 27854 10854 27856 10906
rect 27610 10852 27616 10854
rect 27672 10852 27696 10854
rect 27752 10852 27776 10854
rect 27832 10852 27856 10854
rect 27912 10852 27918 10854
rect 27610 10843 27918 10852
rect 32610 10908 32918 10917
rect 32610 10906 32616 10908
rect 32672 10906 32696 10908
rect 32752 10906 32776 10908
rect 32832 10906 32856 10908
rect 32912 10906 32918 10908
rect 32672 10854 32674 10906
rect 32854 10854 32856 10906
rect 32610 10852 32616 10854
rect 32672 10852 32696 10854
rect 32752 10852 32776 10854
rect 32832 10852 32856 10854
rect 32912 10852 32918 10854
rect 32610 10843 32918 10852
rect 37610 10908 37918 10917
rect 37610 10906 37616 10908
rect 37672 10906 37696 10908
rect 37752 10906 37776 10908
rect 37832 10906 37856 10908
rect 37912 10906 37918 10908
rect 37672 10854 37674 10906
rect 37854 10854 37856 10906
rect 37610 10852 37616 10854
rect 37672 10852 37696 10854
rect 37752 10852 37776 10854
rect 37832 10852 37856 10854
rect 37912 10852 37918 10854
rect 37610 10843 37918 10852
rect 42610 10908 42918 10917
rect 42610 10906 42616 10908
rect 42672 10906 42696 10908
rect 42752 10906 42776 10908
rect 42832 10906 42856 10908
rect 42912 10906 42918 10908
rect 42672 10854 42674 10906
rect 42854 10854 42856 10906
rect 42610 10852 42616 10854
rect 42672 10852 42696 10854
rect 42752 10852 42776 10854
rect 42832 10852 42856 10854
rect 42912 10852 42918 10854
rect 42610 10843 42918 10852
rect 47610 10908 47918 10917
rect 47610 10906 47616 10908
rect 47672 10906 47696 10908
rect 47752 10906 47776 10908
rect 47832 10906 47856 10908
rect 47912 10906 47918 10908
rect 47672 10854 47674 10906
rect 47854 10854 47856 10906
rect 47610 10852 47616 10854
rect 47672 10852 47696 10854
rect 47752 10852 47776 10854
rect 47832 10852 47856 10854
rect 47912 10852 47918 10854
rect 47610 10843 47918 10852
rect 52610 10908 52918 10917
rect 52610 10906 52616 10908
rect 52672 10906 52696 10908
rect 52752 10906 52776 10908
rect 52832 10906 52856 10908
rect 52912 10906 52918 10908
rect 52672 10854 52674 10906
rect 52854 10854 52856 10906
rect 52610 10852 52616 10854
rect 52672 10852 52696 10854
rect 52752 10852 52776 10854
rect 52832 10852 52856 10854
rect 52912 10852 52918 10854
rect 52610 10843 52918 10852
rect 57610 10908 57918 10917
rect 57610 10906 57616 10908
rect 57672 10906 57696 10908
rect 57752 10906 57776 10908
rect 57832 10906 57856 10908
rect 57912 10906 57918 10908
rect 57672 10854 57674 10906
rect 57854 10854 57856 10906
rect 57610 10852 57616 10854
rect 57672 10852 57696 10854
rect 57752 10852 57776 10854
rect 57832 10852 57856 10854
rect 57912 10852 57918 10854
rect 57610 10843 57918 10852
rect 58544 10713 58572 11086
rect 58530 10704 58586 10713
rect 58530 10639 58586 10648
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 21950 10364 22258 10373
rect 21950 10362 21956 10364
rect 22012 10362 22036 10364
rect 22092 10362 22116 10364
rect 22172 10362 22196 10364
rect 22252 10362 22258 10364
rect 22012 10310 22014 10362
rect 22194 10310 22196 10362
rect 21950 10308 21956 10310
rect 22012 10308 22036 10310
rect 22092 10308 22116 10310
rect 22172 10308 22196 10310
rect 22252 10308 22258 10310
rect 21950 10299 22258 10308
rect 26950 10364 27258 10373
rect 26950 10362 26956 10364
rect 27012 10362 27036 10364
rect 27092 10362 27116 10364
rect 27172 10362 27196 10364
rect 27252 10362 27258 10364
rect 27012 10310 27014 10362
rect 27194 10310 27196 10362
rect 26950 10308 26956 10310
rect 27012 10308 27036 10310
rect 27092 10308 27116 10310
rect 27172 10308 27196 10310
rect 27252 10308 27258 10310
rect 26950 10299 27258 10308
rect 31950 10364 32258 10373
rect 31950 10362 31956 10364
rect 32012 10362 32036 10364
rect 32092 10362 32116 10364
rect 32172 10362 32196 10364
rect 32252 10362 32258 10364
rect 32012 10310 32014 10362
rect 32194 10310 32196 10362
rect 31950 10308 31956 10310
rect 32012 10308 32036 10310
rect 32092 10308 32116 10310
rect 32172 10308 32196 10310
rect 32252 10308 32258 10310
rect 31950 10299 32258 10308
rect 36950 10364 37258 10373
rect 36950 10362 36956 10364
rect 37012 10362 37036 10364
rect 37092 10362 37116 10364
rect 37172 10362 37196 10364
rect 37252 10362 37258 10364
rect 37012 10310 37014 10362
rect 37194 10310 37196 10362
rect 36950 10308 36956 10310
rect 37012 10308 37036 10310
rect 37092 10308 37116 10310
rect 37172 10308 37196 10310
rect 37252 10308 37258 10310
rect 36950 10299 37258 10308
rect 41950 10364 42258 10373
rect 41950 10362 41956 10364
rect 42012 10362 42036 10364
rect 42092 10362 42116 10364
rect 42172 10362 42196 10364
rect 42252 10362 42258 10364
rect 42012 10310 42014 10362
rect 42194 10310 42196 10362
rect 41950 10308 41956 10310
rect 42012 10308 42036 10310
rect 42092 10308 42116 10310
rect 42172 10308 42196 10310
rect 42252 10308 42258 10310
rect 41950 10299 42258 10308
rect 46950 10364 47258 10373
rect 46950 10362 46956 10364
rect 47012 10362 47036 10364
rect 47092 10362 47116 10364
rect 47172 10362 47196 10364
rect 47252 10362 47258 10364
rect 47012 10310 47014 10362
rect 47194 10310 47196 10362
rect 46950 10308 46956 10310
rect 47012 10308 47036 10310
rect 47092 10308 47116 10310
rect 47172 10308 47196 10310
rect 47252 10308 47258 10310
rect 46950 10299 47258 10308
rect 51950 10364 52258 10373
rect 51950 10362 51956 10364
rect 52012 10362 52036 10364
rect 52092 10362 52116 10364
rect 52172 10362 52196 10364
rect 52252 10362 52258 10364
rect 52012 10310 52014 10362
rect 52194 10310 52196 10362
rect 51950 10308 51956 10310
rect 52012 10308 52036 10310
rect 52092 10308 52116 10310
rect 52172 10308 52196 10310
rect 52252 10308 52258 10310
rect 51950 10299 52258 10308
rect 56950 10364 57258 10373
rect 56950 10362 56956 10364
rect 57012 10362 57036 10364
rect 57092 10362 57116 10364
rect 57172 10362 57196 10364
rect 57252 10362 57258 10364
rect 57012 10310 57014 10362
rect 57194 10310 57196 10362
rect 56950 10308 56956 10310
rect 57012 10308 57036 10310
rect 57092 10308 57116 10310
rect 57172 10308 57196 10310
rect 57252 10308 57258 10310
rect 56950 10299 57258 10308
rect 58532 10056 58584 10062
rect 58532 9998 58584 10004
rect 58544 9897 58572 9998
rect 58530 9888 58586 9897
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 22610 9820 22918 9829
rect 22610 9818 22616 9820
rect 22672 9818 22696 9820
rect 22752 9818 22776 9820
rect 22832 9818 22856 9820
rect 22912 9818 22918 9820
rect 22672 9766 22674 9818
rect 22854 9766 22856 9818
rect 22610 9764 22616 9766
rect 22672 9764 22696 9766
rect 22752 9764 22776 9766
rect 22832 9764 22856 9766
rect 22912 9764 22918 9766
rect 22610 9755 22918 9764
rect 27610 9820 27918 9829
rect 27610 9818 27616 9820
rect 27672 9818 27696 9820
rect 27752 9818 27776 9820
rect 27832 9818 27856 9820
rect 27912 9818 27918 9820
rect 27672 9766 27674 9818
rect 27854 9766 27856 9818
rect 27610 9764 27616 9766
rect 27672 9764 27696 9766
rect 27752 9764 27776 9766
rect 27832 9764 27856 9766
rect 27912 9764 27918 9766
rect 27610 9755 27918 9764
rect 32610 9820 32918 9829
rect 32610 9818 32616 9820
rect 32672 9818 32696 9820
rect 32752 9818 32776 9820
rect 32832 9818 32856 9820
rect 32912 9818 32918 9820
rect 32672 9766 32674 9818
rect 32854 9766 32856 9818
rect 32610 9764 32616 9766
rect 32672 9764 32696 9766
rect 32752 9764 32776 9766
rect 32832 9764 32856 9766
rect 32912 9764 32918 9766
rect 32610 9755 32918 9764
rect 37610 9820 37918 9829
rect 37610 9818 37616 9820
rect 37672 9818 37696 9820
rect 37752 9818 37776 9820
rect 37832 9818 37856 9820
rect 37912 9818 37918 9820
rect 37672 9766 37674 9818
rect 37854 9766 37856 9818
rect 37610 9764 37616 9766
rect 37672 9764 37696 9766
rect 37752 9764 37776 9766
rect 37832 9764 37856 9766
rect 37912 9764 37918 9766
rect 37610 9755 37918 9764
rect 42610 9820 42918 9829
rect 42610 9818 42616 9820
rect 42672 9818 42696 9820
rect 42752 9818 42776 9820
rect 42832 9818 42856 9820
rect 42912 9818 42918 9820
rect 42672 9766 42674 9818
rect 42854 9766 42856 9818
rect 42610 9764 42616 9766
rect 42672 9764 42696 9766
rect 42752 9764 42776 9766
rect 42832 9764 42856 9766
rect 42912 9764 42918 9766
rect 42610 9755 42918 9764
rect 47610 9820 47918 9829
rect 47610 9818 47616 9820
rect 47672 9818 47696 9820
rect 47752 9818 47776 9820
rect 47832 9818 47856 9820
rect 47912 9818 47918 9820
rect 47672 9766 47674 9818
rect 47854 9766 47856 9818
rect 47610 9764 47616 9766
rect 47672 9764 47696 9766
rect 47752 9764 47776 9766
rect 47832 9764 47856 9766
rect 47912 9764 47918 9766
rect 47610 9755 47918 9764
rect 52610 9820 52918 9829
rect 52610 9818 52616 9820
rect 52672 9818 52696 9820
rect 52752 9818 52776 9820
rect 52832 9818 52856 9820
rect 52912 9818 52918 9820
rect 52672 9766 52674 9818
rect 52854 9766 52856 9818
rect 52610 9764 52616 9766
rect 52672 9764 52696 9766
rect 52752 9764 52776 9766
rect 52832 9764 52856 9766
rect 52912 9764 52918 9766
rect 52610 9755 52918 9764
rect 57610 9820 57918 9829
rect 58530 9823 58586 9832
rect 57610 9818 57616 9820
rect 57672 9818 57696 9820
rect 57752 9818 57776 9820
rect 57832 9818 57856 9820
rect 57912 9818 57918 9820
rect 57672 9766 57674 9818
rect 57854 9766 57856 9818
rect 57610 9764 57616 9766
rect 57672 9764 57696 9766
rect 57752 9764 57776 9766
rect 57832 9764 57856 9766
rect 57912 9764 57918 9766
rect 57610 9755 57918 9764
rect 58532 9376 58584 9382
rect 58532 9318 58584 9324
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 21950 9276 22258 9285
rect 21950 9274 21956 9276
rect 22012 9274 22036 9276
rect 22092 9274 22116 9276
rect 22172 9274 22196 9276
rect 22252 9274 22258 9276
rect 22012 9222 22014 9274
rect 22194 9222 22196 9274
rect 21950 9220 21956 9222
rect 22012 9220 22036 9222
rect 22092 9220 22116 9222
rect 22172 9220 22196 9222
rect 22252 9220 22258 9222
rect 21950 9211 22258 9220
rect 26950 9276 27258 9285
rect 26950 9274 26956 9276
rect 27012 9274 27036 9276
rect 27092 9274 27116 9276
rect 27172 9274 27196 9276
rect 27252 9274 27258 9276
rect 27012 9222 27014 9274
rect 27194 9222 27196 9274
rect 26950 9220 26956 9222
rect 27012 9220 27036 9222
rect 27092 9220 27116 9222
rect 27172 9220 27196 9222
rect 27252 9220 27258 9222
rect 26950 9211 27258 9220
rect 31950 9276 32258 9285
rect 31950 9274 31956 9276
rect 32012 9274 32036 9276
rect 32092 9274 32116 9276
rect 32172 9274 32196 9276
rect 32252 9274 32258 9276
rect 32012 9222 32014 9274
rect 32194 9222 32196 9274
rect 31950 9220 31956 9222
rect 32012 9220 32036 9222
rect 32092 9220 32116 9222
rect 32172 9220 32196 9222
rect 32252 9220 32258 9222
rect 31950 9211 32258 9220
rect 36950 9276 37258 9285
rect 36950 9274 36956 9276
rect 37012 9274 37036 9276
rect 37092 9274 37116 9276
rect 37172 9274 37196 9276
rect 37252 9274 37258 9276
rect 37012 9222 37014 9274
rect 37194 9222 37196 9274
rect 36950 9220 36956 9222
rect 37012 9220 37036 9222
rect 37092 9220 37116 9222
rect 37172 9220 37196 9222
rect 37252 9220 37258 9222
rect 36950 9211 37258 9220
rect 41950 9276 42258 9285
rect 41950 9274 41956 9276
rect 42012 9274 42036 9276
rect 42092 9274 42116 9276
rect 42172 9274 42196 9276
rect 42252 9274 42258 9276
rect 42012 9222 42014 9274
rect 42194 9222 42196 9274
rect 41950 9220 41956 9222
rect 42012 9220 42036 9222
rect 42092 9220 42116 9222
rect 42172 9220 42196 9222
rect 42252 9220 42258 9222
rect 41950 9211 42258 9220
rect 46950 9276 47258 9285
rect 46950 9274 46956 9276
rect 47012 9274 47036 9276
rect 47092 9274 47116 9276
rect 47172 9274 47196 9276
rect 47252 9274 47258 9276
rect 47012 9222 47014 9274
rect 47194 9222 47196 9274
rect 46950 9220 46956 9222
rect 47012 9220 47036 9222
rect 47092 9220 47116 9222
rect 47172 9220 47196 9222
rect 47252 9220 47258 9222
rect 46950 9211 47258 9220
rect 51950 9276 52258 9285
rect 51950 9274 51956 9276
rect 52012 9274 52036 9276
rect 52092 9274 52116 9276
rect 52172 9274 52196 9276
rect 52252 9274 52258 9276
rect 52012 9222 52014 9274
rect 52194 9222 52196 9274
rect 51950 9220 51956 9222
rect 52012 9220 52036 9222
rect 52092 9220 52116 9222
rect 52172 9220 52196 9222
rect 52252 9220 52258 9222
rect 51950 9211 52258 9220
rect 56950 9276 57258 9285
rect 56950 9274 56956 9276
rect 57012 9274 57036 9276
rect 57092 9274 57116 9276
rect 57172 9274 57196 9276
rect 57252 9274 57258 9276
rect 57012 9222 57014 9274
rect 57194 9222 57196 9274
rect 56950 9220 56956 9222
rect 57012 9220 57036 9222
rect 57092 9220 57116 9222
rect 57172 9220 57196 9222
rect 57252 9220 57258 9222
rect 56950 9211 57258 9220
rect 58544 9081 58572 9318
rect 58530 9072 58586 9081
rect 58530 9007 58586 9016
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 22610 8732 22918 8741
rect 22610 8730 22616 8732
rect 22672 8730 22696 8732
rect 22752 8730 22776 8732
rect 22832 8730 22856 8732
rect 22912 8730 22918 8732
rect 22672 8678 22674 8730
rect 22854 8678 22856 8730
rect 22610 8676 22616 8678
rect 22672 8676 22696 8678
rect 22752 8676 22776 8678
rect 22832 8676 22856 8678
rect 22912 8676 22918 8678
rect 22610 8667 22918 8676
rect 27610 8732 27918 8741
rect 27610 8730 27616 8732
rect 27672 8730 27696 8732
rect 27752 8730 27776 8732
rect 27832 8730 27856 8732
rect 27912 8730 27918 8732
rect 27672 8678 27674 8730
rect 27854 8678 27856 8730
rect 27610 8676 27616 8678
rect 27672 8676 27696 8678
rect 27752 8676 27776 8678
rect 27832 8676 27856 8678
rect 27912 8676 27918 8678
rect 27610 8667 27918 8676
rect 32610 8732 32918 8741
rect 32610 8730 32616 8732
rect 32672 8730 32696 8732
rect 32752 8730 32776 8732
rect 32832 8730 32856 8732
rect 32912 8730 32918 8732
rect 32672 8678 32674 8730
rect 32854 8678 32856 8730
rect 32610 8676 32616 8678
rect 32672 8676 32696 8678
rect 32752 8676 32776 8678
rect 32832 8676 32856 8678
rect 32912 8676 32918 8678
rect 32610 8667 32918 8676
rect 37610 8732 37918 8741
rect 37610 8730 37616 8732
rect 37672 8730 37696 8732
rect 37752 8730 37776 8732
rect 37832 8730 37856 8732
rect 37912 8730 37918 8732
rect 37672 8678 37674 8730
rect 37854 8678 37856 8730
rect 37610 8676 37616 8678
rect 37672 8676 37696 8678
rect 37752 8676 37776 8678
rect 37832 8676 37856 8678
rect 37912 8676 37918 8678
rect 37610 8667 37918 8676
rect 42610 8732 42918 8741
rect 42610 8730 42616 8732
rect 42672 8730 42696 8732
rect 42752 8730 42776 8732
rect 42832 8730 42856 8732
rect 42912 8730 42918 8732
rect 42672 8678 42674 8730
rect 42854 8678 42856 8730
rect 42610 8676 42616 8678
rect 42672 8676 42696 8678
rect 42752 8676 42776 8678
rect 42832 8676 42856 8678
rect 42912 8676 42918 8678
rect 42610 8667 42918 8676
rect 47610 8732 47918 8741
rect 47610 8730 47616 8732
rect 47672 8730 47696 8732
rect 47752 8730 47776 8732
rect 47832 8730 47856 8732
rect 47912 8730 47918 8732
rect 47672 8678 47674 8730
rect 47854 8678 47856 8730
rect 47610 8676 47616 8678
rect 47672 8676 47696 8678
rect 47752 8676 47776 8678
rect 47832 8676 47856 8678
rect 47912 8676 47918 8678
rect 47610 8667 47918 8676
rect 52610 8732 52918 8741
rect 52610 8730 52616 8732
rect 52672 8730 52696 8732
rect 52752 8730 52776 8732
rect 52832 8730 52856 8732
rect 52912 8730 52918 8732
rect 52672 8678 52674 8730
rect 52854 8678 52856 8730
rect 52610 8676 52616 8678
rect 52672 8676 52696 8678
rect 52752 8676 52776 8678
rect 52832 8676 52856 8678
rect 52912 8676 52918 8678
rect 52610 8667 52918 8676
rect 57610 8732 57918 8741
rect 57610 8730 57616 8732
rect 57672 8730 57696 8732
rect 57752 8730 57776 8732
rect 57832 8730 57856 8732
rect 57912 8730 57918 8732
rect 57672 8678 57674 8730
rect 57854 8678 57856 8730
rect 57610 8676 57616 8678
rect 57672 8676 57696 8678
rect 57752 8676 57776 8678
rect 57832 8676 57856 8678
rect 57912 8676 57918 8678
rect 57610 8667 57918 8676
rect 58532 8356 58584 8362
rect 58532 8298 58584 8304
rect 58544 8265 58572 8298
rect 58530 8256 58586 8265
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 21950 8188 22258 8197
rect 21950 8186 21956 8188
rect 22012 8186 22036 8188
rect 22092 8186 22116 8188
rect 22172 8186 22196 8188
rect 22252 8186 22258 8188
rect 22012 8134 22014 8186
rect 22194 8134 22196 8186
rect 21950 8132 21956 8134
rect 22012 8132 22036 8134
rect 22092 8132 22116 8134
rect 22172 8132 22196 8134
rect 22252 8132 22258 8134
rect 21950 8123 22258 8132
rect 26950 8188 27258 8197
rect 26950 8186 26956 8188
rect 27012 8186 27036 8188
rect 27092 8186 27116 8188
rect 27172 8186 27196 8188
rect 27252 8186 27258 8188
rect 27012 8134 27014 8186
rect 27194 8134 27196 8186
rect 26950 8132 26956 8134
rect 27012 8132 27036 8134
rect 27092 8132 27116 8134
rect 27172 8132 27196 8134
rect 27252 8132 27258 8134
rect 26950 8123 27258 8132
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 36950 8188 37258 8197
rect 36950 8186 36956 8188
rect 37012 8186 37036 8188
rect 37092 8186 37116 8188
rect 37172 8186 37196 8188
rect 37252 8186 37258 8188
rect 37012 8134 37014 8186
rect 37194 8134 37196 8186
rect 36950 8132 36956 8134
rect 37012 8132 37036 8134
rect 37092 8132 37116 8134
rect 37172 8132 37196 8134
rect 37252 8132 37258 8134
rect 36950 8123 37258 8132
rect 41950 8188 42258 8197
rect 41950 8186 41956 8188
rect 42012 8186 42036 8188
rect 42092 8186 42116 8188
rect 42172 8186 42196 8188
rect 42252 8186 42258 8188
rect 42012 8134 42014 8186
rect 42194 8134 42196 8186
rect 41950 8132 41956 8134
rect 42012 8132 42036 8134
rect 42092 8132 42116 8134
rect 42172 8132 42196 8134
rect 42252 8132 42258 8134
rect 41950 8123 42258 8132
rect 46950 8188 47258 8197
rect 46950 8186 46956 8188
rect 47012 8186 47036 8188
rect 47092 8186 47116 8188
rect 47172 8186 47196 8188
rect 47252 8186 47258 8188
rect 47012 8134 47014 8186
rect 47194 8134 47196 8186
rect 46950 8132 46956 8134
rect 47012 8132 47036 8134
rect 47092 8132 47116 8134
rect 47172 8132 47196 8134
rect 47252 8132 47258 8134
rect 46950 8123 47258 8132
rect 51950 8188 52258 8197
rect 51950 8186 51956 8188
rect 52012 8186 52036 8188
rect 52092 8186 52116 8188
rect 52172 8186 52196 8188
rect 52252 8186 52258 8188
rect 52012 8134 52014 8186
rect 52194 8134 52196 8186
rect 51950 8132 51956 8134
rect 52012 8132 52036 8134
rect 52092 8132 52116 8134
rect 52172 8132 52196 8134
rect 52252 8132 52258 8134
rect 51950 8123 52258 8132
rect 56950 8188 57258 8197
rect 58530 8191 58586 8200
rect 56950 8186 56956 8188
rect 57012 8186 57036 8188
rect 57092 8186 57116 8188
rect 57172 8186 57196 8188
rect 57252 8186 57258 8188
rect 57012 8134 57014 8186
rect 57194 8134 57196 8186
rect 56950 8132 56956 8134
rect 57012 8132 57036 8134
rect 57092 8132 57116 8134
rect 57172 8132 57196 8134
rect 57252 8132 57258 8134
rect 56950 8123 57258 8132
rect 58532 7880 58584 7886
rect 58532 7822 58584 7828
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 22610 7644 22918 7653
rect 22610 7642 22616 7644
rect 22672 7642 22696 7644
rect 22752 7642 22776 7644
rect 22832 7642 22856 7644
rect 22912 7642 22918 7644
rect 22672 7590 22674 7642
rect 22854 7590 22856 7642
rect 22610 7588 22616 7590
rect 22672 7588 22696 7590
rect 22752 7588 22776 7590
rect 22832 7588 22856 7590
rect 22912 7588 22918 7590
rect 22610 7579 22918 7588
rect 27610 7644 27918 7653
rect 27610 7642 27616 7644
rect 27672 7642 27696 7644
rect 27752 7642 27776 7644
rect 27832 7642 27856 7644
rect 27912 7642 27918 7644
rect 27672 7590 27674 7642
rect 27854 7590 27856 7642
rect 27610 7588 27616 7590
rect 27672 7588 27696 7590
rect 27752 7588 27776 7590
rect 27832 7588 27856 7590
rect 27912 7588 27918 7590
rect 27610 7579 27918 7588
rect 32610 7644 32918 7653
rect 32610 7642 32616 7644
rect 32672 7642 32696 7644
rect 32752 7642 32776 7644
rect 32832 7642 32856 7644
rect 32912 7642 32918 7644
rect 32672 7590 32674 7642
rect 32854 7590 32856 7642
rect 32610 7588 32616 7590
rect 32672 7588 32696 7590
rect 32752 7588 32776 7590
rect 32832 7588 32856 7590
rect 32912 7588 32918 7590
rect 32610 7579 32918 7588
rect 37610 7644 37918 7653
rect 37610 7642 37616 7644
rect 37672 7642 37696 7644
rect 37752 7642 37776 7644
rect 37832 7642 37856 7644
rect 37912 7642 37918 7644
rect 37672 7590 37674 7642
rect 37854 7590 37856 7642
rect 37610 7588 37616 7590
rect 37672 7588 37696 7590
rect 37752 7588 37776 7590
rect 37832 7588 37856 7590
rect 37912 7588 37918 7590
rect 37610 7579 37918 7588
rect 42610 7644 42918 7653
rect 42610 7642 42616 7644
rect 42672 7642 42696 7644
rect 42752 7642 42776 7644
rect 42832 7642 42856 7644
rect 42912 7642 42918 7644
rect 42672 7590 42674 7642
rect 42854 7590 42856 7642
rect 42610 7588 42616 7590
rect 42672 7588 42696 7590
rect 42752 7588 42776 7590
rect 42832 7588 42856 7590
rect 42912 7588 42918 7590
rect 42610 7579 42918 7588
rect 47610 7644 47918 7653
rect 47610 7642 47616 7644
rect 47672 7642 47696 7644
rect 47752 7642 47776 7644
rect 47832 7642 47856 7644
rect 47912 7642 47918 7644
rect 47672 7590 47674 7642
rect 47854 7590 47856 7642
rect 47610 7588 47616 7590
rect 47672 7588 47696 7590
rect 47752 7588 47776 7590
rect 47832 7588 47856 7590
rect 47912 7588 47918 7590
rect 47610 7579 47918 7588
rect 52610 7644 52918 7653
rect 52610 7642 52616 7644
rect 52672 7642 52696 7644
rect 52752 7642 52776 7644
rect 52832 7642 52856 7644
rect 52912 7642 52918 7644
rect 52672 7590 52674 7642
rect 52854 7590 52856 7642
rect 52610 7588 52616 7590
rect 52672 7588 52696 7590
rect 52752 7588 52776 7590
rect 52832 7588 52856 7590
rect 52912 7588 52918 7590
rect 52610 7579 52918 7588
rect 57610 7644 57918 7653
rect 57610 7642 57616 7644
rect 57672 7642 57696 7644
rect 57752 7642 57776 7644
rect 57832 7642 57856 7644
rect 57912 7642 57918 7644
rect 57672 7590 57674 7642
rect 57854 7590 57856 7642
rect 57610 7588 57616 7590
rect 57672 7588 57696 7590
rect 57752 7588 57776 7590
rect 57832 7588 57856 7590
rect 57912 7588 57918 7590
rect 57610 7579 57918 7588
rect 58544 7449 58572 7822
rect 58530 7440 58586 7449
rect 58530 7375 58586 7384
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 21950 7100 22258 7109
rect 21950 7098 21956 7100
rect 22012 7098 22036 7100
rect 22092 7098 22116 7100
rect 22172 7098 22196 7100
rect 22252 7098 22258 7100
rect 22012 7046 22014 7098
rect 22194 7046 22196 7098
rect 21950 7044 21956 7046
rect 22012 7044 22036 7046
rect 22092 7044 22116 7046
rect 22172 7044 22196 7046
rect 22252 7044 22258 7046
rect 21950 7035 22258 7044
rect 26950 7100 27258 7109
rect 26950 7098 26956 7100
rect 27012 7098 27036 7100
rect 27092 7098 27116 7100
rect 27172 7098 27196 7100
rect 27252 7098 27258 7100
rect 27012 7046 27014 7098
rect 27194 7046 27196 7098
rect 26950 7044 26956 7046
rect 27012 7044 27036 7046
rect 27092 7044 27116 7046
rect 27172 7044 27196 7046
rect 27252 7044 27258 7046
rect 26950 7035 27258 7044
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 36950 7100 37258 7109
rect 36950 7098 36956 7100
rect 37012 7098 37036 7100
rect 37092 7098 37116 7100
rect 37172 7098 37196 7100
rect 37252 7098 37258 7100
rect 37012 7046 37014 7098
rect 37194 7046 37196 7098
rect 36950 7044 36956 7046
rect 37012 7044 37036 7046
rect 37092 7044 37116 7046
rect 37172 7044 37196 7046
rect 37252 7044 37258 7046
rect 36950 7035 37258 7044
rect 41950 7100 42258 7109
rect 41950 7098 41956 7100
rect 42012 7098 42036 7100
rect 42092 7098 42116 7100
rect 42172 7098 42196 7100
rect 42252 7098 42258 7100
rect 42012 7046 42014 7098
rect 42194 7046 42196 7098
rect 41950 7044 41956 7046
rect 42012 7044 42036 7046
rect 42092 7044 42116 7046
rect 42172 7044 42196 7046
rect 42252 7044 42258 7046
rect 41950 7035 42258 7044
rect 46950 7100 47258 7109
rect 46950 7098 46956 7100
rect 47012 7098 47036 7100
rect 47092 7098 47116 7100
rect 47172 7098 47196 7100
rect 47252 7098 47258 7100
rect 47012 7046 47014 7098
rect 47194 7046 47196 7098
rect 46950 7044 46956 7046
rect 47012 7044 47036 7046
rect 47092 7044 47116 7046
rect 47172 7044 47196 7046
rect 47252 7044 47258 7046
rect 46950 7035 47258 7044
rect 51950 7100 52258 7109
rect 51950 7098 51956 7100
rect 52012 7098 52036 7100
rect 52092 7098 52116 7100
rect 52172 7098 52196 7100
rect 52252 7098 52258 7100
rect 52012 7046 52014 7098
rect 52194 7046 52196 7098
rect 51950 7044 51956 7046
rect 52012 7044 52036 7046
rect 52092 7044 52116 7046
rect 52172 7044 52196 7046
rect 52252 7044 52258 7046
rect 51950 7035 52258 7044
rect 56950 7100 57258 7109
rect 56950 7098 56956 7100
rect 57012 7098 57036 7100
rect 57092 7098 57116 7100
rect 57172 7098 57196 7100
rect 57252 7098 57258 7100
rect 57012 7046 57014 7098
rect 57194 7046 57196 7098
rect 56950 7044 56956 7046
rect 57012 7044 57036 7046
rect 57092 7044 57116 7046
rect 57172 7044 57196 7046
rect 57252 7044 57258 7046
rect 56950 7035 57258 7044
rect 58532 6792 58584 6798
rect 58532 6734 58584 6740
rect 58544 6633 58572 6734
rect 58530 6624 58586 6633
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 22610 6556 22918 6565
rect 22610 6554 22616 6556
rect 22672 6554 22696 6556
rect 22752 6554 22776 6556
rect 22832 6554 22856 6556
rect 22912 6554 22918 6556
rect 22672 6502 22674 6554
rect 22854 6502 22856 6554
rect 22610 6500 22616 6502
rect 22672 6500 22696 6502
rect 22752 6500 22776 6502
rect 22832 6500 22856 6502
rect 22912 6500 22918 6502
rect 22610 6491 22918 6500
rect 27610 6556 27918 6565
rect 27610 6554 27616 6556
rect 27672 6554 27696 6556
rect 27752 6554 27776 6556
rect 27832 6554 27856 6556
rect 27912 6554 27918 6556
rect 27672 6502 27674 6554
rect 27854 6502 27856 6554
rect 27610 6500 27616 6502
rect 27672 6500 27696 6502
rect 27752 6500 27776 6502
rect 27832 6500 27856 6502
rect 27912 6500 27918 6502
rect 27610 6491 27918 6500
rect 32610 6556 32918 6565
rect 32610 6554 32616 6556
rect 32672 6554 32696 6556
rect 32752 6554 32776 6556
rect 32832 6554 32856 6556
rect 32912 6554 32918 6556
rect 32672 6502 32674 6554
rect 32854 6502 32856 6554
rect 32610 6500 32616 6502
rect 32672 6500 32696 6502
rect 32752 6500 32776 6502
rect 32832 6500 32856 6502
rect 32912 6500 32918 6502
rect 32610 6491 32918 6500
rect 37610 6556 37918 6565
rect 37610 6554 37616 6556
rect 37672 6554 37696 6556
rect 37752 6554 37776 6556
rect 37832 6554 37856 6556
rect 37912 6554 37918 6556
rect 37672 6502 37674 6554
rect 37854 6502 37856 6554
rect 37610 6500 37616 6502
rect 37672 6500 37696 6502
rect 37752 6500 37776 6502
rect 37832 6500 37856 6502
rect 37912 6500 37918 6502
rect 37610 6491 37918 6500
rect 42610 6556 42918 6565
rect 42610 6554 42616 6556
rect 42672 6554 42696 6556
rect 42752 6554 42776 6556
rect 42832 6554 42856 6556
rect 42912 6554 42918 6556
rect 42672 6502 42674 6554
rect 42854 6502 42856 6554
rect 42610 6500 42616 6502
rect 42672 6500 42696 6502
rect 42752 6500 42776 6502
rect 42832 6500 42856 6502
rect 42912 6500 42918 6502
rect 42610 6491 42918 6500
rect 47610 6556 47918 6565
rect 47610 6554 47616 6556
rect 47672 6554 47696 6556
rect 47752 6554 47776 6556
rect 47832 6554 47856 6556
rect 47912 6554 47918 6556
rect 47672 6502 47674 6554
rect 47854 6502 47856 6554
rect 47610 6500 47616 6502
rect 47672 6500 47696 6502
rect 47752 6500 47776 6502
rect 47832 6500 47856 6502
rect 47912 6500 47918 6502
rect 47610 6491 47918 6500
rect 52610 6556 52918 6565
rect 52610 6554 52616 6556
rect 52672 6554 52696 6556
rect 52752 6554 52776 6556
rect 52832 6554 52856 6556
rect 52912 6554 52918 6556
rect 52672 6502 52674 6554
rect 52854 6502 52856 6554
rect 52610 6500 52616 6502
rect 52672 6500 52696 6502
rect 52752 6500 52776 6502
rect 52832 6500 52856 6502
rect 52912 6500 52918 6502
rect 52610 6491 52918 6500
rect 57610 6556 57918 6565
rect 58530 6559 58586 6568
rect 57610 6554 57616 6556
rect 57672 6554 57696 6556
rect 57752 6554 57776 6556
rect 57832 6554 57856 6556
rect 57912 6554 57918 6556
rect 57672 6502 57674 6554
rect 57854 6502 57856 6554
rect 57610 6500 57616 6502
rect 57672 6500 57696 6502
rect 57752 6500 57776 6502
rect 57832 6500 57856 6502
rect 57912 6500 57918 6502
rect 57610 6491 57918 6500
rect 58532 6112 58584 6118
rect 58532 6054 58584 6060
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 21950 6012 22258 6021
rect 21950 6010 21956 6012
rect 22012 6010 22036 6012
rect 22092 6010 22116 6012
rect 22172 6010 22196 6012
rect 22252 6010 22258 6012
rect 22012 5958 22014 6010
rect 22194 5958 22196 6010
rect 21950 5956 21956 5958
rect 22012 5956 22036 5958
rect 22092 5956 22116 5958
rect 22172 5956 22196 5958
rect 22252 5956 22258 5958
rect 21950 5947 22258 5956
rect 26950 6012 27258 6021
rect 26950 6010 26956 6012
rect 27012 6010 27036 6012
rect 27092 6010 27116 6012
rect 27172 6010 27196 6012
rect 27252 6010 27258 6012
rect 27012 5958 27014 6010
rect 27194 5958 27196 6010
rect 26950 5956 26956 5958
rect 27012 5956 27036 5958
rect 27092 5956 27116 5958
rect 27172 5956 27196 5958
rect 27252 5956 27258 5958
rect 26950 5947 27258 5956
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 36950 6012 37258 6021
rect 36950 6010 36956 6012
rect 37012 6010 37036 6012
rect 37092 6010 37116 6012
rect 37172 6010 37196 6012
rect 37252 6010 37258 6012
rect 37012 5958 37014 6010
rect 37194 5958 37196 6010
rect 36950 5956 36956 5958
rect 37012 5956 37036 5958
rect 37092 5956 37116 5958
rect 37172 5956 37196 5958
rect 37252 5956 37258 5958
rect 36950 5947 37258 5956
rect 41950 6012 42258 6021
rect 41950 6010 41956 6012
rect 42012 6010 42036 6012
rect 42092 6010 42116 6012
rect 42172 6010 42196 6012
rect 42252 6010 42258 6012
rect 42012 5958 42014 6010
rect 42194 5958 42196 6010
rect 41950 5956 41956 5958
rect 42012 5956 42036 5958
rect 42092 5956 42116 5958
rect 42172 5956 42196 5958
rect 42252 5956 42258 5958
rect 41950 5947 42258 5956
rect 46950 6012 47258 6021
rect 46950 6010 46956 6012
rect 47012 6010 47036 6012
rect 47092 6010 47116 6012
rect 47172 6010 47196 6012
rect 47252 6010 47258 6012
rect 47012 5958 47014 6010
rect 47194 5958 47196 6010
rect 46950 5956 46956 5958
rect 47012 5956 47036 5958
rect 47092 5956 47116 5958
rect 47172 5956 47196 5958
rect 47252 5956 47258 5958
rect 46950 5947 47258 5956
rect 51950 6012 52258 6021
rect 51950 6010 51956 6012
rect 52012 6010 52036 6012
rect 52092 6010 52116 6012
rect 52172 6010 52196 6012
rect 52252 6010 52258 6012
rect 52012 5958 52014 6010
rect 52194 5958 52196 6010
rect 51950 5956 51956 5958
rect 52012 5956 52036 5958
rect 52092 5956 52116 5958
rect 52172 5956 52196 5958
rect 52252 5956 52258 5958
rect 51950 5947 52258 5956
rect 56950 6012 57258 6021
rect 56950 6010 56956 6012
rect 57012 6010 57036 6012
rect 57092 6010 57116 6012
rect 57172 6010 57196 6012
rect 57252 6010 57258 6012
rect 57012 5958 57014 6010
rect 57194 5958 57196 6010
rect 56950 5956 56956 5958
rect 57012 5956 57036 5958
rect 57092 5956 57116 5958
rect 57172 5956 57196 5958
rect 57252 5956 57258 5958
rect 56950 5947 57258 5956
rect 58544 5817 58572 6054
rect 58530 5808 58586 5817
rect 58530 5743 58586 5752
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 22610 5468 22918 5477
rect 22610 5466 22616 5468
rect 22672 5466 22696 5468
rect 22752 5466 22776 5468
rect 22832 5466 22856 5468
rect 22912 5466 22918 5468
rect 22672 5414 22674 5466
rect 22854 5414 22856 5466
rect 22610 5412 22616 5414
rect 22672 5412 22696 5414
rect 22752 5412 22776 5414
rect 22832 5412 22856 5414
rect 22912 5412 22918 5414
rect 22610 5403 22918 5412
rect 27610 5468 27918 5477
rect 27610 5466 27616 5468
rect 27672 5466 27696 5468
rect 27752 5466 27776 5468
rect 27832 5466 27856 5468
rect 27912 5466 27918 5468
rect 27672 5414 27674 5466
rect 27854 5414 27856 5466
rect 27610 5412 27616 5414
rect 27672 5412 27696 5414
rect 27752 5412 27776 5414
rect 27832 5412 27856 5414
rect 27912 5412 27918 5414
rect 27610 5403 27918 5412
rect 32610 5468 32918 5477
rect 32610 5466 32616 5468
rect 32672 5466 32696 5468
rect 32752 5466 32776 5468
rect 32832 5466 32856 5468
rect 32912 5466 32918 5468
rect 32672 5414 32674 5466
rect 32854 5414 32856 5466
rect 32610 5412 32616 5414
rect 32672 5412 32696 5414
rect 32752 5412 32776 5414
rect 32832 5412 32856 5414
rect 32912 5412 32918 5414
rect 32610 5403 32918 5412
rect 37610 5468 37918 5477
rect 37610 5466 37616 5468
rect 37672 5466 37696 5468
rect 37752 5466 37776 5468
rect 37832 5466 37856 5468
rect 37912 5466 37918 5468
rect 37672 5414 37674 5466
rect 37854 5414 37856 5466
rect 37610 5412 37616 5414
rect 37672 5412 37696 5414
rect 37752 5412 37776 5414
rect 37832 5412 37856 5414
rect 37912 5412 37918 5414
rect 37610 5403 37918 5412
rect 42610 5468 42918 5477
rect 42610 5466 42616 5468
rect 42672 5466 42696 5468
rect 42752 5466 42776 5468
rect 42832 5466 42856 5468
rect 42912 5466 42918 5468
rect 42672 5414 42674 5466
rect 42854 5414 42856 5466
rect 42610 5412 42616 5414
rect 42672 5412 42696 5414
rect 42752 5412 42776 5414
rect 42832 5412 42856 5414
rect 42912 5412 42918 5414
rect 42610 5403 42918 5412
rect 47610 5468 47918 5477
rect 47610 5466 47616 5468
rect 47672 5466 47696 5468
rect 47752 5466 47776 5468
rect 47832 5466 47856 5468
rect 47912 5466 47918 5468
rect 47672 5414 47674 5466
rect 47854 5414 47856 5466
rect 47610 5412 47616 5414
rect 47672 5412 47696 5414
rect 47752 5412 47776 5414
rect 47832 5412 47856 5414
rect 47912 5412 47918 5414
rect 47610 5403 47918 5412
rect 52610 5468 52918 5477
rect 52610 5466 52616 5468
rect 52672 5466 52696 5468
rect 52752 5466 52776 5468
rect 52832 5466 52856 5468
rect 52912 5466 52918 5468
rect 52672 5414 52674 5466
rect 52854 5414 52856 5466
rect 52610 5412 52616 5414
rect 52672 5412 52696 5414
rect 52752 5412 52776 5414
rect 52832 5412 52856 5414
rect 52912 5412 52918 5414
rect 52610 5403 52918 5412
rect 57610 5468 57918 5477
rect 57610 5466 57616 5468
rect 57672 5466 57696 5468
rect 57752 5466 57776 5468
rect 57832 5466 57856 5468
rect 57912 5466 57918 5468
rect 57672 5414 57674 5466
rect 57854 5414 57856 5466
rect 57610 5412 57616 5414
rect 57672 5412 57696 5414
rect 57752 5412 57776 5414
rect 57832 5412 57856 5414
rect 57912 5412 57918 5414
rect 57610 5403 57918 5412
rect 58532 5024 58584 5030
rect 58530 4992 58532 5001
rect 58584 4992 58586 5001
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 21950 4924 22258 4933
rect 21950 4922 21956 4924
rect 22012 4922 22036 4924
rect 22092 4922 22116 4924
rect 22172 4922 22196 4924
rect 22252 4922 22258 4924
rect 22012 4870 22014 4922
rect 22194 4870 22196 4922
rect 21950 4868 21956 4870
rect 22012 4868 22036 4870
rect 22092 4868 22116 4870
rect 22172 4868 22196 4870
rect 22252 4868 22258 4870
rect 21950 4859 22258 4868
rect 26950 4924 27258 4933
rect 26950 4922 26956 4924
rect 27012 4922 27036 4924
rect 27092 4922 27116 4924
rect 27172 4922 27196 4924
rect 27252 4922 27258 4924
rect 27012 4870 27014 4922
rect 27194 4870 27196 4922
rect 26950 4868 26956 4870
rect 27012 4868 27036 4870
rect 27092 4868 27116 4870
rect 27172 4868 27196 4870
rect 27252 4868 27258 4870
rect 26950 4859 27258 4868
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 36950 4924 37258 4933
rect 36950 4922 36956 4924
rect 37012 4922 37036 4924
rect 37092 4922 37116 4924
rect 37172 4922 37196 4924
rect 37252 4922 37258 4924
rect 37012 4870 37014 4922
rect 37194 4870 37196 4922
rect 36950 4868 36956 4870
rect 37012 4868 37036 4870
rect 37092 4868 37116 4870
rect 37172 4868 37196 4870
rect 37252 4868 37258 4870
rect 36950 4859 37258 4868
rect 41950 4924 42258 4933
rect 41950 4922 41956 4924
rect 42012 4922 42036 4924
rect 42092 4922 42116 4924
rect 42172 4922 42196 4924
rect 42252 4922 42258 4924
rect 42012 4870 42014 4922
rect 42194 4870 42196 4922
rect 41950 4868 41956 4870
rect 42012 4868 42036 4870
rect 42092 4868 42116 4870
rect 42172 4868 42196 4870
rect 42252 4868 42258 4870
rect 41950 4859 42258 4868
rect 46950 4924 47258 4933
rect 46950 4922 46956 4924
rect 47012 4922 47036 4924
rect 47092 4922 47116 4924
rect 47172 4922 47196 4924
rect 47252 4922 47258 4924
rect 47012 4870 47014 4922
rect 47194 4870 47196 4922
rect 46950 4868 46956 4870
rect 47012 4868 47036 4870
rect 47092 4868 47116 4870
rect 47172 4868 47196 4870
rect 47252 4868 47258 4870
rect 46950 4859 47258 4868
rect 51950 4924 52258 4933
rect 51950 4922 51956 4924
rect 52012 4922 52036 4924
rect 52092 4922 52116 4924
rect 52172 4922 52196 4924
rect 52252 4922 52258 4924
rect 52012 4870 52014 4922
rect 52194 4870 52196 4922
rect 51950 4868 51956 4870
rect 52012 4868 52036 4870
rect 52092 4868 52116 4870
rect 52172 4868 52196 4870
rect 52252 4868 52258 4870
rect 51950 4859 52258 4868
rect 56950 4924 57258 4933
rect 58530 4927 58586 4936
rect 56950 4922 56956 4924
rect 57012 4922 57036 4924
rect 57092 4922 57116 4924
rect 57172 4922 57196 4924
rect 57252 4922 57258 4924
rect 57012 4870 57014 4922
rect 57194 4870 57196 4922
rect 56950 4868 56956 4870
rect 57012 4868 57036 4870
rect 57092 4868 57116 4870
rect 57172 4868 57196 4870
rect 57252 4868 57258 4870
rect 56950 4859 57258 4868
rect 58532 4616 58584 4622
rect 58532 4558 58584 4564
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 22610 4380 22918 4389
rect 22610 4378 22616 4380
rect 22672 4378 22696 4380
rect 22752 4378 22776 4380
rect 22832 4378 22856 4380
rect 22912 4378 22918 4380
rect 22672 4326 22674 4378
rect 22854 4326 22856 4378
rect 22610 4324 22616 4326
rect 22672 4324 22696 4326
rect 22752 4324 22776 4326
rect 22832 4324 22856 4326
rect 22912 4324 22918 4326
rect 22610 4315 22918 4324
rect 27610 4380 27918 4389
rect 27610 4378 27616 4380
rect 27672 4378 27696 4380
rect 27752 4378 27776 4380
rect 27832 4378 27856 4380
rect 27912 4378 27918 4380
rect 27672 4326 27674 4378
rect 27854 4326 27856 4378
rect 27610 4324 27616 4326
rect 27672 4324 27696 4326
rect 27752 4324 27776 4326
rect 27832 4324 27856 4326
rect 27912 4324 27918 4326
rect 27610 4315 27918 4324
rect 32610 4380 32918 4389
rect 32610 4378 32616 4380
rect 32672 4378 32696 4380
rect 32752 4378 32776 4380
rect 32832 4378 32856 4380
rect 32912 4378 32918 4380
rect 32672 4326 32674 4378
rect 32854 4326 32856 4378
rect 32610 4324 32616 4326
rect 32672 4324 32696 4326
rect 32752 4324 32776 4326
rect 32832 4324 32856 4326
rect 32912 4324 32918 4326
rect 32610 4315 32918 4324
rect 37610 4380 37918 4389
rect 37610 4378 37616 4380
rect 37672 4378 37696 4380
rect 37752 4378 37776 4380
rect 37832 4378 37856 4380
rect 37912 4378 37918 4380
rect 37672 4326 37674 4378
rect 37854 4326 37856 4378
rect 37610 4324 37616 4326
rect 37672 4324 37696 4326
rect 37752 4324 37776 4326
rect 37832 4324 37856 4326
rect 37912 4324 37918 4326
rect 37610 4315 37918 4324
rect 42610 4380 42918 4389
rect 42610 4378 42616 4380
rect 42672 4378 42696 4380
rect 42752 4378 42776 4380
rect 42832 4378 42856 4380
rect 42912 4378 42918 4380
rect 42672 4326 42674 4378
rect 42854 4326 42856 4378
rect 42610 4324 42616 4326
rect 42672 4324 42696 4326
rect 42752 4324 42776 4326
rect 42832 4324 42856 4326
rect 42912 4324 42918 4326
rect 42610 4315 42918 4324
rect 47610 4380 47918 4389
rect 47610 4378 47616 4380
rect 47672 4378 47696 4380
rect 47752 4378 47776 4380
rect 47832 4378 47856 4380
rect 47912 4378 47918 4380
rect 47672 4326 47674 4378
rect 47854 4326 47856 4378
rect 47610 4324 47616 4326
rect 47672 4324 47696 4326
rect 47752 4324 47776 4326
rect 47832 4324 47856 4326
rect 47912 4324 47918 4326
rect 47610 4315 47918 4324
rect 52610 4380 52918 4389
rect 52610 4378 52616 4380
rect 52672 4378 52696 4380
rect 52752 4378 52776 4380
rect 52832 4378 52856 4380
rect 52912 4378 52918 4380
rect 52672 4326 52674 4378
rect 52854 4326 52856 4378
rect 52610 4324 52616 4326
rect 52672 4324 52696 4326
rect 52752 4324 52776 4326
rect 52832 4324 52856 4326
rect 52912 4324 52918 4326
rect 52610 4315 52918 4324
rect 57610 4380 57918 4389
rect 57610 4378 57616 4380
rect 57672 4378 57696 4380
rect 57752 4378 57776 4380
rect 57832 4378 57856 4380
rect 57912 4378 57918 4380
rect 57672 4326 57674 4378
rect 57854 4326 57856 4378
rect 57610 4324 57616 4326
rect 57672 4324 57696 4326
rect 57752 4324 57776 4326
rect 57832 4324 57856 4326
rect 57912 4324 57918 4326
rect 57610 4315 57918 4324
rect 58544 4185 58572 4558
rect 58530 4176 58586 4185
rect 58530 4111 58586 4120
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 21950 3836 22258 3845
rect 21950 3834 21956 3836
rect 22012 3834 22036 3836
rect 22092 3834 22116 3836
rect 22172 3834 22196 3836
rect 22252 3834 22258 3836
rect 22012 3782 22014 3834
rect 22194 3782 22196 3834
rect 21950 3780 21956 3782
rect 22012 3780 22036 3782
rect 22092 3780 22116 3782
rect 22172 3780 22196 3782
rect 22252 3780 22258 3782
rect 21950 3771 22258 3780
rect 26950 3836 27258 3845
rect 26950 3834 26956 3836
rect 27012 3834 27036 3836
rect 27092 3834 27116 3836
rect 27172 3834 27196 3836
rect 27252 3834 27258 3836
rect 27012 3782 27014 3834
rect 27194 3782 27196 3834
rect 26950 3780 26956 3782
rect 27012 3780 27036 3782
rect 27092 3780 27116 3782
rect 27172 3780 27196 3782
rect 27252 3780 27258 3782
rect 26950 3771 27258 3780
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 36950 3836 37258 3845
rect 36950 3834 36956 3836
rect 37012 3834 37036 3836
rect 37092 3834 37116 3836
rect 37172 3834 37196 3836
rect 37252 3834 37258 3836
rect 37012 3782 37014 3834
rect 37194 3782 37196 3834
rect 36950 3780 36956 3782
rect 37012 3780 37036 3782
rect 37092 3780 37116 3782
rect 37172 3780 37196 3782
rect 37252 3780 37258 3782
rect 36950 3771 37258 3780
rect 41950 3836 42258 3845
rect 41950 3834 41956 3836
rect 42012 3834 42036 3836
rect 42092 3834 42116 3836
rect 42172 3834 42196 3836
rect 42252 3834 42258 3836
rect 42012 3782 42014 3834
rect 42194 3782 42196 3834
rect 41950 3780 41956 3782
rect 42012 3780 42036 3782
rect 42092 3780 42116 3782
rect 42172 3780 42196 3782
rect 42252 3780 42258 3782
rect 41950 3771 42258 3780
rect 46950 3836 47258 3845
rect 46950 3834 46956 3836
rect 47012 3834 47036 3836
rect 47092 3834 47116 3836
rect 47172 3834 47196 3836
rect 47252 3834 47258 3836
rect 47012 3782 47014 3834
rect 47194 3782 47196 3834
rect 46950 3780 46956 3782
rect 47012 3780 47036 3782
rect 47092 3780 47116 3782
rect 47172 3780 47196 3782
rect 47252 3780 47258 3782
rect 46950 3771 47258 3780
rect 51950 3836 52258 3845
rect 51950 3834 51956 3836
rect 52012 3834 52036 3836
rect 52092 3834 52116 3836
rect 52172 3834 52196 3836
rect 52252 3834 52258 3836
rect 52012 3782 52014 3834
rect 52194 3782 52196 3834
rect 51950 3780 51956 3782
rect 52012 3780 52036 3782
rect 52092 3780 52116 3782
rect 52172 3780 52196 3782
rect 52252 3780 52258 3782
rect 51950 3771 52258 3780
rect 56950 3836 57258 3845
rect 56950 3834 56956 3836
rect 57012 3834 57036 3836
rect 57092 3834 57116 3836
rect 57172 3834 57196 3836
rect 57252 3834 57258 3836
rect 57012 3782 57014 3834
rect 57194 3782 57196 3834
rect 56950 3780 56956 3782
rect 57012 3780 57036 3782
rect 57092 3780 57116 3782
rect 57172 3780 57196 3782
rect 57252 3780 57258 3782
rect 56950 3771 57258 3780
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 22610 3292 22918 3301
rect 22610 3290 22616 3292
rect 22672 3290 22696 3292
rect 22752 3290 22776 3292
rect 22832 3290 22856 3292
rect 22912 3290 22918 3292
rect 22672 3238 22674 3290
rect 22854 3238 22856 3290
rect 22610 3236 22616 3238
rect 22672 3236 22696 3238
rect 22752 3236 22776 3238
rect 22832 3236 22856 3238
rect 22912 3236 22918 3238
rect 22610 3227 22918 3236
rect 27610 3292 27918 3301
rect 27610 3290 27616 3292
rect 27672 3290 27696 3292
rect 27752 3290 27776 3292
rect 27832 3290 27856 3292
rect 27912 3290 27918 3292
rect 27672 3238 27674 3290
rect 27854 3238 27856 3290
rect 27610 3236 27616 3238
rect 27672 3236 27696 3238
rect 27752 3236 27776 3238
rect 27832 3236 27856 3238
rect 27912 3236 27918 3238
rect 27610 3227 27918 3236
rect 32610 3292 32918 3301
rect 32610 3290 32616 3292
rect 32672 3290 32696 3292
rect 32752 3290 32776 3292
rect 32832 3290 32856 3292
rect 32912 3290 32918 3292
rect 32672 3238 32674 3290
rect 32854 3238 32856 3290
rect 32610 3236 32616 3238
rect 32672 3236 32696 3238
rect 32752 3236 32776 3238
rect 32832 3236 32856 3238
rect 32912 3236 32918 3238
rect 32610 3227 32918 3236
rect 37610 3292 37918 3301
rect 37610 3290 37616 3292
rect 37672 3290 37696 3292
rect 37752 3290 37776 3292
rect 37832 3290 37856 3292
rect 37912 3290 37918 3292
rect 37672 3238 37674 3290
rect 37854 3238 37856 3290
rect 37610 3236 37616 3238
rect 37672 3236 37696 3238
rect 37752 3236 37776 3238
rect 37832 3236 37856 3238
rect 37912 3236 37918 3238
rect 37610 3227 37918 3236
rect 42610 3292 42918 3301
rect 42610 3290 42616 3292
rect 42672 3290 42696 3292
rect 42752 3290 42776 3292
rect 42832 3290 42856 3292
rect 42912 3290 42918 3292
rect 42672 3238 42674 3290
rect 42854 3238 42856 3290
rect 42610 3236 42616 3238
rect 42672 3236 42696 3238
rect 42752 3236 42776 3238
rect 42832 3236 42856 3238
rect 42912 3236 42918 3238
rect 42610 3227 42918 3236
rect 47610 3292 47918 3301
rect 47610 3290 47616 3292
rect 47672 3290 47696 3292
rect 47752 3290 47776 3292
rect 47832 3290 47856 3292
rect 47912 3290 47918 3292
rect 47672 3238 47674 3290
rect 47854 3238 47856 3290
rect 47610 3236 47616 3238
rect 47672 3236 47696 3238
rect 47752 3236 47776 3238
rect 47832 3236 47856 3238
rect 47912 3236 47918 3238
rect 47610 3227 47918 3236
rect 52610 3292 52918 3301
rect 52610 3290 52616 3292
rect 52672 3290 52696 3292
rect 52752 3290 52776 3292
rect 52832 3290 52856 3292
rect 52912 3290 52918 3292
rect 52672 3238 52674 3290
rect 52854 3238 52856 3290
rect 52610 3236 52616 3238
rect 52672 3236 52696 3238
rect 52752 3236 52776 3238
rect 52832 3236 52856 3238
rect 52912 3236 52918 3238
rect 52610 3227 52918 3236
rect 57610 3292 57918 3301
rect 57610 3290 57616 3292
rect 57672 3290 57696 3292
rect 57752 3290 57776 3292
rect 57832 3290 57856 3292
rect 57912 3290 57918 3292
rect 57672 3238 57674 3290
rect 57854 3238 57856 3290
rect 57610 3236 57616 3238
rect 57672 3236 57696 3238
rect 57752 3236 57776 3238
rect 57832 3236 57856 3238
rect 57912 3236 57918 3238
rect 57610 3227 57918 3236
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 21950 2748 22258 2757
rect 21950 2746 21956 2748
rect 22012 2746 22036 2748
rect 22092 2746 22116 2748
rect 22172 2746 22196 2748
rect 22252 2746 22258 2748
rect 22012 2694 22014 2746
rect 22194 2694 22196 2746
rect 21950 2692 21956 2694
rect 22012 2692 22036 2694
rect 22092 2692 22116 2694
rect 22172 2692 22196 2694
rect 22252 2692 22258 2694
rect 21950 2683 22258 2692
rect 26950 2748 27258 2757
rect 26950 2746 26956 2748
rect 27012 2746 27036 2748
rect 27092 2746 27116 2748
rect 27172 2746 27196 2748
rect 27252 2746 27258 2748
rect 27012 2694 27014 2746
rect 27194 2694 27196 2746
rect 26950 2692 26956 2694
rect 27012 2692 27036 2694
rect 27092 2692 27116 2694
rect 27172 2692 27196 2694
rect 27252 2692 27258 2694
rect 26950 2683 27258 2692
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 36950 2748 37258 2757
rect 36950 2746 36956 2748
rect 37012 2746 37036 2748
rect 37092 2746 37116 2748
rect 37172 2746 37196 2748
rect 37252 2746 37258 2748
rect 37012 2694 37014 2746
rect 37194 2694 37196 2746
rect 36950 2692 36956 2694
rect 37012 2692 37036 2694
rect 37092 2692 37116 2694
rect 37172 2692 37196 2694
rect 37252 2692 37258 2694
rect 36950 2683 37258 2692
rect 41950 2748 42258 2757
rect 41950 2746 41956 2748
rect 42012 2746 42036 2748
rect 42092 2746 42116 2748
rect 42172 2746 42196 2748
rect 42252 2746 42258 2748
rect 42012 2694 42014 2746
rect 42194 2694 42196 2746
rect 41950 2692 41956 2694
rect 42012 2692 42036 2694
rect 42092 2692 42116 2694
rect 42172 2692 42196 2694
rect 42252 2692 42258 2694
rect 41950 2683 42258 2692
rect 46950 2748 47258 2757
rect 46950 2746 46956 2748
rect 47012 2746 47036 2748
rect 47092 2746 47116 2748
rect 47172 2746 47196 2748
rect 47252 2746 47258 2748
rect 47012 2694 47014 2746
rect 47194 2694 47196 2746
rect 46950 2692 46956 2694
rect 47012 2692 47036 2694
rect 47092 2692 47116 2694
rect 47172 2692 47196 2694
rect 47252 2692 47258 2694
rect 46950 2683 47258 2692
rect 51950 2748 52258 2757
rect 51950 2746 51956 2748
rect 52012 2746 52036 2748
rect 52092 2746 52116 2748
rect 52172 2746 52196 2748
rect 52252 2746 52258 2748
rect 52012 2694 52014 2746
rect 52194 2694 52196 2746
rect 51950 2692 51956 2694
rect 52012 2692 52036 2694
rect 52092 2692 52116 2694
rect 52172 2692 52196 2694
rect 52252 2692 52258 2694
rect 51950 2683 52258 2692
rect 56950 2748 57258 2757
rect 56950 2746 56956 2748
rect 57012 2746 57036 2748
rect 57092 2746 57116 2748
rect 57172 2746 57196 2748
rect 57252 2746 57258 2748
rect 57012 2694 57014 2746
rect 57194 2694 57196 2746
rect 56950 2692 56956 2694
rect 57012 2692 57036 2694
rect 57092 2692 57116 2694
rect 57172 2692 57196 2694
rect 57252 2692 57258 2694
rect 56950 2683 57258 2692
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 17610 2204 17918 2213
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
rect 22610 2204 22918 2213
rect 22610 2202 22616 2204
rect 22672 2202 22696 2204
rect 22752 2202 22776 2204
rect 22832 2202 22856 2204
rect 22912 2202 22918 2204
rect 22672 2150 22674 2202
rect 22854 2150 22856 2202
rect 22610 2148 22616 2150
rect 22672 2148 22696 2150
rect 22752 2148 22776 2150
rect 22832 2148 22856 2150
rect 22912 2148 22918 2150
rect 22610 2139 22918 2148
rect 27610 2204 27918 2213
rect 27610 2202 27616 2204
rect 27672 2202 27696 2204
rect 27752 2202 27776 2204
rect 27832 2202 27856 2204
rect 27912 2202 27918 2204
rect 27672 2150 27674 2202
rect 27854 2150 27856 2202
rect 27610 2148 27616 2150
rect 27672 2148 27696 2150
rect 27752 2148 27776 2150
rect 27832 2148 27856 2150
rect 27912 2148 27918 2150
rect 27610 2139 27918 2148
rect 32610 2204 32918 2213
rect 32610 2202 32616 2204
rect 32672 2202 32696 2204
rect 32752 2202 32776 2204
rect 32832 2202 32856 2204
rect 32912 2202 32918 2204
rect 32672 2150 32674 2202
rect 32854 2150 32856 2202
rect 32610 2148 32616 2150
rect 32672 2148 32696 2150
rect 32752 2148 32776 2150
rect 32832 2148 32856 2150
rect 32912 2148 32918 2150
rect 32610 2139 32918 2148
rect 37610 2204 37918 2213
rect 37610 2202 37616 2204
rect 37672 2202 37696 2204
rect 37752 2202 37776 2204
rect 37832 2202 37856 2204
rect 37912 2202 37918 2204
rect 37672 2150 37674 2202
rect 37854 2150 37856 2202
rect 37610 2148 37616 2150
rect 37672 2148 37696 2150
rect 37752 2148 37776 2150
rect 37832 2148 37856 2150
rect 37912 2148 37918 2150
rect 37610 2139 37918 2148
rect 42610 2204 42918 2213
rect 42610 2202 42616 2204
rect 42672 2202 42696 2204
rect 42752 2202 42776 2204
rect 42832 2202 42856 2204
rect 42912 2202 42918 2204
rect 42672 2150 42674 2202
rect 42854 2150 42856 2202
rect 42610 2148 42616 2150
rect 42672 2148 42696 2150
rect 42752 2148 42776 2150
rect 42832 2148 42856 2150
rect 42912 2148 42918 2150
rect 42610 2139 42918 2148
rect 47610 2204 47918 2213
rect 47610 2202 47616 2204
rect 47672 2202 47696 2204
rect 47752 2202 47776 2204
rect 47832 2202 47856 2204
rect 47912 2202 47918 2204
rect 47672 2150 47674 2202
rect 47854 2150 47856 2202
rect 47610 2148 47616 2150
rect 47672 2148 47696 2150
rect 47752 2148 47776 2150
rect 47832 2148 47856 2150
rect 47912 2148 47918 2150
rect 47610 2139 47918 2148
rect 52610 2204 52918 2213
rect 52610 2202 52616 2204
rect 52672 2202 52696 2204
rect 52752 2202 52776 2204
rect 52832 2202 52856 2204
rect 52912 2202 52918 2204
rect 52672 2150 52674 2202
rect 52854 2150 52856 2202
rect 52610 2148 52616 2150
rect 52672 2148 52696 2150
rect 52752 2148 52776 2150
rect 52832 2148 52856 2150
rect 52912 2148 52918 2150
rect 52610 2139 52918 2148
rect 57610 2204 57918 2213
rect 57610 2202 57616 2204
rect 57672 2202 57696 2204
rect 57752 2202 57776 2204
rect 57832 2202 57856 2204
rect 57912 2202 57918 2204
rect 57672 2150 57674 2202
rect 57854 2150 57856 2202
rect 57610 2148 57616 2150
rect 57672 2148 57696 2150
rect 57752 2148 57776 2150
rect 57832 2148 57856 2150
rect 57912 2148 57918 2150
rect 57610 2139 57918 2148
<< via2 >>
rect 2616 57690 2672 57692
rect 2696 57690 2752 57692
rect 2776 57690 2832 57692
rect 2856 57690 2912 57692
rect 2616 57638 2662 57690
rect 2662 57638 2672 57690
rect 2696 57638 2726 57690
rect 2726 57638 2738 57690
rect 2738 57638 2752 57690
rect 2776 57638 2790 57690
rect 2790 57638 2802 57690
rect 2802 57638 2832 57690
rect 2856 57638 2866 57690
rect 2866 57638 2912 57690
rect 2616 57636 2672 57638
rect 2696 57636 2752 57638
rect 2776 57636 2832 57638
rect 2856 57636 2912 57638
rect 7616 57690 7672 57692
rect 7696 57690 7752 57692
rect 7776 57690 7832 57692
rect 7856 57690 7912 57692
rect 7616 57638 7662 57690
rect 7662 57638 7672 57690
rect 7696 57638 7726 57690
rect 7726 57638 7738 57690
rect 7738 57638 7752 57690
rect 7776 57638 7790 57690
rect 7790 57638 7802 57690
rect 7802 57638 7832 57690
rect 7856 57638 7866 57690
rect 7866 57638 7912 57690
rect 7616 57636 7672 57638
rect 7696 57636 7752 57638
rect 7776 57636 7832 57638
rect 7856 57636 7912 57638
rect 12616 57690 12672 57692
rect 12696 57690 12752 57692
rect 12776 57690 12832 57692
rect 12856 57690 12912 57692
rect 12616 57638 12662 57690
rect 12662 57638 12672 57690
rect 12696 57638 12726 57690
rect 12726 57638 12738 57690
rect 12738 57638 12752 57690
rect 12776 57638 12790 57690
rect 12790 57638 12802 57690
rect 12802 57638 12832 57690
rect 12856 57638 12866 57690
rect 12866 57638 12912 57690
rect 12616 57636 12672 57638
rect 12696 57636 12752 57638
rect 12776 57636 12832 57638
rect 12856 57636 12912 57638
rect 17616 57690 17672 57692
rect 17696 57690 17752 57692
rect 17776 57690 17832 57692
rect 17856 57690 17912 57692
rect 17616 57638 17662 57690
rect 17662 57638 17672 57690
rect 17696 57638 17726 57690
rect 17726 57638 17738 57690
rect 17738 57638 17752 57690
rect 17776 57638 17790 57690
rect 17790 57638 17802 57690
rect 17802 57638 17832 57690
rect 17856 57638 17866 57690
rect 17866 57638 17912 57690
rect 17616 57636 17672 57638
rect 17696 57636 17752 57638
rect 17776 57636 17832 57638
rect 17856 57636 17912 57638
rect 22616 57690 22672 57692
rect 22696 57690 22752 57692
rect 22776 57690 22832 57692
rect 22856 57690 22912 57692
rect 22616 57638 22662 57690
rect 22662 57638 22672 57690
rect 22696 57638 22726 57690
rect 22726 57638 22738 57690
rect 22738 57638 22752 57690
rect 22776 57638 22790 57690
rect 22790 57638 22802 57690
rect 22802 57638 22832 57690
rect 22856 57638 22866 57690
rect 22866 57638 22912 57690
rect 22616 57636 22672 57638
rect 22696 57636 22752 57638
rect 22776 57636 22832 57638
rect 22856 57636 22912 57638
rect 27616 57690 27672 57692
rect 27696 57690 27752 57692
rect 27776 57690 27832 57692
rect 27856 57690 27912 57692
rect 27616 57638 27662 57690
rect 27662 57638 27672 57690
rect 27696 57638 27726 57690
rect 27726 57638 27738 57690
rect 27738 57638 27752 57690
rect 27776 57638 27790 57690
rect 27790 57638 27802 57690
rect 27802 57638 27832 57690
rect 27856 57638 27866 57690
rect 27866 57638 27912 57690
rect 27616 57636 27672 57638
rect 27696 57636 27752 57638
rect 27776 57636 27832 57638
rect 27856 57636 27912 57638
rect 32616 57690 32672 57692
rect 32696 57690 32752 57692
rect 32776 57690 32832 57692
rect 32856 57690 32912 57692
rect 32616 57638 32662 57690
rect 32662 57638 32672 57690
rect 32696 57638 32726 57690
rect 32726 57638 32738 57690
rect 32738 57638 32752 57690
rect 32776 57638 32790 57690
rect 32790 57638 32802 57690
rect 32802 57638 32832 57690
rect 32856 57638 32866 57690
rect 32866 57638 32912 57690
rect 32616 57636 32672 57638
rect 32696 57636 32752 57638
rect 32776 57636 32832 57638
rect 32856 57636 32912 57638
rect 37616 57690 37672 57692
rect 37696 57690 37752 57692
rect 37776 57690 37832 57692
rect 37856 57690 37912 57692
rect 37616 57638 37662 57690
rect 37662 57638 37672 57690
rect 37696 57638 37726 57690
rect 37726 57638 37738 57690
rect 37738 57638 37752 57690
rect 37776 57638 37790 57690
rect 37790 57638 37802 57690
rect 37802 57638 37832 57690
rect 37856 57638 37866 57690
rect 37866 57638 37912 57690
rect 37616 57636 37672 57638
rect 37696 57636 37752 57638
rect 37776 57636 37832 57638
rect 37856 57636 37912 57638
rect 42616 57690 42672 57692
rect 42696 57690 42752 57692
rect 42776 57690 42832 57692
rect 42856 57690 42912 57692
rect 42616 57638 42662 57690
rect 42662 57638 42672 57690
rect 42696 57638 42726 57690
rect 42726 57638 42738 57690
rect 42738 57638 42752 57690
rect 42776 57638 42790 57690
rect 42790 57638 42802 57690
rect 42802 57638 42832 57690
rect 42856 57638 42866 57690
rect 42866 57638 42912 57690
rect 42616 57636 42672 57638
rect 42696 57636 42752 57638
rect 42776 57636 42832 57638
rect 42856 57636 42912 57638
rect 47616 57690 47672 57692
rect 47696 57690 47752 57692
rect 47776 57690 47832 57692
rect 47856 57690 47912 57692
rect 47616 57638 47662 57690
rect 47662 57638 47672 57690
rect 47696 57638 47726 57690
rect 47726 57638 47738 57690
rect 47738 57638 47752 57690
rect 47776 57638 47790 57690
rect 47790 57638 47802 57690
rect 47802 57638 47832 57690
rect 47856 57638 47866 57690
rect 47866 57638 47912 57690
rect 47616 57636 47672 57638
rect 47696 57636 47752 57638
rect 47776 57636 47832 57638
rect 47856 57636 47912 57638
rect 52616 57690 52672 57692
rect 52696 57690 52752 57692
rect 52776 57690 52832 57692
rect 52856 57690 52912 57692
rect 52616 57638 52662 57690
rect 52662 57638 52672 57690
rect 52696 57638 52726 57690
rect 52726 57638 52738 57690
rect 52738 57638 52752 57690
rect 52776 57638 52790 57690
rect 52790 57638 52802 57690
rect 52802 57638 52832 57690
rect 52856 57638 52866 57690
rect 52866 57638 52912 57690
rect 52616 57636 52672 57638
rect 52696 57636 52752 57638
rect 52776 57636 52832 57638
rect 52856 57636 52912 57638
rect 57616 57690 57672 57692
rect 57696 57690 57752 57692
rect 57776 57690 57832 57692
rect 57856 57690 57912 57692
rect 57616 57638 57662 57690
rect 57662 57638 57672 57690
rect 57696 57638 57726 57690
rect 57726 57638 57738 57690
rect 57738 57638 57752 57690
rect 57776 57638 57790 57690
rect 57790 57638 57802 57690
rect 57802 57638 57832 57690
rect 57856 57638 57866 57690
rect 57866 57638 57912 57690
rect 57616 57636 57672 57638
rect 57696 57636 57752 57638
rect 57776 57636 57832 57638
rect 57856 57636 57912 57638
rect 1956 57146 2012 57148
rect 2036 57146 2092 57148
rect 2116 57146 2172 57148
rect 2196 57146 2252 57148
rect 1956 57094 2002 57146
rect 2002 57094 2012 57146
rect 2036 57094 2066 57146
rect 2066 57094 2078 57146
rect 2078 57094 2092 57146
rect 2116 57094 2130 57146
rect 2130 57094 2142 57146
rect 2142 57094 2172 57146
rect 2196 57094 2206 57146
rect 2206 57094 2252 57146
rect 1956 57092 2012 57094
rect 2036 57092 2092 57094
rect 2116 57092 2172 57094
rect 2196 57092 2252 57094
rect 6956 57146 7012 57148
rect 7036 57146 7092 57148
rect 7116 57146 7172 57148
rect 7196 57146 7252 57148
rect 6956 57094 7002 57146
rect 7002 57094 7012 57146
rect 7036 57094 7066 57146
rect 7066 57094 7078 57146
rect 7078 57094 7092 57146
rect 7116 57094 7130 57146
rect 7130 57094 7142 57146
rect 7142 57094 7172 57146
rect 7196 57094 7206 57146
rect 7206 57094 7252 57146
rect 6956 57092 7012 57094
rect 7036 57092 7092 57094
rect 7116 57092 7172 57094
rect 7196 57092 7252 57094
rect 11956 57146 12012 57148
rect 12036 57146 12092 57148
rect 12116 57146 12172 57148
rect 12196 57146 12252 57148
rect 11956 57094 12002 57146
rect 12002 57094 12012 57146
rect 12036 57094 12066 57146
rect 12066 57094 12078 57146
rect 12078 57094 12092 57146
rect 12116 57094 12130 57146
rect 12130 57094 12142 57146
rect 12142 57094 12172 57146
rect 12196 57094 12206 57146
rect 12206 57094 12252 57146
rect 11956 57092 12012 57094
rect 12036 57092 12092 57094
rect 12116 57092 12172 57094
rect 12196 57092 12252 57094
rect 16956 57146 17012 57148
rect 17036 57146 17092 57148
rect 17116 57146 17172 57148
rect 17196 57146 17252 57148
rect 16956 57094 17002 57146
rect 17002 57094 17012 57146
rect 17036 57094 17066 57146
rect 17066 57094 17078 57146
rect 17078 57094 17092 57146
rect 17116 57094 17130 57146
rect 17130 57094 17142 57146
rect 17142 57094 17172 57146
rect 17196 57094 17206 57146
rect 17206 57094 17252 57146
rect 16956 57092 17012 57094
rect 17036 57092 17092 57094
rect 17116 57092 17172 57094
rect 17196 57092 17252 57094
rect 21956 57146 22012 57148
rect 22036 57146 22092 57148
rect 22116 57146 22172 57148
rect 22196 57146 22252 57148
rect 21956 57094 22002 57146
rect 22002 57094 22012 57146
rect 22036 57094 22066 57146
rect 22066 57094 22078 57146
rect 22078 57094 22092 57146
rect 22116 57094 22130 57146
rect 22130 57094 22142 57146
rect 22142 57094 22172 57146
rect 22196 57094 22206 57146
rect 22206 57094 22252 57146
rect 21956 57092 22012 57094
rect 22036 57092 22092 57094
rect 22116 57092 22172 57094
rect 22196 57092 22252 57094
rect 26956 57146 27012 57148
rect 27036 57146 27092 57148
rect 27116 57146 27172 57148
rect 27196 57146 27252 57148
rect 26956 57094 27002 57146
rect 27002 57094 27012 57146
rect 27036 57094 27066 57146
rect 27066 57094 27078 57146
rect 27078 57094 27092 57146
rect 27116 57094 27130 57146
rect 27130 57094 27142 57146
rect 27142 57094 27172 57146
rect 27196 57094 27206 57146
rect 27206 57094 27252 57146
rect 26956 57092 27012 57094
rect 27036 57092 27092 57094
rect 27116 57092 27172 57094
rect 27196 57092 27252 57094
rect 31956 57146 32012 57148
rect 32036 57146 32092 57148
rect 32116 57146 32172 57148
rect 32196 57146 32252 57148
rect 31956 57094 32002 57146
rect 32002 57094 32012 57146
rect 32036 57094 32066 57146
rect 32066 57094 32078 57146
rect 32078 57094 32092 57146
rect 32116 57094 32130 57146
rect 32130 57094 32142 57146
rect 32142 57094 32172 57146
rect 32196 57094 32206 57146
rect 32206 57094 32252 57146
rect 31956 57092 32012 57094
rect 32036 57092 32092 57094
rect 32116 57092 32172 57094
rect 32196 57092 32252 57094
rect 36956 57146 37012 57148
rect 37036 57146 37092 57148
rect 37116 57146 37172 57148
rect 37196 57146 37252 57148
rect 36956 57094 37002 57146
rect 37002 57094 37012 57146
rect 37036 57094 37066 57146
rect 37066 57094 37078 57146
rect 37078 57094 37092 57146
rect 37116 57094 37130 57146
rect 37130 57094 37142 57146
rect 37142 57094 37172 57146
rect 37196 57094 37206 57146
rect 37206 57094 37252 57146
rect 36956 57092 37012 57094
rect 37036 57092 37092 57094
rect 37116 57092 37172 57094
rect 37196 57092 37252 57094
rect 41956 57146 42012 57148
rect 42036 57146 42092 57148
rect 42116 57146 42172 57148
rect 42196 57146 42252 57148
rect 41956 57094 42002 57146
rect 42002 57094 42012 57146
rect 42036 57094 42066 57146
rect 42066 57094 42078 57146
rect 42078 57094 42092 57146
rect 42116 57094 42130 57146
rect 42130 57094 42142 57146
rect 42142 57094 42172 57146
rect 42196 57094 42206 57146
rect 42206 57094 42252 57146
rect 41956 57092 42012 57094
rect 42036 57092 42092 57094
rect 42116 57092 42172 57094
rect 42196 57092 42252 57094
rect 46956 57146 47012 57148
rect 47036 57146 47092 57148
rect 47116 57146 47172 57148
rect 47196 57146 47252 57148
rect 46956 57094 47002 57146
rect 47002 57094 47012 57146
rect 47036 57094 47066 57146
rect 47066 57094 47078 57146
rect 47078 57094 47092 57146
rect 47116 57094 47130 57146
rect 47130 57094 47142 57146
rect 47142 57094 47172 57146
rect 47196 57094 47206 57146
rect 47206 57094 47252 57146
rect 46956 57092 47012 57094
rect 47036 57092 47092 57094
rect 47116 57092 47172 57094
rect 47196 57092 47252 57094
rect 51956 57146 52012 57148
rect 52036 57146 52092 57148
rect 52116 57146 52172 57148
rect 52196 57146 52252 57148
rect 51956 57094 52002 57146
rect 52002 57094 52012 57146
rect 52036 57094 52066 57146
rect 52066 57094 52078 57146
rect 52078 57094 52092 57146
rect 52116 57094 52130 57146
rect 52130 57094 52142 57146
rect 52142 57094 52172 57146
rect 52196 57094 52206 57146
rect 52206 57094 52252 57146
rect 51956 57092 52012 57094
rect 52036 57092 52092 57094
rect 52116 57092 52172 57094
rect 52196 57092 52252 57094
rect 56956 57146 57012 57148
rect 57036 57146 57092 57148
rect 57116 57146 57172 57148
rect 57196 57146 57252 57148
rect 56956 57094 57002 57146
rect 57002 57094 57012 57146
rect 57036 57094 57066 57146
rect 57066 57094 57078 57146
rect 57078 57094 57092 57146
rect 57116 57094 57130 57146
rect 57130 57094 57142 57146
rect 57142 57094 57172 57146
rect 57196 57094 57206 57146
rect 57206 57094 57252 57146
rect 56956 57092 57012 57094
rect 57036 57092 57092 57094
rect 57116 57092 57172 57094
rect 57196 57092 57252 57094
rect 2616 56602 2672 56604
rect 2696 56602 2752 56604
rect 2776 56602 2832 56604
rect 2856 56602 2912 56604
rect 2616 56550 2662 56602
rect 2662 56550 2672 56602
rect 2696 56550 2726 56602
rect 2726 56550 2738 56602
rect 2738 56550 2752 56602
rect 2776 56550 2790 56602
rect 2790 56550 2802 56602
rect 2802 56550 2832 56602
rect 2856 56550 2866 56602
rect 2866 56550 2912 56602
rect 2616 56548 2672 56550
rect 2696 56548 2752 56550
rect 2776 56548 2832 56550
rect 2856 56548 2912 56550
rect 7616 56602 7672 56604
rect 7696 56602 7752 56604
rect 7776 56602 7832 56604
rect 7856 56602 7912 56604
rect 7616 56550 7662 56602
rect 7662 56550 7672 56602
rect 7696 56550 7726 56602
rect 7726 56550 7738 56602
rect 7738 56550 7752 56602
rect 7776 56550 7790 56602
rect 7790 56550 7802 56602
rect 7802 56550 7832 56602
rect 7856 56550 7866 56602
rect 7866 56550 7912 56602
rect 7616 56548 7672 56550
rect 7696 56548 7752 56550
rect 7776 56548 7832 56550
rect 7856 56548 7912 56550
rect 12616 56602 12672 56604
rect 12696 56602 12752 56604
rect 12776 56602 12832 56604
rect 12856 56602 12912 56604
rect 12616 56550 12662 56602
rect 12662 56550 12672 56602
rect 12696 56550 12726 56602
rect 12726 56550 12738 56602
rect 12738 56550 12752 56602
rect 12776 56550 12790 56602
rect 12790 56550 12802 56602
rect 12802 56550 12832 56602
rect 12856 56550 12866 56602
rect 12866 56550 12912 56602
rect 12616 56548 12672 56550
rect 12696 56548 12752 56550
rect 12776 56548 12832 56550
rect 12856 56548 12912 56550
rect 17616 56602 17672 56604
rect 17696 56602 17752 56604
rect 17776 56602 17832 56604
rect 17856 56602 17912 56604
rect 17616 56550 17662 56602
rect 17662 56550 17672 56602
rect 17696 56550 17726 56602
rect 17726 56550 17738 56602
rect 17738 56550 17752 56602
rect 17776 56550 17790 56602
rect 17790 56550 17802 56602
rect 17802 56550 17832 56602
rect 17856 56550 17866 56602
rect 17866 56550 17912 56602
rect 17616 56548 17672 56550
rect 17696 56548 17752 56550
rect 17776 56548 17832 56550
rect 17856 56548 17912 56550
rect 22616 56602 22672 56604
rect 22696 56602 22752 56604
rect 22776 56602 22832 56604
rect 22856 56602 22912 56604
rect 22616 56550 22662 56602
rect 22662 56550 22672 56602
rect 22696 56550 22726 56602
rect 22726 56550 22738 56602
rect 22738 56550 22752 56602
rect 22776 56550 22790 56602
rect 22790 56550 22802 56602
rect 22802 56550 22832 56602
rect 22856 56550 22866 56602
rect 22866 56550 22912 56602
rect 22616 56548 22672 56550
rect 22696 56548 22752 56550
rect 22776 56548 22832 56550
rect 22856 56548 22912 56550
rect 27616 56602 27672 56604
rect 27696 56602 27752 56604
rect 27776 56602 27832 56604
rect 27856 56602 27912 56604
rect 27616 56550 27662 56602
rect 27662 56550 27672 56602
rect 27696 56550 27726 56602
rect 27726 56550 27738 56602
rect 27738 56550 27752 56602
rect 27776 56550 27790 56602
rect 27790 56550 27802 56602
rect 27802 56550 27832 56602
rect 27856 56550 27866 56602
rect 27866 56550 27912 56602
rect 27616 56548 27672 56550
rect 27696 56548 27752 56550
rect 27776 56548 27832 56550
rect 27856 56548 27912 56550
rect 32616 56602 32672 56604
rect 32696 56602 32752 56604
rect 32776 56602 32832 56604
rect 32856 56602 32912 56604
rect 32616 56550 32662 56602
rect 32662 56550 32672 56602
rect 32696 56550 32726 56602
rect 32726 56550 32738 56602
rect 32738 56550 32752 56602
rect 32776 56550 32790 56602
rect 32790 56550 32802 56602
rect 32802 56550 32832 56602
rect 32856 56550 32866 56602
rect 32866 56550 32912 56602
rect 32616 56548 32672 56550
rect 32696 56548 32752 56550
rect 32776 56548 32832 56550
rect 32856 56548 32912 56550
rect 37616 56602 37672 56604
rect 37696 56602 37752 56604
rect 37776 56602 37832 56604
rect 37856 56602 37912 56604
rect 37616 56550 37662 56602
rect 37662 56550 37672 56602
rect 37696 56550 37726 56602
rect 37726 56550 37738 56602
rect 37738 56550 37752 56602
rect 37776 56550 37790 56602
rect 37790 56550 37802 56602
rect 37802 56550 37832 56602
rect 37856 56550 37866 56602
rect 37866 56550 37912 56602
rect 37616 56548 37672 56550
rect 37696 56548 37752 56550
rect 37776 56548 37832 56550
rect 37856 56548 37912 56550
rect 42616 56602 42672 56604
rect 42696 56602 42752 56604
rect 42776 56602 42832 56604
rect 42856 56602 42912 56604
rect 42616 56550 42662 56602
rect 42662 56550 42672 56602
rect 42696 56550 42726 56602
rect 42726 56550 42738 56602
rect 42738 56550 42752 56602
rect 42776 56550 42790 56602
rect 42790 56550 42802 56602
rect 42802 56550 42832 56602
rect 42856 56550 42866 56602
rect 42866 56550 42912 56602
rect 42616 56548 42672 56550
rect 42696 56548 42752 56550
rect 42776 56548 42832 56550
rect 42856 56548 42912 56550
rect 47616 56602 47672 56604
rect 47696 56602 47752 56604
rect 47776 56602 47832 56604
rect 47856 56602 47912 56604
rect 47616 56550 47662 56602
rect 47662 56550 47672 56602
rect 47696 56550 47726 56602
rect 47726 56550 47738 56602
rect 47738 56550 47752 56602
rect 47776 56550 47790 56602
rect 47790 56550 47802 56602
rect 47802 56550 47832 56602
rect 47856 56550 47866 56602
rect 47866 56550 47912 56602
rect 47616 56548 47672 56550
rect 47696 56548 47752 56550
rect 47776 56548 47832 56550
rect 47856 56548 47912 56550
rect 52616 56602 52672 56604
rect 52696 56602 52752 56604
rect 52776 56602 52832 56604
rect 52856 56602 52912 56604
rect 52616 56550 52662 56602
rect 52662 56550 52672 56602
rect 52696 56550 52726 56602
rect 52726 56550 52738 56602
rect 52738 56550 52752 56602
rect 52776 56550 52790 56602
rect 52790 56550 52802 56602
rect 52802 56550 52832 56602
rect 52856 56550 52866 56602
rect 52866 56550 52912 56602
rect 52616 56548 52672 56550
rect 52696 56548 52752 56550
rect 52776 56548 52832 56550
rect 52856 56548 52912 56550
rect 57616 56602 57672 56604
rect 57696 56602 57752 56604
rect 57776 56602 57832 56604
rect 57856 56602 57912 56604
rect 57616 56550 57662 56602
rect 57662 56550 57672 56602
rect 57696 56550 57726 56602
rect 57726 56550 57738 56602
rect 57738 56550 57752 56602
rect 57776 56550 57790 56602
rect 57790 56550 57802 56602
rect 57802 56550 57832 56602
rect 57856 56550 57866 56602
rect 57866 56550 57912 56602
rect 57616 56548 57672 56550
rect 57696 56548 57752 56550
rect 57776 56548 57832 56550
rect 57856 56548 57912 56550
rect 1956 56058 2012 56060
rect 2036 56058 2092 56060
rect 2116 56058 2172 56060
rect 2196 56058 2252 56060
rect 1956 56006 2002 56058
rect 2002 56006 2012 56058
rect 2036 56006 2066 56058
rect 2066 56006 2078 56058
rect 2078 56006 2092 56058
rect 2116 56006 2130 56058
rect 2130 56006 2142 56058
rect 2142 56006 2172 56058
rect 2196 56006 2206 56058
rect 2206 56006 2252 56058
rect 1956 56004 2012 56006
rect 2036 56004 2092 56006
rect 2116 56004 2172 56006
rect 2196 56004 2252 56006
rect 6956 56058 7012 56060
rect 7036 56058 7092 56060
rect 7116 56058 7172 56060
rect 7196 56058 7252 56060
rect 6956 56006 7002 56058
rect 7002 56006 7012 56058
rect 7036 56006 7066 56058
rect 7066 56006 7078 56058
rect 7078 56006 7092 56058
rect 7116 56006 7130 56058
rect 7130 56006 7142 56058
rect 7142 56006 7172 56058
rect 7196 56006 7206 56058
rect 7206 56006 7252 56058
rect 6956 56004 7012 56006
rect 7036 56004 7092 56006
rect 7116 56004 7172 56006
rect 7196 56004 7252 56006
rect 11956 56058 12012 56060
rect 12036 56058 12092 56060
rect 12116 56058 12172 56060
rect 12196 56058 12252 56060
rect 11956 56006 12002 56058
rect 12002 56006 12012 56058
rect 12036 56006 12066 56058
rect 12066 56006 12078 56058
rect 12078 56006 12092 56058
rect 12116 56006 12130 56058
rect 12130 56006 12142 56058
rect 12142 56006 12172 56058
rect 12196 56006 12206 56058
rect 12206 56006 12252 56058
rect 11956 56004 12012 56006
rect 12036 56004 12092 56006
rect 12116 56004 12172 56006
rect 12196 56004 12252 56006
rect 16956 56058 17012 56060
rect 17036 56058 17092 56060
rect 17116 56058 17172 56060
rect 17196 56058 17252 56060
rect 16956 56006 17002 56058
rect 17002 56006 17012 56058
rect 17036 56006 17066 56058
rect 17066 56006 17078 56058
rect 17078 56006 17092 56058
rect 17116 56006 17130 56058
rect 17130 56006 17142 56058
rect 17142 56006 17172 56058
rect 17196 56006 17206 56058
rect 17206 56006 17252 56058
rect 16956 56004 17012 56006
rect 17036 56004 17092 56006
rect 17116 56004 17172 56006
rect 17196 56004 17252 56006
rect 21956 56058 22012 56060
rect 22036 56058 22092 56060
rect 22116 56058 22172 56060
rect 22196 56058 22252 56060
rect 21956 56006 22002 56058
rect 22002 56006 22012 56058
rect 22036 56006 22066 56058
rect 22066 56006 22078 56058
rect 22078 56006 22092 56058
rect 22116 56006 22130 56058
rect 22130 56006 22142 56058
rect 22142 56006 22172 56058
rect 22196 56006 22206 56058
rect 22206 56006 22252 56058
rect 21956 56004 22012 56006
rect 22036 56004 22092 56006
rect 22116 56004 22172 56006
rect 22196 56004 22252 56006
rect 26956 56058 27012 56060
rect 27036 56058 27092 56060
rect 27116 56058 27172 56060
rect 27196 56058 27252 56060
rect 26956 56006 27002 56058
rect 27002 56006 27012 56058
rect 27036 56006 27066 56058
rect 27066 56006 27078 56058
rect 27078 56006 27092 56058
rect 27116 56006 27130 56058
rect 27130 56006 27142 56058
rect 27142 56006 27172 56058
rect 27196 56006 27206 56058
rect 27206 56006 27252 56058
rect 26956 56004 27012 56006
rect 27036 56004 27092 56006
rect 27116 56004 27172 56006
rect 27196 56004 27252 56006
rect 31956 56058 32012 56060
rect 32036 56058 32092 56060
rect 32116 56058 32172 56060
rect 32196 56058 32252 56060
rect 31956 56006 32002 56058
rect 32002 56006 32012 56058
rect 32036 56006 32066 56058
rect 32066 56006 32078 56058
rect 32078 56006 32092 56058
rect 32116 56006 32130 56058
rect 32130 56006 32142 56058
rect 32142 56006 32172 56058
rect 32196 56006 32206 56058
rect 32206 56006 32252 56058
rect 31956 56004 32012 56006
rect 32036 56004 32092 56006
rect 32116 56004 32172 56006
rect 32196 56004 32252 56006
rect 36956 56058 37012 56060
rect 37036 56058 37092 56060
rect 37116 56058 37172 56060
rect 37196 56058 37252 56060
rect 36956 56006 37002 56058
rect 37002 56006 37012 56058
rect 37036 56006 37066 56058
rect 37066 56006 37078 56058
rect 37078 56006 37092 56058
rect 37116 56006 37130 56058
rect 37130 56006 37142 56058
rect 37142 56006 37172 56058
rect 37196 56006 37206 56058
rect 37206 56006 37252 56058
rect 36956 56004 37012 56006
rect 37036 56004 37092 56006
rect 37116 56004 37172 56006
rect 37196 56004 37252 56006
rect 41956 56058 42012 56060
rect 42036 56058 42092 56060
rect 42116 56058 42172 56060
rect 42196 56058 42252 56060
rect 41956 56006 42002 56058
rect 42002 56006 42012 56058
rect 42036 56006 42066 56058
rect 42066 56006 42078 56058
rect 42078 56006 42092 56058
rect 42116 56006 42130 56058
rect 42130 56006 42142 56058
rect 42142 56006 42172 56058
rect 42196 56006 42206 56058
rect 42206 56006 42252 56058
rect 41956 56004 42012 56006
rect 42036 56004 42092 56006
rect 42116 56004 42172 56006
rect 42196 56004 42252 56006
rect 46956 56058 47012 56060
rect 47036 56058 47092 56060
rect 47116 56058 47172 56060
rect 47196 56058 47252 56060
rect 46956 56006 47002 56058
rect 47002 56006 47012 56058
rect 47036 56006 47066 56058
rect 47066 56006 47078 56058
rect 47078 56006 47092 56058
rect 47116 56006 47130 56058
rect 47130 56006 47142 56058
rect 47142 56006 47172 56058
rect 47196 56006 47206 56058
rect 47206 56006 47252 56058
rect 46956 56004 47012 56006
rect 47036 56004 47092 56006
rect 47116 56004 47172 56006
rect 47196 56004 47252 56006
rect 51956 56058 52012 56060
rect 52036 56058 52092 56060
rect 52116 56058 52172 56060
rect 52196 56058 52252 56060
rect 51956 56006 52002 56058
rect 52002 56006 52012 56058
rect 52036 56006 52066 56058
rect 52066 56006 52078 56058
rect 52078 56006 52092 56058
rect 52116 56006 52130 56058
rect 52130 56006 52142 56058
rect 52142 56006 52172 56058
rect 52196 56006 52206 56058
rect 52206 56006 52252 56058
rect 51956 56004 52012 56006
rect 52036 56004 52092 56006
rect 52116 56004 52172 56006
rect 52196 56004 52252 56006
rect 56956 56058 57012 56060
rect 57036 56058 57092 56060
rect 57116 56058 57172 56060
rect 57196 56058 57252 56060
rect 56956 56006 57002 56058
rect 57002 56006 57012 56058
rect 57036 56006 57066 56058
rect 57066 56006 57078 56058
rect 57078 56006 57092 56058
rect 57116 56006 57130 56058
rect 57130 56006 57142 56058
rect 57142 56006 57172 56058
rect 57196 56006 57206 56058
rect 57206 56006 57252 56058
rect 56956 56004 57012 56006
rect 57036 56004 57092 56006
rect 57116 56004 57172 56006
rect 57196 56004 57252 56006
rect 58530 55528 58586 55584
rect 2616 55514 2672 55516
rect 2696 55514 2752 55516
rect 2776 55514 2832 55516
rect 2856 55514 2912 55516
rect 2616 55462 2662 55514
rect 2662 55462 2672 55514
rect 2696 55462 2726 55514
rect 2726 55462 2738 55514
rect 2738 55462 2752 55514
rect 2776 55462 2790 55514
rect 2790 55462 2802 55514
rect 2802 55462 2832 55514
rect 2856 55462 2866 55514
rect 2866 55462 2912 55514
rect 2616 55460 2672 55462
rect 2696 55460 2752 55462
rect 2776 55460 2832 55462
rect 2856 55460 2912 55462
rect 7616 55514 7672 55516
rect 7696 55514 7752 55516
rect 7776 55514 7832 55516
rect 7856 55514 7912 55516
rect 7616 55462 7662 55514
rect 7662 55462 7672 55514
rect 7696 55462 7726 55514
rect 7726 55462 7738 55514
rect 7738 55462 7752 55514
rect 7776 55462 7790 55514
rect 7790 55462 7802 55514
rect 7802 55462 7832 55514
rect 7856 55462 7866 55514
rect 7866 55462 7912 55514
rect 7616 55460 7672 55462
rect 7696 55460 7752 55462
rect 7776 55460 7832 55462
rect 7856 55460 7912 55462
rect 12616 55514 12672 55516
rect 12696 55514 12752 55516
rect 12776 55514 12832 55516
rect 12856 55514 12912 55516
rect 12616 55462 12662 55514
rect 12662 55462 12672 55514
rect 12696 55462 12726 55514
rect 12726 55462 12738 55514
rect 12738 55462 12752 55514
rect 12776 55462 12790 55514
rect 12790 55462 12802 55514
rect 12802 55462 12832 55514
rect 12856 55462 12866 55514
rect 12866 55462 12912 55514
rect 12616 55460 12672 55462
rect 12696 55460 12752 55462
rect 12776 55460 12832 55462
rect 12856 55460 12912 55462
rect 17616 55514 17672 55516
rect 17696 55514 17752 55516
rect 17776 55514 17832 55516
rect 17856 55514 17912 55516
rect 17616 55462 17662 55514
rect 17662 55462 17672 55514
rect 17696 55462 17726 55514
rect 17726 55462 17738 55514
rect 17738 55462 17752 55514
rect 17776 55462 17790 55514
rect 17790 55462 17802 55514
rect 17802 55462 17832 55514
rect 17856 55462 17866 55514
rect 17866 55462 17912 55514
rect 17616 55460 17672 55462
rect 17696 55460 17752 55462
rect 17776 55460 17832 55462
rect 17856 55460 17912 55462
rect 22616 55514 22672 55516
rect 22696 55514 22752 55516
rect 22776 55514 22832 55516
rect 22856 55514 22912 55516
rect 22616 55462 22662 55514
rect 22662 55462 22672 55514
rect 22696 55462 22726 55514
rect 22726 55462 22738 55514
rect 22738 55462 22752 55514
rect 22776 55462 22790 55514
rect 22790 55462 22802 55514
rect 22802 55462 22832 55514
rect 22856 55462 22866 55514
rect 22866 55462 22912 55514
rect 22616 55460 22672 55462
rect 22696 55460 22752 55462
rect 22776 55460 22832 55462
rect 22856 55460 22912 55462
rect 27616 55514 27672 55516
rect 27696 55514 27752 55516
rect 27776 55514 27832 55516
rect 27856 55514 27912 55516
rect 27616 55462 27662 55514
rect 27662 55462 27672 55514
rect 27696 55462 27726 55514
rect 27726 55462 27738 55514
rect 27738 55462 27752 55514
rect 27776 55462 27790 55514
rect 27790 55462 27802 55514
rect 27802 55462 27832 55514
rect 27856 55462 27866 55514
rect 27866 55462 27912 55514
rect 27616 55460 27672 55462
rect 27696 55460 27752 55462
rect 27776 55460 27832 55462
rect 27856 55460 27912 55462
rect 32616 55514 32672 55516
rect 32696 55514 32752 55516
rect 32776 55514 32832 55516
rect 32856 55514 32912 55516
rect 32616 55462 32662 55514
rect 32662 55462 32672 55514
rect 32696 55462 32726 55514
rect 32726 55462 32738 55514
rect 32738 55462 32752 55514
rect 32776 55462 32790 55514
rect 32790 55462 32802 55514
rect 32802 55462 32832 55514
rect 32856 55462 32866 55514
rect 32866 55462 32912 55514
rect 32616 55460 32672 55462
rect 32696 55460 32752 55462
rect 32776 55460 32832 55462
rect 32856 55460 32912 55462
rect 37616 55514 37672 55516
rect 37696 55514 37752 55516
rect 37776 55514 37832 55516
rect 37856 55514 37912 55516
rect 37616 55462 37662 55514
rect 37662 55462 37672 55514
rect 37696 55462 37726 55514
rect 37726 55462 37738 55514
rect 37738 55462 37752 55514
rect 37776 55462 37790 55514
rect 37790 55462 37802 55514
rect 37802 55462 37832 55514
rect 37856 55462 37866 55514
rect 37866 55462 37912 55514
rect 37616 55460 37672 55462
rect 37696 55460 37752 55462
rect 37776 55460 37832 55462
rect 37856 55460 37912 55462
rect 42616 55514 42672 55516
rect 42696 55514 42752 55516
rect 42776 55514 42832 55516
rect 42856 55514 42912 55516
rect 42616 55462 42662 55514
rect 42662 55462 42672 55514
rect 42696 55462 42726 55514
rect 42726 55462 42738 55514
rect 42738 55462 42752 55514
rect 42776 55462 42790 55514
rect 42790 55462 42802 55514
rect 42802 55462 42832 55514
rect 42856 55462 42866 55514
rect 42866 55462 42912 55514
rect 42616 55460 42672 55462
rect 42696 55460 42752 55462
rect 42776 55460 42832 55462
rect 42856 55460 42912 55462
rect 47616 55514 47672 55516
rect 47696 55514 47752 55516
rect 47776 55514 47832 55516
rect 47856 55514 47912 55516
rect 47616 55462 47662 55514
rect 47662 55462 47672 55514
rect 47696 55462 47726 55514
rect 47726 55462 47738 55514
rect 47738 55462 47752 55514
rect 47776 55462 47790 55514
rect 47790 55462 47802 55514
rect 47802 55462 47832 55514
rect 47856 55462 47866 55514
rect 47866 55462 47912 55514
rect 47616 55460 47672 55462
rect 47696 55460 47752 55462
rect 47776 55460 47832 55462
rect 47856 55460 47912 55462
rect 52616 55514 52672 55516
rect 52696 55514 52752 55516
rect 52776 55514 52832 55516
rect 52856 55514 52912 55516
rect 52616 55462 52662 55514
rect 52662 55462 52672 55514
rect 52696 55462 52726 55514
rect 52726 55462 52738 55514
rect 52738 55462 52752 55514
rect 52776 55462 52790 55514
rect 52790 55462 52802 55514
rect 52802 55462 52832 55514
rect 52856 55462 52866 55514
rect 52866 55462 52912 55514
rect 52616 55460 52672 55462
rect 52696 55460 52752 55462
rect 52776 55460 52832 55462
rect 52856 55460 52912 55462
rect 57616 55514 57672 55516
rect 57696 55514 57752 55516
rect 57776 55514 57832 55516
rect 57856 55514 57912 55516
rect 57616 55462 57662 55514
rect 57662 55462 57672 55514
rect 57696 55462 57726 55514
rect 57726 55462 57738 55514
rect 57738 55462 57752 55514
rect 57776 55462 57790 55514
rect 57790 55462 57802 55514
rect 57802 55462 57832 55514
rect 57856 55462 57866 55514
rect 57866 55462 57912 55514
rect 57616 55460 57672 55462
rect 57696 55460 57752 55462
rect 57776 55460 57832 55462
rect 57856 55460 57912 55462
rect 1956 54970 2012 54972
rect 2036 54970 2092 54972
rect 2116 54970 2172 54972
rect 2196 54970 2252 54972
rect 1956 54918 2002 54970
rect 2002 54918 2012 54970
rect 2036 54918 2066 54970
rect 2066 54918 2078 54970
rect 2078 54918 2092 54970
rect 2116 54918 2130 54970
rect 2130 54918 2142 54970
rect 2142 54918 2172 54970
rect 2196 54918 2206 54970
rect 2206 54918 2252 54970
rect 1956 54916 2012 54918
rect 2036 54916 2092 54918
rect 2116 54916 2172 54918
rect 2196 54916 2252 54918
rect 6956 54970 7012 54972
rect 7036 54970 7092 54972
rect 7116 54970 7172 54972
rect 7196 54970 7252 54972
rect 6956 54918 7002 54970
rect 7002 54918 7012 54970
rect 7036 54918 7066 54970
rect 7066 54918 7078 54970
rect 7078 54918 7092 54970
rect 7116 54918 7130 54970
rect 7130 54918 7142 54970
rect 7142 54918 7172 54970
rect 7196 54918 7206 54970
rect 7206 54918 7252 54970
rect 6956 54916 7012 54918
rect 7036 54916 7092 54918
rect 7116 54916 7172 54918
rect 7196 54916 7252 54918
rect 11956 54970 12012 54972
rect 12036 54970 12092 54972
rect 12116 54970 12172 54972
rect 12196 54970 12252 54972
rect 11956 54918 12002 54970
rect 12002 54918 12012 54970
rect 12036 54918 12066 54970
rect 12066 54918 12078 54970
rect 12078 54918 12092 54970
rect 12116 54918 12130 54970
rect 12130 54918 12142 54970
rect 12142 54918 12172 54970
rect 12196 54918 12206 54970
rect 12206 54918 12252 54970
rect 11956 54916 12012 54918
rect 12036 54916 12092 54918
rect 12116 54916 12172 54918
rect 12196 54916 12252 54918
rect 16956 54970 17012 54972
rect 17036 54970 17092 54972
rect 17116 54970 17172 54972
rect 17196 54970 17252 54972
rect 16956 54918 17002 54970
rect 17002 54918 17012 54970
rect 17036 54918 17066 54970
rect 17066 54918 17078 54970
rect 17078 54918 17092 54970
rect 17116 54918 17130 54970
rect 17130 54918 17142 54970
rect 17142 54918 17172 54970
rect 17196 54918 17206 54970
rect 17206 54918 17252 54970
rect 16956 54916 17012 54918
rect 17036 54916 17092 54918
rect 17116 54916 17172 54918
rect 17196 54916 17252 54918
rect 21956 54970 22012 54972
rect 22036 54970 22092 54972
rect 22116 54970 22172 54972
rect 22196 54970 22252 54972
rect 21956 54918 22002 54970
rect 22002 54918 22012 54970
rect 22036 54918 22066 54970
rect 22066 54918 22078 54970
rect 22078 54918 22092 54970
rect 22116 54918 22130 54970
rect 22130 54918 22142 54970
rect 22142 54918 22172 54970
rect 22196 54918 22206 54970
rect 22206 54918 22252 54970
rect 21956 54916 22012 54918
rect 22036 54916 22092 54918
rect 22116 54916 22172 54918
rect 22196 54916 22252 54918
rect 26956 54970 27012 54972
rect 27036 54970 27092 54972
rect 27116 54970 27172 54972
rect 27196 54970 27252 54972
rect 26956 54918 27002 54970
rect 27002 54918 27012 54970
rect 27036 54918 27066 54970
rect 27066 54918 27078 54970
rect 27078 54918 27092 54970
rect 27116 54918 27130 54970
rect 27130 54918 27142 54970
rect 27142 54918 27172 54970
rect 27196 54918 27206 54970
rect 27206 54918 27252 54970
rect 26956 54916 27012 54918
rect 27036 54916 27092 54918
rect 27116 54916 27172 54918
rect 27196 54916 27252 54918
rect 31956 54970 32012 54972
rect 32036 54970 32092 54972
rect 32116 54970 32172 54972
rect 32196 54970 32252 54972
rect 31956 54918 32002 54970
rect 32002 54918 32012 54970
rect 32036 54918 32066 54970
rect 32066 54918 32078 54970
rect 32078 54918 32092 54970
rect 32116 54918 32130 54970
rect 32130 54918 32142 54970
rect 32142 54918 32172 54970
rect 32196 54918 32206 54970
rect 32206 54918 32252 54970
rect 31956 54916 32012 54918
rect 32036 54916 32092 54918
rect 32116 54916 32172 54918
rect 32196 54916 32252 54918
rect 36956 54970 37012 54972
rect 37036 54970 37092 54972
rect 37116 54970 37172 54972
rect 37196 54970 37252 54972
rect 36956 54918 37002 54970
rect 37002 54918 37012 54970
rect 37036 54918 37066 54970
rect 37066 54918 37078 54970
rect 37078 54918 37092 54970
rect 37116 54918 37130 54970
rect 37130 54918 37142 54970
rect 37142 54918 37172 54970
rect 37196 54918 37206 54970
rect 37206 54918 37252 54970
rect 36956 54916 37012 54918
rect 37036 54916 37092 54918
rect 37116 54916 37172 54918
rect 37196 54916 37252 54918
rect 41956 54970 42012 54972
rect 42036 54970 42092 54972
rect 42116 54970 42172 54972
rect 42196 54970 42252 54972
rect 41956 54918 42002 54970
rect 42002 54918 42012 54970
rect 42036 54918 42066 54970
rect 42066 54918 42078 54970
rect 42078 54918 42092 54970
rect 42116 54918 42130 54970
rect 42130 54918 42142 54970
rect 42142 54918 42172 54970
rect 42196 54918 42206 54970
rect 42206 54918 42252 54970
rect 41956 54916 42012 54918
rect 42036 54916 42092 54918
rect 42116 54916 42172 54918
rect 42196 54916 42252 54918
rect 46956 54970 47012 54972
rect 47036 54970 47092 54972
rect 47116 54970 47172 54972
rect 47196 54970 47252 54972
rect 46956 54918 47002 54970
rect 47002 54918 47012 54970
rect 47036 54918 47066 54970
rect 47066 54918 47078 54970
rect 47078 54918 47092 54970
rect 47116 54918 47130 54970
rect 47130 54918 47142 54970
rect 47142 54918 47172 54970
rect 47196 54918 47206 54970
rect 47206 54918 47252 54970
rect 46956 54916 47012 54918
rect 47036 54916 47092 54918
rect 47116 54916 47172 54918
rect 47196 54916 47252 54918
rect 51956 54970 52012 54972
rect 52036 54970 52092 54972
rect 52116 54970 52172 54972
rect 52196 54970 52252 54972
rect 51956 54918 52002 54970
rect 52002 54918 52012 54970
rect 52036 54918 52066 54970
rect 52066 54918 52078 54970
rect 52078 54918 52092 54970
rect 52116 54918 52130 54970
rect 52130 54918 52142 54970
rect 52142 54918 52172 54970
rect 52196 54918 52206 54970
rect 52206 54918 52252 54970
rect 51956 54916 52012 54918
rect 52036 54916 52092 54918
rect 52116 54916 52172 54918
rect 52196 54916 52252 54918
rect 56956 54970 57012 54972
rect 57036 54970 57092 54972
rect 57116 54970 57172 54972
rect 57196 54970 57252 54972
rect 56956 54918 57002 54970
rect 57002 54918 57012 54970
rect 57036 54918 57066 54970
rect 57066 54918 57078 54970
rect 57078 54918 57092 54970
rect 57116 54918 57130 54970
rect 57130 54918 57142 54970
rect 57142 54918 57172 54970
rect 57196 54918 57206 54970
rect 57206 54918 57252 54970
rect 56956 54916 57012 54918
rect 57036 54916 57092 54918
rect 57116 54916 57172 54918
rect 57196 54916 57252 54918
rect 58530 54712 58586 54768
rect 2616 54426 2672 54428
rect 2696 54426 2752 54428
rect 2776 54426 2832 54428
rect 2856 54426 2912 54428
rect 2616 54374 2662 54426
rect 2662 54374 2672 54426
rect 2696 54374 2726 54426
rect 2726 54374 2738 54426
rect 2738 54374 2752 54426
rect 2776 54374 2790 54426
rect 2790 54374 2802 54426
rect 2802 54374 2832 54426
rect 2856 54374 2866 54426
rect 2866 54374 2912 54426
rect 2616 54372 2672 54374
rect 2696 54372 2752 54374
rect 2776 54372 2832 54374
rect 2856 54372 2912 54374
rect 7616 54426 7672 54428
rect 7696 54426 7752 54428
rect 7776 54426 7832 54428
rect 7856 54426 7912 54428
rect 7616 54374 7662 54426
rect 7662 54374 7672 54426
rect 7696 54374 7726 54426
rect 7726 54374 7738 54426
rect 7738 54374 7752 54426
rect 7776 54374 7790 54426
rect 7790 54374 7802 54426
rect 7802 54374 7832 54426
rect 7856 54374 7866 54426
rect 7866 54374 7912 54426
rect 7616 54372 7672 54374
rect 7696 54372 7752 54374
rect 7776 54372 7832 54374
rect 7856 54372 7912 54374
rect 12616 54426 12672 54428
rect 12696 54426 12752 54428
rect 12776 54426 12832 54428
rect 12856 54426 12912 54428
rect 12616 54374 12662 54426
rect 12662 54374 12672 54426
rect 12696 54374 12726 54426
rect 12726 54374 12738 54426
rect 12738 54374 12752 54426
rect 12776 54374 12790 54426
rect 12790 54374 12802 54426
rect 12802 54374 12832 54426
rect 12856 54374 12866 54426
rect 12866 54374 12912 54426
rect 12616 54372 12672 54374
rect 12696 54372 12752 54374
rect 12776 54372 12832 54374
rect 12856 54372 12912 54374
rect 17616 54426 17672 54428
rect 17696 54426 17752 54428
rect 17776 54426 17832 54428
rect 17856 54426 17912 54428
rect 17616 54374 17662 54426
rect 17662 54374 17672 54426
rect 17696 54374 17726 54426
rect 17726 54374 17738 54426
rect 17738 54374 17752 54426
rect 17776 54374 17790 54426
rect 17790 54374 17802 54426
rect 17802 54374 17832 54426
rect 17856 54374 17866 54426
rect 17866 54374 17912 54426
rect 17616 54372 17672 54374
rect 17696 54372 17752 54374
rect 17776 54372 17832 54374
rect 17856 54372 17912 54374
rect 22616 54426 22672 54428
rect 22696 54426 22752 54428
rect 22776 54426 22832 54428
rect 22856 54426 22912 54428
rect 22616 54374 22662 54426
rect 22662 54374 22672 54426
rect 22696 54374 22726 54426
rect 22726 54374 22738 54426
rect 22738 54374 22752 54426
rect 22776 54374 22790 54426
rect 22790 54374 22802 54426
rect 22802 54374 22832 54426
rect 22856 54374 22866 54426
rect 22866 54374 22912 54426
rect 22616 54372 22672 54374
rect 22696 54372 22752 54374
rect 22776 54372 22832 54374
rect 22856 54372 22912 54374
rect 27616 54426 27672 54428
rect 27696 54426 27752 54428
rect 27776 54426 27832 54428
rect 27856 54426 27912 54428
rect 27616 54374 27662 54426
rect 27662 54374 27672 54426
rect 27696 54374 27726 54426
rect 27726 54374 27738 54426
rect 27738 54374 27752 54426
rect 27776 54374 27790 54426
rect 27790 54374 27802 54426
rect 27802 54374 27832 54426
rect 27856 54374 27866 54426
rect 27866 54374 27912 54426
rect 27616 54372 27672 54374
rect 27696 54372 27752 54374
rect 27776 54372 27832 54374
rect 27856 54372 27912 54374
rect 32616 54426 32672 54428
rect 32696 54426 32752 54428
rect 32776 54426 32832 54428
rect 32856 54426 32912 54428
rect 32616 54374 32662 54426
rect 32662 54374 32672 54426
rect 32696 54374 32726 54426
rect 32726 54374 32738 54426
rect 32738 54374 32752 54426
rect 32776 54374 32790 54426
rect 32790 54374 32802 54426
rect 32802 54374 32832 54426
rect 32856 54374 32866 54426
rect 32866 54374 32912 54426
rect 32616 54372 32672 54374
rect 32696 54372 32752 54374
rect 32776 54372 32832 54374
rect 32856 54372 32912 54374
rect 37616 54426 37672 54428
rect 37696 54426 37752 54428
rect 37776 54426 37832 54428
rect 37856 54426 37912 54428
rect 37616 54374 37662 54426
rect 37662 54374 37672 54426
rect 37696 54374 37726 54426
rect 37726 54374 37738 54426
rect 37738 54374 37752 54426
rect 37776 54374 37790 54426
rect 37790 54374 37802 54426
rect 37802 54374 37832 54426
rect 37856 54374 37866 54426
rect 37866 54374 37912 54426
rect 37616 54372 37672 54374
rect 37696 54372 37752 54374
rect 37776 54372 37832 54374
rect 37856 54372 37912 54374
rect 42616 54426 42672 54428
rect 42696 54426 42752 54428
rect 42776 54426 42832 54428
rect 42856 54426 42912 54428
rect 42616 54374 42662 54426
rect 42662 54374 42672 54426
rect 42696 54374 42726 54426
rect 42726 54374 42738 54426
rect 42738 54374 42752 54426
rect 42776 54374 42790 54426
rect 42790 54374 42802 54426
rect 42802 54374 42832 54426
rect 42856 54374 42866 54426
rect 42866 54374 42912 54426
rect 42616 54372 42672 54374
rect 42696 54372 42752 54374
rect 42776 54372 42832 54374
rect 42856 54372 42912 54374
rect 47616 54426 47672 54428
rect 47696 54426 47752 54428
rect 47776 54426 47832 54428
rect 47856 54426 47912 54428
rect 47616 54374 47662 54426
rect 47662 54374 47672 54426
rect 47696 54374 47726 54426
rect 47726 54374 47738 54426
rect 47738 54374 47752 54426
rect 47776 54374 47790 54426
rect 47790 54374 47802 54426
rect 47802 54374 47832 54426
rect 47856 54374 47866 54426
rect 47866 54374 47912 54426
rect 47616 54372 47672 54374
rect 47696 54372 47752 54374
rect 47776 54372 47832 54374
rect 47856 54372 47912 54374
rect 52616 54426 52672 54428
rect 52696 54426 52752 54428
rect 52776 54426 52832 54428
rect 52856 54426 52912 54428
rect 52616 54374 52662 54426
rect 52662 54374 52672 54426
rect 52696 54374 52726 54426
rect 52726 54374 52738 54426
rect 52738 54374 52752 54426
rect 52776 54374 52790 54426
rect 52790 54374 52802 54426
rect 52802 54374 52832 54426
rect 52856 54374 52866 54426
rect 52866 54374 52912 54426
rect 52616 54372 52672 54374
rect 52696 54372 52752 54374
rect 52776 54372 52832 54374
rect 52856 54372 52912 54374
rect 57616 54426 57672 54428
rect 57696 54426 57752 54428
rect 57776 54426 57832 54428
rect 57856 54426 57912 54428
rect 57616 54374 57662 54426
rect 57662 54374 57672 54426
rect 57696 54374 57726 54426
rect 57726 54374 57738 54426
rect 57738 54374 57752 54426
rect 57776 54374 57790 54426
rect 57790 54374 57802 54426
rect 57802 54374 57832 54426
rect 57856 54374 57866 54426
rect 57866 54374 57912 54426
rect 57616 54372 57672 54374
rect 57696 54372 57752 54374
rect 57776 54372 57832 54374
rect 57856 54372 57912 54374
rect 58530 53932 58532 53952
rect 58532 53932 58584 53952
rect 58584 53932 58586 53952
rect 58530 53896 58586 53932
rect 1956 53882 2012 53884
rect 2036 53882 2092 53884
rect 2116 53882 2172 53884
rect 2196 53882 2252 53884
rect 1956 53830 2002 53882
rect 2002 53830 2012 53882
rect 2036 53830 2066 53882
rect 2066 53830 2078 53882
rect 2078 53830 2092 53882
rect 2116 53830 2130 53882
rect 2130 53830 2142 53882
rect 2142 53830 2172 53882
rect 2196 53830 2206 53882
rect 2206 53830 2252 53882
rect 1956 53828 2012 53830
rect 2036 53828 2092 53830
rect 2116 53828 2172 53830
rect 2196 53828 2252 53830
rect 6956 53882 7012 53884
rect 7036 53882 7092 53884
rect 7116 53882 7172 53884
rect 7196 53882 7252 53884
rect 6956 53830 7002 53882
rect 7002 53830 7012 53882
rect 7036 53830 7066 53882
rect 7066 53830 7078 53882
rect 7078 53830 7092 53882
rect 7116 53830 7130 53882
rect 7130 53830 7142 53882
rect 7142 53830 7172 53882
rect 7196 53830 7206 53882
rect 7206 53830 7252 53882
rect 6956 53828 7012 53830
rect 7036 53828 7092 53830
rect 7116 53828 7172 53830
rect 7196 53828 7252 53830
rect 11956 53882 12012 53884
rect 12036 53882 12092 53884
rect 12116 53882 12172 53884
rect 12196 53882 12252 53884
rect 11956 53830 12002 53882
rect 12002 53830 12012 53882
rect 12036 53830 12066 53882
rect 12066 53830 12078 53882
rect 12078 53830 12092 53882
rect 12116 53830 12130 53882
rect 12130 53830 12142 53882
rect 12142 53830 12172 53882
rect 12196 53830 12206 53882
rect 12206 53830 12252 53882
rect 11956 53828 12012 53830
rect 12036 53828 12092 53830
rect 12116 53828 12172 53830
rect 12196 53828 12252 53830
rect 16956 53882 17012 53884
rect 17036 53882 17092 53884
rect 17116 53882 17172 53884
rect 17196 53882 17252 53884
rect 16956 53830 17002 53882
rect 17002 53830 17012 53882
rect 17036 53830 17066 53882
rect 17066 53830 17078 53882
rect 17078 53830 17092 53882
rect 17116 53830 17130 53882
rect 17130 53830 17142 53882
rect 17142 53830 17172 53882
rect 17196 53830 17206 53882
rect 17206 53830 17252 53882
rect 16956 53828 17012 53830
rect 17036 53828 17092 53830
rect 17116 53828 17172 53830
rect 17196 53828 17252 53830
rect 21956 53882 22012 53884
rect 22036 53882 22092 53884
rect 22116 53882 22172 53884
rect 22196 53882 22252 53884
rect 21956 53830 22002 53882
rect 22002 53830 22012 53882
rect 22036 53830 22066 53882
rect 22066 53830 22078 53882
rect 22078 53830 22092 53882
rect 22116 53830 22130 53882
rect 22130 53830 22142 53882
rect 22142 53830 22172 53882
rect 22196 53830 22206 53882
rect 22206 53830 22252 53882
rect 21956 53828 22012 53830
rect 22036 53828 22092 53830
rect 22116 53828 22172 53830
rect 22196 53828 22252 53830
rect 26956 53882 27012 53884
rect 27036 53882 27092 53884
rect 27116 53882 27172 53884
rect 27196 53882 27252 53884
rect 26956 53830 27002 53882
rect 27002 53830 27012 53882
rect 27036 53830 27066 53882
rect 27066 53830 27078 53882
rect 27078 53830 27092 53882
rect 27116 53830 27130 53882
rect 27130 53830 27142 53882
rect 27142 53830 27172 53882
rect 27196 53830 27206 53882
rect 27206 53830 27252 53882
rect 26956 53828 27012 53830
rect 27036 53828 27092 53830
rect 27116 53828 27172 53830
rect 27196 53828 27252 53830
rect 31956 53882 32012 53884
rect 32036 53882 32092 53884
rect 32116 53882 32172 53884
rect 32196 53882 32252 53884
rect 31956 53830 32002 53882
rect 32002 53830 32012 53882
rect 32036 53830 32066 53882
rect 32066 53830 32078 53882
rect 32078 53830 32092 53882
rect 32116 53830 32130 53882
rect 32130 53830 32142 53882
rect 32142 53830 32172 53882
rect 32196 53830 32206 53882
rect 32206 53830 32252 53882
rect 31956 53828 32012 53830
rect 32036 53828 32092 53830
rect 32116 53828 32172 53830
rect 32196 53828 32252 53830
rect 36956 53882 37012 53884
rect 37036 53882 37092 53884
rect 37116 53882 37172 53884
rect 37196 53882 37252 53884
rect 36956 53830 37002 53882
rect 37002 53830 37012 53882
rect 37036 53830 37066 53882
rect 37066 53830 37078 53882
rect 37078 53830 37092 53882
rect 37116 53830 37130 53882
rect 37130 53830 37142 53882
rect 37142 53830 37172 53882
rect 37196 53830 37206 53882
rect 37206 53830 37252 53882
rect 36956 53828 37012 53830
rect 37036 53828 37092 53830
rect 37116 53828 37172 53830
rect 37196 53828 37252 53830
rect 41956 53882 42012 53884
rect 42036 53882 42092 53884
rect 42116 53882 42172 53884
rect 42196 53882 42252 53884
rect 41956 53830 42002 53882
rect 42002 53830 42012 53882
rect 42036 53830 42066 53882
rect 42066 53830 42078 53882
rect 42078 53830 42092 53882
rect 42116 53830 42130 53882
rect 42130 53830 42142 53882
rect 42142 53830 42172 53882
rect 42196 53830 42206 53882
rect 42206 53830 42252 53882
rect 41956 53828 42012 53830
rect 42036 53828 42092 53830
rect 42116 53828 42172 53830
rect 42196 53828 42252 53830
rect 46956 53882 47012 53884
rect 47036 53882 47092 53884
rect 47116 53882 47172 53884
rect 47196 53882 47252 53884
rect 46956 53830 47002 53882
rect 47002 53830 47012 53882
rect 47036 53830 47066 53882
rect 47066 53830 47078 53882
rect 47078 53830 47092 53882
rect 47116 53830 47130 53882
rect 47130 53830 47142 53882
rect 47142 53830 47172 53882
rect 47196 53830 47206 53882
rect 47206 53830 47252 53882
rect 46956 53828 47012 53830
rect 47036 53828 47092 53830
rect 47116 53828 47172 53830
rect 47196 53828 47252 53830
rect 51956 53882 52012 53884
rect 52036 53882 52092 53884
rect 52116 53882 52172 53884
rect 52196 53882 52252 53884
rect 51956 53830 52002 53882
rect 52002 53830 52012 53882
rect 52036 53830 52066 53882
rect 52066 53830 52078 53882
rect 52078 53830 52092 53882
rect 52116 53830 52130 53882
rect 52130 53830 52142 53882
rect 52142 53830 52172 53882
rect 52196 53830 52206 53882
rect 52206 53830 52252 53882
rect 51956 53828 52012 53830
rect 52036 53828 52092 53830
rect 52116 53828 52172 53830
rect 52196 53828 52252 53830
rect 56956 53882 57012 53884
rect 57036 53882 57092 53884
rect 57116 53882 57172 53884
rect 57196 53882 57252 53884
rect 56956 53830 57002 53882
rect 57002 53830 57012 53882
rect 57036 53830 57066 53882
rect 57066 53830 57078 53882
rect 57078 53830 57092 53882
rect 57116 53830 57130 53882
rect 57130 53830 57142 53882
rect 57142 53830 57172 53882
rect 57196 53830 57206 53882
rect 57206 53830 57252 53882
rect 56956 53828 57012 53830
rect 57036 53828 57092 53830
rect 57116 53828 57172 53830
rect 57196 53828 57252 53830
rect 2616 53338 2672 53340
rect 2696 53338 2752 53340
rect 2776 53338 2832 53340
rect 2856 53338 2912 53340
rect 2616 53286 2662 53338
rect 2662 53286 2672 53338
rect 2696 53286 2726 53338
rect 2726 53286 2738 53338
rect 2738 53286 2752 53338
rect 2776 53286 2790 53338
rect 2790 53286 2802 53338
rect 2802 53286 2832 53338
rect 2856 53286 2866 53338
rect 2866 53286 2912 53338
rect 2616 53284 2672 53286
rect 2696 53284 2752 53286
rect 2776 53284 2832 53286
rect 2856 53284 2912 53286
rect 7616 53338 7672 53340
rect 7696 53338 7752 53340
rect 7776 53338 7832 53340
rect 7856 53338 7912 53340
rect 7616 53286 7662 53338
rect 7662 53286 7672 53338
rect 7696 53286 7726 53338
rect 7726 53286 7738 53338
rect 7738 53286 7752 53338
rect 7776 53286 7790 53338
rect 7790 53286 7802 53338
rect 7802 53286 7832 53338
rect 7856 53286 7866 53338
rect 7866 53286 7912 53338
rect 7616 53284 7672 53286
rect 7696 53284 7752 53286
rect 7776 53284 7832 53286
rect 7856 53284 7912 53286
rect 12616 53338 12672 53340
rect 12696 53338 12752 53340
rect 12776 53338 12832 53340
rect 12856 53338 12912 53340
rect 12616 53286 12662 53338
rect 12662 53286 12672 53338
rect 12696 53286 12726 53338
rect 12726 53286 12738 53338
rect 12738 53286 12752 53338
rect 12776 53286 12790 53338
rect 12790 53286 12802 53338
rect 12802 53286 12832 53338
rect 12856 53286 12866 53338
rect 12866 53286 12912 53338
rect 12616 53284 12672 53286
rect 12696 53284 12752 53286
rect 12776 53284 12832 53286
rect 12856 53284 12912 53286
rect 17616 53338 17672 53340
rect 17696 53338 17752 53340
rect 17776 53338 17832 53340
rect 17856 53338 17912 53340
rect 17616 53286 17662 53338
rect 17662 53286 17672 53338
rect 17696 53286 17726 53338
rect 17726 53286 17738 53338
rect 17738 53286 17752 53338
rect 17776 53286 17790 53338
rect 17790 53286 17802 53338
rect 17802 53286 17832 53338
rect 17856 53286 17866 53338
rect 17866 53286 17912 53338
rect 17616 53284 17672 53286
rect 17696 53284 17752 53286
rect 17776 53284 17832 53286
rect 17856 53284 17912 53286
rect 22616 53338 22672 53340
rect 22696 53338 22752 53340
rect 22776 53338 22832 53340
rect 22856 53338 22912 53340
rect 22616 53286 22662 53338
rect 22662 53286 22672 53338
rect 22696 53286 22726 53338
rect 22726 53286 22738 53338
rect 22738 53286 22752 53338
rect 22776 53286 22790 53338
rect 22790 53286 22802 53338
rect 22802 53286 22832 53338
rect 22856 53286 22866 53338
rect 22866 53286 22912 53338
rect 22616 53284 22672 53286
rect 22696 53284 22752 53286
rect 22776 53284 22832 53286
rect 22856 53284 22912 53286
rect 27616 53338 27672 53340
rect 27696 53338 27752 53340
rect 27776 53338 27832 53340
rect 27856 53338 27912 53340
rect 27616 53286 27662 53338
rect 27662 53286 27672 53338
rect 27696 53286 27726 53338
rect 27726 53286 27738 53338
rect 27738 53286 27752 53338
rect 27776 53286 27790 53338
rect 27790 53286 27802 53338
rect 27802 53286 27832 53338
rect 27856 53286 27866 53338
rect 27866 53286 27912 53338
rect 27616 53284 27672 53286
rect 27696 53284 27752 53286
rect 27776 53284 27832 53286
rect 27856 53284 27912 53286
rect 32616 53338 32672 53340
rect 32696 53338 32752 53340
rect 32776 53338 32832 53340
rect 32856 53338 32912 53340
rect 32616 53286 32662 53338
rect 32662 53286 32672 53338
rect 32696 53286 32726 53338
rect 32726 53286 32738 53338
rect 32738 53286 32752 53338
rect 32776 53286 32790 53338
rect 32790 53286 32802 53338
rect 32802 53286 32832 53338
rect 32856 53286 32866 53338
rect 32866 53286 32912 53338
rect 32616 53284 32672 53286
rect 32696 53284 32752 53286
rect 32776 53284 32832 53286
rect 32856 53284 32912 53286
rect 37616 53338 37672 53340
rect 37696 53338 37752 53340
rect 37776 53338 37832 53340
rect 37856 53338 37912 53340
rect 37616 53286 37662 53338
rect 37662 53286 37672 53338
rect 37696 53286 37726 53338
rect 37726 53286 37738 53338
rect 37738 53286 37752 53338
rect 37776 53286 37790 53338
rect 37790 53286 37802 53338
rect 37802 53286 37832 53338
rect 37856 53286 37866 53338
rect 37866 53286 37912 53338
rect 37616 53284 37672 53286
rect 37696 53284 37752 53286
rect 37776 53284 37832 53286
rect 37856 53284 37912 53286
rect 42616 53338 42672 53340
rect 42696 53338 42752 53340
rect 42776 53338 42832 53340
rect 42856 53338 42912 53340
rect 42616 53286 42662 53338
rect 42662 53286 42672 53338
rect 42696 53286 42726 53338
rect 42726 53286 42738 53338
rect 42738 53286 42752 53338
rect 42776 53286 42790 53338
rect 42790 53286 42802 53338
rect 42802 53286 42832 53338
rect 42856 53286 42866 53338
rect 42866 53286 42912 53338
rect 42616 53284 42672 53286
rect 42696 53284 42752 53286
rect 42776 53284 42832 53286
rect 42856 53284 42912 53286
rect 47616 53338 47672 53340
rect 47696 53338 47752 53340
rect 47776 53338 47832 53340
rect 47856 53338 47912 53340
rect 47616 53286 47662 53338
rect 47662 53286 47672 53338
rect 47696 53286 47726 53338
rect 47726 53286 47738 53338
rect 47738 53286 47752 53338
rect 47776 53286 47790 53338
rect 47790 53286 47802 53338
rect 47802 53286 47832 53338
rect 47856 53286 47866 53338
rect 47866 53286 47912 53338
rect 47616 53284 47672 53286
rect 47696 53284 47752 53286
rect 47776 53284 47832 53286
rect 47856 53284 47912 53286
rect 52616 53338 52672 53340
rect 52696 53338 52752 53340
rect 52776 53338 52832 53340
rect 52856 53338 52912 53340
rect 52616 53286 52662 53338
rect 52662 53286 52672 53338
rect 52696 53286 52726 53338
rect 52726 53286 52738 53338
rect 52738 53286 52752 53338
rect 52776 53286 52790 53338
rect 52790 53286 52802 53338
rect 52802 53286 52832 53338
rect 52856 53286 52866 53338
rect 52866 53286 52912 53338
rect 52616 53284 52672 53286
rect 52696 53284 52752 53286
rect 52776 53284 52832 53286
rect 52856 53284 52912 53286
rect 57616 53338 57672 53340
rect 57696 53338 57752 53340
rect 57776 53338 57832 53340
rect 57856 53338 57912 53340
rect 57616 53286 57662 53338
rect 57662 53286 57672 53338
rect 57696 53286 57726 53338
rect 57726 53286 57738 53338
rect 57738 53286 57752 53338
rect 57776 53286 57790 53338
rect 57790 53286 57802 53338
rect 57802 53286 57832 53338
rect 57856 53286 57866 53338
rect 57866 53286 57912 53338
rect 57616 53284 57672 53286
rect 57696 53284 57752 53286
rect 57776 53284 57832 53286
rect 57856 53284 57912 53286
rect 58530 53080 58586 53136
rect 1956 52794 2012 52796
rect 2036 52794 2092 52796
rect 2116 52794 2172 52796
rect 2196 52794 2252 52796
rect 1956 52742 2002 52794
rect 2002 52742 2012 52794
rect 2036 52742 2066 52794
rect 2066 52742 2078 52794
rect 2078 52742 2092 52794
rect 2116 52742 2130 52794
rect 2130 52742 2142 52794
rect 2142 52742 2172 52794
rect 2196 52742 2206 52794
rect 2206 52742 2252 52794
rect 1956 52740 2012 52742
rect 2036 52740 2092 52742
rect 2116 52740 2172 52742
rect 2196 52740 2252 52742
rect 6956 52794 7012 52796
rect 7036 52794 7092 52796
rect 7116 52794 7172 52796
rect 7196 52794 7252 52796
rect 6956 52742 7002 52794
rect 7002 52742 7012 52794
rect 7036 52742 7066 52794
rect 7066 52742 7078 52794
rect 7078 52742 7092 52794
rect 7116 52742 7130 52794
rect 7130 52742 7142 52794
rect 7142 52742 7172 52794
rect 7196 52742 7206 52794
rect 7206 52742 7252 52794
rect 6956 52740 7012 52742
rect 7036 52740 7092 52742
rect 7116 52740 7172 52742
rect 7196 52740 7252 52742
rect 11956 52794 12012 52796
rect 12036 52794 12092 52796
rect 12116 52794 12172 52796
rect 12196 52794 12252 52796
rect 11956 52742 12002 52794
rect 12002 52742 12012 52794
rect 12036 52742 12066 52794
rect 12066 52742 12078 52794
rect 12078 52742 12092 52794
rect 12116 52742 12130 52794
rect 12130 52742 12142 52794
rect 12142 52742 12172 52794
rect 12196 52742 12206 52794
rect 12206 52742 12252 52794
rect 11956 52740 12012 52742
rect 12036 52740 12092 52742
rect 12116 52740 12172 52742
rect 12196 52740 12252 52742
rect 16956 52794 17012 52796
rect 17036 52794 17092 52796
rect 17116 52794 17172 52796
rect 17196 52794 17252 52796
rect 16956 52742 17002 52794
rect 17002 52742 17012 52794
rect 17036 52742 17066 52794
rect 17066 52742 17078 52794
rect 17078 52742 17092 52794
rect 17116 52742 17130 52794
rect 17130 52742 17142 52794
rect 17142 52742 17172 52794
rect 17196 52742 17206 52794
rect 17206 52742 17252 52794
rect 16956 52740 17012 52742
rect 17036 52740 17092 52742
rect 17116 52740 17172 52742
rect 17196 52740 17252 52742
rect 21956 52794 22012 52796
rect 22036 52794 22092 52796
rect 22116 52794 22172 52796
rect 22196 52794 22252 52796
rect 21956 52742 22002 52794
rect 22002 52742 22012 52794
rect 22036 52742 22066 52794
rect 22066 52742 22078 52794
rect 22078 52742 22092 52794
rect 22116 52742 22130 52794
rect 22130 52742 22142 52794
rect 22142 52742 22172 52794
rect 22196 52742 22206 52794
rect 22206 52742 22252 52794
rect 21956 52740 22012 52742
rect 22036 52740 22092 52742
rect 22116 52740 22172 52742
rect 22196 52740 22252 52742
rect 26956 52794 27012 52796
rect 27036 52794 27092 52796
rect 27116 52794 27172 52796
rect 27196 52794 27252 52796
rect 26956 52742 27002 52794
rect 27002 52742 27012 52794
rect 27036 52742 27066 52794
rect 27066 52742 27078 52794
rect 27078 52742 27092 52794
rect 27116 52742 27130 52794
rect 27130 52742 27142 52794
rect 27142 52742 27172 52794
rect 27196 52742 27206 52794
rect 27206 52742 27252 52794
rect 26956 52740 27012 52742
rect 27036 52740 27092 52742
rect 27116 52740 27172 52742
rect 27196 52740 27252 52742
rect 31956 52794 32012 52796
rect 32036 52794 32092 52796
rect 32116 52794 32172 52796
rect 32196 52794 32252 52796
rect 31956 52742 32002 52794
rect 32002 52742 32012 52794
rect 32036 52742 32066 52794
rect 32066 52742 32078 52794
rect 32078 52742 32092 52794
rect 32116 52742 32130 52794
rect 32130 52742 32142 52794
rect 32142 52742 32172 52794
rect 32196 52742 32206 52794
rect 32206 52742 32252 52794
rect 31956 52740 32012 52742
rect 32036 52740 32092 52742
rect 32116 52740 32172 52742
rect 32196 52740 32252 52742
rect 36956 52794 37012 52796
rect 37036 52794 37092 52796
rect 37116 52794 37172 52796
rect 37196 52794 37252 52796
rect 36956 52742 37002 52794
rect 37002 52742 37012 52794
rect 37036 52742 37066 52794
rect 37066 52742 37078 52794
rect 37078 52742 37092 52794
rect 37116 52742 37130 52794
rect 37130 52742 37142 52794
rect 37142 52742 37172 52794
rect 37196 52742 37206 52794
rect 37206 52742 37252 52794
rect 36956 52740 37012 52742
rect 37036 52740 37092 52742
rect 37116 52740 37172 52742
rect 37196 52740 37252 52742
rect 41956 52794 42012 52796
rect 42036 52794 42092 52796
rect 42116 52794 42172 52796
rect 42196 52794 42252 52796
rect 41956 52742 42002 52794
rect 42002 52742 42012 52794
rect 42036 52742 42066 52794
rect 42066 52742 42078 52794
rect 42078 52742 42092 52794
rect 42116 52742 42130 52794
rect 42130 52742 42142 52794
rect 42142 52742 42172 52794
rect 42196 52742 42206 52794
rect 42206 52742 42252 52794
rect 41956 52740 42012 52742
rect 42036 52740 42092 52742
rect 42116 52740 42172 52742
rect 42196 52740 42252 52742
rect 46956 52794 47012 52796
rect 47036 52794 47092 52796
rect 47116 52794 47172 52796
rect 47196 52794 47252 52796
rect 46956 52742 47002 52794
rect 47002 52742 47012 52794
rect 47036 52742 47066 52794
rect 47066 52742 47078 52794
rect 47078 52742 47092 52794
rect 47116 52742 47130 52794
rect 47130 52742 47142 52794
rect 47142 52742 47172 52794
rect 47196 52742 47206 52794
rect 47206 52742 47252 52794
rect 46956 52740 47012 52742
rect 47036 52740 47092 52742
rect 47116 52740 47172 52742
rect 47196 52740 47252 52742
rect 51956 52794 52012 52796
rect 52036 52794 52092 52796
rect 52116 52794 52172 52796
rect 52196 52794 52252 52796
rect 51956 52742 52002 52794
rect 52002 52742 52012 52794
rect 52036 52742 52066 52794
rect 52066 52742 52078 52794
rect 52078 52742 52092 52794
rect 52116 52742 52130 52794
rect 52130 52742 52142 52794
rect 52142 52742 52172 52794
rect 52196 52742 52206 52794
rect 52206 52742 52252 52794
rect 51956 52740 52012 52742
rect 52036 52740 52092 52742
rect 52116 52740 52172 52742
rect 52196 52740 52252 52742
rect 56956 52794 57012 52796
rect 57036 52794 57092 52796
rect 57116 52794 57172 52796
rect 57196 52794 57252 52796
rect 56956 52742 57002 52794
rect 57002 52742 57012 52794
rect 57036 52742 57066 52794
rect 57066 52742 57078 52794
rect 57078 52742 57092 52794
rect 57116 52742 57130 52794
rect 57130 52742 57142 52794
rect 57142 52742 57172 52794
rect 57196 52742 57206 52794
rect 57206 52742 57252 52794
rect 56956 52740 57012 52742
rect 57036 52740 57092 52742
rect 57116 52740 57172 52742
rect 57196 52740 57252 52742
rect 58530 52264 58586 52320
rect 2616 52250 2672 52252
rect 2696 52250 2752 52252
rect 2776 52250 2832 52252
rect 2856 52250 2912 52252
rect 2616 52198 2662 52250
rect 2662 52198 2672 52250
rect 2696 52198 2726 52250
rect 2726 52198 2738 52250
rect 2738 52198 2752 52250
rect 2776 52198 2790 52250
rect 2790 52198 2802 52250
rect 2802 52198 2832 52250
rect 2856 52198 2866 52250
rect 2866 52198 2912 52250
rect 2616 52196 2672 52198
rect 2696 52196 2752 52198
rect 2776 52196 2832 52198
rect 2856 52196 2912 52198
rect 7616 52250 7672 52252
rect 7696 52250 7752 52252
rect 7776 52250 7832 52252
rect 7856 52250 7912 52252
rect 7616 52198 7662 52250
rect 7662 52198 7672 52250
rect 7696 52198 7726 52250
rect 7726 52198 7738 52250
rect 7738 52198 7752 52250
rect 7776 52198 7790 52250
rect 7790 52198 7802 52250
rect 7802 52198 7832 52250
rect 7856 52198 7866 52250
rect 7866 52198 7912 52250
rect 7616 52196 7672 52198
rect 7696 52196 7752 52198
rect 7776 52196 7832 52198
rect 7856 52196 7912 52198
rect 12616 52250 12672 52252
rect 12696 52250 12752 52252
rect 12776 52250 12832 52252
rect 12856 52250 12912 52252
rect 12616 52198 12662 52250
rect 12662 52198 12672 52250
rect 12696 52198 12726 52250
rect 12726 52198 12738 52250
rect 12738 52198 12752 52250
rect 12776 52198 12790 52250
rect 12790 52198 12802 52250
rect 12802 52198 12832 52250
rect 12856 52198 12866 52250
rect 12866 52198 12912 52250
rect 12616 52196 12672 52198
rect 12696 52196 12752 52198
rect 12776 52196 12832 52198
rect 12856 52196 12912 52198
rect 17616 52250 17672 52252
rect 17696 52250 17752 52252
rect 17776 52250 17832 52252
rect 17856 52250 17912 52252
rect 17616 52198 17662 52250
rect 17662 52198 17672 52250
rect 17696 52198 17726 52250
rect 17726 52198 17738 52250
rect 17738 52198 17752 52250
rect 17776 52198 17790 52250
rect 17790 52198 17802 52250
rect 17802 52198 17832 52250
rect 17856 52198 17866 52250
rect 17866 52198 17912 52250
rect 17616 52196 17672 52198
rect 17696 52196 17752 52198
rect 17776 52196 17832 52198
rect 17856 52196 17912 52198
rect 22616 52250 22672 52252
rect 22696 52250 22752 52252
rect 22776 52250 22832 52252
rect 22856 52250 22912 52252
rect 22616 52198 22662 52250
rect 22662 52198 22672 52250
rect 22696 52198 22726 52250
rect 22726 52198 22738 52250
rect 22738 52198 22752 52250
rect 22776 52198 22790 52250
rect 22790 52198 22802 52250
rect 22802 52198 22832 52250
rect 22856 52198 22866 52250
rect 22866 52198 22912 52250
rect 22616 52196 22672 52198
rect 22696 52196 22752 52198
rect 22776 52196 22832 52198
rect 22856 52196 22912 52198
rect 27616 52250 27672 52252
rect 27696 52250 27752 52252
rect 27776 52250 27832 52252
rect 27856 52250 27912 52252
rect 27616 52198 27662 52250
rect 27662 52198 27672 52250
rect 27696 52198 27726 52250
rect 27726 52198 27738 52250
rect 27738 52198 27752 52250
rect 27776 52198 27790 52250
rect 27790 52198 27802 52250
rect 27802 52198 27832 52250
rect 27856 52198 27866 52250
rect 27866 52198 27912 52250
rect 27616 52196 27672 52198
rect 27696 52196 27752 52198
rect 27776 52196 27832 52198
rect 27856 52196 27912 52198
rect 32616 52250 32672 52252
rect 32696 52250 32752 52252
rect 32776 52250 32832 52252
rect 32856 52250 32912 52252
rect 32616 52198 32662 52250
rect 32662 52198 32672 52250
rect 32696 52198 32726 52250
rect 32726 52198 32738 52250
rect 32738 52198 32752 52250
rect 32776 52198 32790 52250
rect 32790 52198 32802 52250
rect 32802 52198 32832 52250
rect 32856 52198 32866 52250
rect 32866 52198 32912 52250
rect 32616 52196 32672 52198
rect 32696 52196 32752 52198
rect 32776 52196 32832 52198
rect 32856 52196 32912 52198
rect 37616 52250 37672 52252
rect 37696 52250 37752 52252
rect 37776 52250 37832 52252
rect 37856 52250 37912 52252
rect 37616 52198 37662 52250
rect 37662 52198 37672 52250
rect 37696 52198 37726 52250
rect 37726 52198 37738 52250
rect 37738 52198 37752 52250
rect 37776 52198 37790 52250
rect 37790 52198 37802 52250
rect 37802 52198 37832 52250
rect 37856 52198 37866 52250
rect 37866 52198 37912 52250
rect 37616 52196 37672 52198
rect 37696 52196 37752 52198
rect 37776 52196 37832 52198
rect 37856 52196 37912 52198
rect 42616 52250 42672 52252
rect 42696 52250 42752 52252
rect 42776 52250 42832 52252
rect 42856 52250 42912 52252
rect 42616 52198 42662 52250
rect 42662 52198 42672 52250
rect 42696 52198 42726 52250
rect 42726 52198 42738 52250
rect 42738 52198 42752 52250
rect 42776 52198 42790 52250
rect 42790 52198 42802 52250
rect 42802 52198 42832 52250
rect 42856 52198 42866 52250
rect 42866 52198 42912 52250
rect 42616 52196 42672 52198
rect 42696 52196 42752 52198
rect 42776 52196 42832 52198
rect 42856 52196 42912 52198
rect 47616 52250 47672 52252
rect 47696 52250 47752 52252
rect 47776 52250 47832 52252
rect 47856 52250 47912 52252
rect 47616 52198 47662 52250
rect 47662 52198 47672 52250
rect 47696 52198 47726 52250
rect 47726 52198 47738 52250
rect 47738 52198 47752 52250
rect 47776 52198 47790 52250
rect 47790 52198 47802 52250
rect 47802 52198 47832 52250
rect 47856 52198 47866 52250
rect 47866 52198 47912 52250
rect 47616 52196 47672 52198
rect 47696 52196 47752 52198
rect 47776 52196 47832 52198
rect 47856 52196 47912 52198
rect 52616 52250 52672 52252
rect 52696 52250 52752 52252
rect 52776 52250 52832 52252
rect 52856 52250 52912 52252
rect 52616 52198 52662 52250
rect 52662 52198 52672 52250
rect 52696 52198 52726 52250
rect 52726 52198 52738 52250
rect 52738 52198 52752 52250
rect 52776 52198 52790 52250
rect 52790 52198 52802 52250
rect 52802 52198 52832 52250
rect 52856 52198 52866 52250
rect 52866 52198 52912 52250
rect 52616 52196 52672 52198
rect 52696 52196 52752 52198
rect 52776 52196 52832 52198
rect 52856 52196 52912 52198
rect 57616 52250 57672 52252
rect 57696 52250 57752 52252
rect 57776 52250 57832 52252
rect 57856 52250 57912 52252
rect 57616 52198 57662 52250
rect 57662 52198 57672 52250
rect 57696 52198 57726 52250
rect 57726 52198 57738 52250
rect 57738 52198 57752 52250
rect 57776 52198 57790 52250
rect 57790 52198 57802 52250
rect 57802 52198 57832 52250
rect 57856 52198 57866 52250
rect 57866 52198 57912 52250
rect 57616 52196 57672 52198
rect 57696 52196 57752 52198
rect 57776 52196 57832 52198
rect 57856 52196 57912 52198
rect 1956 51706 2012 51708
rect 2036 51706 2092 51708
rect 2116 51706 2172 51708
rect 2196 51706 2252 51708
rect 1956 51654 2002 51706
rect 2002 51654 2012 51706
rect 2036 51654 2066 51706
rect 2066 51654 2078 51706
rect 2078 51654 2092 51706
rect 2116 51654 2130 51706
rect 2130 51654 2142 51706
rect 2142 51654 2172 51706
rect 2196 51654 2206 51706
rect 2206 51654 2252 51706
rect 1956 51652 2012 51654
rect 2036 51652 2092 51654
rect 2116 51652 2172 51654
rect 2196 51652 2252 51654
rect 6956 51706 7012 51708
rect 7036 51706 7092 51708
rect 7116 51706 7172 51708
rect 7196 51706 7252 51708
rect 6956 51654 7002 51706
rect 7002 51654 7012 51706
rect 7036 51654 7066 51706
rect 7066 51654 7078 51706
rect 7078 51654 7092 51706
rect 7116 51654 7130 51706
rect 7130 51654 7142 51706
rect 7142 51654 7172 51706
rect 7196 51654 7206 51706
rect 7206 51654 7252 51706
rect 6956 51652 7012 51654
rect 7036 51652 7092 51654
rect 7116 51652 7172 51654
rect 7196 51652 7252 51654
rect 11956 51706 12012 51708
rect 12036 51706 12092 51708
rect 12116 51706 12172 51708
rect 12196 51706 12252 51708
rect 11956 51654 12002 51706
rect 12002 51654 12012 51706
rect 12036 51654 12066 51706
rect 12066 51654 12078 51706
rect 12078 51654 12092 51706
rect 12116 51654 12130 51706
rect 12130 51654 12142 51706
rect 12142 51654 12172 51706
rect 12196 51654 12206 51706
rect 12206 51654 12252 51706
rect 11956 51652 12012 51654
rect 12036 51652 12092 51654
rect 12116 51652 12172 51654
rect 12196 51652 12252 51654
rect 16956 51706 17012 51708
rect 17036 51706 17092 51708
rect 17116 51706 17172 51708
rect 17196 51706 17252 51708
rect 16956 51654 17002 51706
rect 17002 51654 17012 51706
rect 17036 51654 17066 51706
rect 17066 51654 17078 51706
rect 17078 51654 17092 51706
rect 17116 51654 17130 51706
rect 17130 51654 17142 51706
rect 17142 51654 17172 51706
rect 17196 51654 17206 51706
rect 17206 51654 17252 51706
rect 16956 51652 17012 51654
rect 17036 51652 17092 51654
rect 17116 51652 17172 51654
rect 17196 51652 17252 51654
rect 21956 51706 22012 51708
rect 22036 51706 22092 51708
rect 22116 51706 22172 51708
rect 22196 51706 22252 51708
rect 21956 51654 22002 51706
rect 22002 51654 22012 51706
rect 22036 51654 22066 51706
rect 22066 51654 22078 51706
rect 22078 51654 22092 51706
rect 22116 51654 22130 51706
rect 22130 51654 22142 51706
rect 22142 51654 22172 51706
rect 22196 51654 22206 51706
rect 22206 51654 22252 51706
rect 21956 51652 22012 51654
rect 22036 51652 22092 51654
rect 22116 51652 22172 51654
rect 22196 51652 22252 51654
rect 26956 51706 27012 51708
rect 27036 51706 27092 51708
rect 27116 51706 27172 51708
rect 27196 51706 27252 51708
rect 26956 51654 27002 51706
rect 27002 51654 27012 51706
rect 27036 51654 27066 51706
rect 27066 51654 27078 51706
rect 27078 51654 27092 51706
rect 27116 51654 27130 51706
rect 27130 51654 27142 51706
rect 27142 51654 27172 51706
rect 27196 51654 27206 51706
rect 27206 51654 27252 51706
rect 26956 51652 27012 51654
rect 27036 51652 27092 51654
rect 27116 51652 27172 51654
rect 27196 51652 27252 51654
rect 31956 51706 32012 51708
rect 32036 51706 32092 51708
rect 32116 51706 32172 51708
rect 32196 51706 32252 51708
rect 31956 51654 32002 51706
rect 32002 51654 32012 51706
rect 32036 51654 32066 51706
rect 32066 51654 32078 51706
rect 32078 51654 32092 51706
rect 32116 51654 32130 51706
rect 32130 51654 32142 51706
rect 32142 51654 32172 51706
rect 32196 51654 32206 51706
rect 32206 51654 32252 51706
rect 31956 51652 32012 51654
rect 32036 51652 32092 51654
rect 32116 51652 32172 51654
rect 32196 51652 32252 51654
rect 36956 51706 37012 51708
rect 37036 51706 37092 51708
rect 37116 51706 37172 51708
rect 37196 51706 37252 51708
rect 36956 51654 37002 51706
rect 37002 51654 37012 51706
rect 37036 51654 37066 51706
rect 37066 51654 37078 51706
rect 37078 51654 37092 51706
rect 37116 51654 37130 51706
rect 37130 51654 37142 51706
rect 37142 51654 37172 51706
rect 37196 51654 37206 51706
rect 37206 51654 37252 51706
rect 36956 51652 37012 51654
rect 37036 51652 37092 51654
rect 37116 51652 37172 51654
rect 37196 51652 37252 51654
rect 41956 51706 42012 51708
rect 42036 51706 42092 51708
rect 42116 51706 42172 51708
rect 42196 51706 42252 51708
rect 41956 51654 42002 51706
rect 42002 51654 42012 51706
rect 42036 51654 42066 51706
rect 42066 51654 42078 51706
rect 42078 51654 42092 51706
rect 42116 51654 42130 51706
rect 42130 51654 42142 51706
rect 42142 51654 42172 51706
rect 42196 51654 42206 51706
rect 42206 51654 42252 51706
rect 41956 51652 42012 51654
rect 42036 51652 42092 51654
rect 42116 51652 42172 51654
rect 42196 51652 42252 51654
rect 46956 51706 47012 51708
rect 47036 51706 47092 51708
rect 47116 51706 47172 51708
rect 47196 51706 47252 51708
rect 46956 51654 47002 51706
rect 47002 51654 47012 51706
rect 47036 51654 47066 51706
rect 47066 51654 47078 51706
rect 47078 51654 47092 51706
rect 47116 51654 47130 51706
rect 47130 51654 47142 51706
rect 47142 51654 47172 51706
rect 47196 51654 47206 51706
rect 47206 51654 47252 51706
rect 46956 51652 47012 51654
rect 47036 51652 47092 51654
rect 47116 51652 47172 51654
rect 47196 51652 47252 51654
rect 51956 51706 52012 51708
rect 52036 51706 52092 51708
rect 52116 51706 52172 51708
rect 52196 51706 52252 51708
rect 51956 51654 52002 51706
rect 52002 51654 52012 51706
rect 52036 51654 52066 51706
rect 52066 51654 52078 51706
rect 52078 51654 52092 51706
rect 52116 51654 52130 51706
rect 52130 51654 52142 51706
rect 52142 51654 52172 51706
rect 52196 51654 52206 51706
rect 52206 51654 52252 51706
rect 51956 51652 52012 51654
rect 52036 51652 52092 51654
rect 52116 51652 52172 51654
rect 52196 51652 52252 51654
rect 56956 51706 57012 51708
rect 57036 51706 57092 51708
rect 57116 51706 57172 51708
rect 57196 51706 57252 51708
rect 56956 51654 57002 51706
rect 57002 51654 57012 51706
rect 57036 51654 57066 51706
rect 57066 51654 57078 51706
rect 57078 51654 57092 51706
rect 57116 51654 57130 51706
rect 57130 51654 57142 51706
rect 57142 51654 57172 51706
rect 57196 51654 57206 51706
rect 57206 51654 57252 51706
rect 56956 51652 57012 51654
rect 57036 51652 57092 51654
rect 57116 51652 57172 51654
rect 57196 51652 57252 51654
rect 58530 51448 58586 51504
rect 2616 51162 2672 51164
rect 2696 51162 2752 51164
rect 2776 51162 2832 51164
rect 2856 51162 2912 51164
rect 2616 51110 2662 51162
rect 2662 51110 2672 51162
rect 2696 51110 2726 51162
rect 2726 51110 2738 51162
rect 2738 51110 2752 51162
rect 2776 51110 2790 51162
rect 2790 51110 2802 51162
rect 2802 51110 2832 51162
rect 2856 51110 2866 51162
rect 2866 51110 2912 51162
rect 2616 51108 2672 51110
rect 2696 51108 2752 51110
rect 2776 51108 2832 51110
rect 2856 51108 2912 51110
rect 7616 51162 7672 51164
rect 7696 51162 7752 51164
rect 7776 51162 7832 51164
rect 7856 51162 7912 51164
rect 7616 51110 7662 51162
rect 7662 51110 7672 51162
rect 7696 51110 7726 51162
rect 7726 51110 7738 51162
rect 7738 51110 7752 51162
rect 7776 51110 7790 51162
rect 7790 51110 7802 51162
rect 7802 51110 7832 51162
rect 7856 51110 7866 51162
rect 7866 51110 7912 51162
rect 7616 51108 7672 51110
rect 7696 51108 7752 51110
rect 7776 51108 7832 51110
rect 7856 51108 7912 51110
rect 12616 51162 12672 51164
rect 12696 51162 12752 51164
rect 12776 51162 12832 51164
rect 12856 51162 12912 51164
rect 12616 51110 12662 51162
rect 12662 51110 12672 51162
rect 12696 51110 12726 51162
rect 12726 51110 12738 51162
rect 12738 51110 12752 51162
rect 12776 51110 12790 51162
rect 12790 51110 12802 51162
rect 12802 51110 12832 51162
rect 12856 51110 12866 51162
rect 12866 51110 12912 51162
rect 12616 51108 12672 51110
rect 12696 51108 12752 51110
rect 12776 51108 12832 51110
rect 12856 51108 12912 51110
rect 17616 51162 17672 51164
rect 17696 51162 17752 51164
rect 17776 51162 17832 51164
rect 17856 51162 17912 51164
rect 17616 51110 17662 51162
rect 17662 51110 17672 51162
rect 17696 51110 17726 51162
rect 17726 51110 17738 51162
rect 17738 51110 17752 51162
rect 17776 51110 17790 51162
rect 17790 51110 17802 51162
rect 17802 51110 17832 51162
rect 17856 51110 17866 51162
rect 17866 51110 17912 51162
rect 17616 51108 17672 51110
rect 17696 51108 17752 51110
rect 17776 51108 17832 51110
rect 17856 51108 17912 51110
rect 22616 51162 22672 51164
rect 22696 51162 22752 51164
rect 22776 51162 22832 51164
rect 22856 51162 22912 51164
rect 22616 51110 22662 51162
rect 22662 51110 22672 51162
rect 22696 51110 22726 51162
rect 22726 51110 22738 51162
rect 22738 51110 22752 51162
rect 22776 51110 22790 51162
rect 22790 51110 22802 51162
rect 22802 51110 22832 51162
rect 22856 51110 22866 51162
rect 22866 51110 22912 51162
rect 22616 51108 22672 51110
rect 22696 51108 22752 51110
rect 22776 51108 22832 51110
rect 22856 51108 22912 51110
rect 27616 51162 27672 51164
rect 27696 51162 27752 51164
rect 27776 51162 27832 51164
rect 27856 51162 27912 51164
rect 27616 51110 27662 51162
rect 27662 51110 27672 51162
rect 27696 51110 27726 51162
rect 27726 51110 27738 51162
rect 27738 51110 27752 51162
rect 27776 51110 27790 51162
rect 27790 51110 27802 51162
rect 27802 51110 27832 51162
rect 27856 51110 27866 51162
rect 27866 51110 27912 51162
rect 27616 51108 27672 51110
rect 27696 51108 27752 51110
rect 27776 51108 27832 51110
rect 27856 51108 27912 51110
rect 32616 51162 32672 51164
rect 32696 51162 32752 51164
rect 32776 51162 32832 51164
rect 32856 51162 32912 51164
rect 32616 51110 32662 51162
rect 32662 51110 32672 51162
rect 32696 51110 32726 51162
rect 32726 51110 32738 51162
rect 32738 51110 32752 51162
rect 32776 51110 32790 51162
rect 32790 51110 32802 51162
rect 32802 51110 32832 51162
rect 32856 51110 32866 51162
rect 32866 51110 32912 51162
rect 32616 51108 32672 51110
rect 32696 51108 32752 51110
rect 32776 51108 32832 51110
rect 32856 51108 32912 51110
rect 37616 51162 37672 51164
rect 37696 51162 37752 51164
rect 37776 51162 37832 51164
rect 37856 51162 37912 51164
rect 37616 51110 37662 51162
rect 37662 51110 37672 51162
rect 37696 51110 37726 51162
rect 37726 51110 37738 51162
rect 37738 51110 37752 51162
rect 37776 51110 37790 51162
rect 37790 51110 37802 51162
rect 37802 51110 37832 51162
rect 37856 51110 37866 51162
rect 37866 51110 37912 51162
rect 37616 51108 37672 51110
rect 37696 51108 37752 51110
rect 37776 51108 37832 51110
rect 37856 51108 37912 51110
rect 42616 51162 42672 51164
rect 42696 51162 42752 51164
rect 42776 51162 42832 51164
rect 42856 51162 42912 51164
rect 42616 51110 42662 51162
rect 42662 51110 42672 51162
rect 42696 51110 42726 51162
rect 42726 51110 42738 51162
rect 42738 51110 42752 51162
rect 42776 51110 42790 51162
rect 42790 51110 42802 51162
rect 42802 51110 42832 51162
rect 42856 51110 42866 51162
rect 42866 51110 42912 51162
rect 42616 51108 42672 51110
rect 42696 51108 42752 51110
rect 42776 51108 42832 51110
rect 42856 51108 42912 51110
rect 47616 51162 47672 51164
rect 47696 51162 47752 51164
rect 47776 51162 47832 51164
rect 47856 51162 47912 51164
rect 47616 51110 47662 51162
rect 47662 51110 47672 51162
rect 47696 51110 47726 51162
rect 47726 51110 47738 51162
rect 47738 51110 47752 51162
rect 47776 51110 47790 51162
rect 47790 51110 47802 51162
rect 47802 51110 47832 51162
rect 47856 51110 47866 51162
rect 47866 51110 47912 51162
rect 47616 51108 47672 51110
rect 47696 51108 47752 51110
rect 47776 51108 47832 51110
rect 47856 51108 47912 51110
rect 52616 51162 52672 51164
rect 52696 51162 52752 51164
rect 52776 51162 52832 51164
rect 52856 51162 52912 51164
rect 52616 51110 52662 51162
rect 52662 51110 52672 51162
rect 52696 51110 52726 51162
rect 52726 51110 52738 51162
rect 52738 51110 52752 51162
rect 52776 51110 52790 51162
rect 52790 51110 52802 51162
rect 52802 51110 52832 51162
rect 52856 51110 52866 51162
rect 52866 51110 52912 51162
rect 52616 51108 52672 51110
rect 52696 51108 52752 51110
rect 52776 51108 52832 51110
rect 52856 51108 52912 51110
rect 57616 51162 57672 51164
rect 57696 51162 57752 51164
rect 57776 51162 57832 51164
rect 57856 51162 57912 51164
rect 57616 51110 57662 51162
rect 57662 51110 57672 51162
rect 57696 51110 57726 51162
rect 57726 51110 57738 51162
rect 57738 51110 57752 51162
rect 57776 51110 57790 51162
rect 57790 51110 57802 51162
rect 57802 51110 57832 51162
rect 57856 51110 57866 51162
rect 57866 51110 57912 51162
rect 57616 51108 57672 51110
rect 57696 51108 57752 51110
rect 57776 51108 57832 51110
rect 57856 51108 57912 51110
rect 58530 50668 58532 50688
rect 58532 50668 58584 50688
rect 58584 50668 58586 50688
rect 58530 50632 58586 50668
rect 1956 50618 2012 50620
rect 2036 50618 2092 50620
rect 2116 50618 2172 50620
rect 2196 50618 2252 50620
rect 1956 50566 2002 50618
rect 2002 50566 2012 50618
rect 2036 50566 2066 50618
rect 2066 50566 2078 50618
rect 2078 50566 2092 50618
rect 2116 50566 2130 50618
rect 2130 50566 2142 50618
rect 2142 50566 2172 50618
rect 2196 50566 2206 50618
rect 2206 50566 2252 50618
rect 1956 50564 2012 50566
rect 2036 50564 2092 50566
rect 2116 50564 2172 50566
rect 2196 50564 2252 50566
rect 6956 50618 7012 50620
rect 7036 50618 7092 50620
rect 7116 50618 7172 50620
rect 7196 50618 7252 50620
rect 6956 50566 7002 50618
rect 7002 50566 7012 50618
rect 7036 50566 7066 50618
rect 7066 50566 7078 50618
rect 7078 50566 7092 50618
rect 7116 50566 7130 50618
rect 7130 50566 7142 50618
rect 7142 50566 7172 50618
rect 7196 50566 7206 50618
rect 7206 50566 7252 50618
rect 6956 50564 7012 50566
rect 7036 50564 7092 50566
rect 7116 50564 7172 50566
rect 7196 50564 7252 50566
rect 11956 50618 12012 50620
rect 12036 50618 12092 50620
rect 12116 50618 12172 50620
rect 12196 50618 12252 50620
rect 11956 50566 12002 50618
rect 12002 50566 12012 50618
rect 12036 50566 12066 50618
rect 12066 50566 12078 50618
rect 12078 50566 12092 50618
rect 12116 50566 12130 50618
rect 12130 50566 12142 50618
rect 12142 50566 12172 50618
rect 12196 50566 12206 50618
rect 12206 50566 12252 50618
rect 11956 50564 12012 50566
rect 12036 50564 12092 50566
rect 12116 50564 12172 50566
rect 12196 50564 12252 50566
rect 16956 50618 17012 50620
rect 17036 50618 17092 50620
rect 17116 50618 17172 50620
rect 17196 50618 17252 50620
rect 16956 50566 17002 50618
rect 17002 50566 17012 50618
rect 17036 50566 17066 50618
rect 17066 50566 17078 50618
rect 17078 50566 17092 50618
rect 17116 50566 17130 50618
rect 17130 50566 17142 50618
rect 17142 50566 17172 50618
rect 17196 50566 17206 50618
rect 17206 50566 17252 50618
rect 16956 50564 17012 50566
rect 17036 50564 17092 50566
rect 17116 50564 17172 50566
rect 17196 50564 17252 50566
rect 21956 50618 22012 50620
rect 22036 50618 22092 50620
rect 22116 50618 22172 50620
rect 22196 50618 22252 50620
rect 21956 50566 22002 50618
rect 22002 50566 22012 50618
rect 22036 50566 22066 50618
rect 22066 50566 22078 50618
rect 22078 50566 22092 50618
rect 22116 50566 22130 50618
rect 22130 50566 22142 50618
rect 22142 50566 22172 50618
rect 22196 50566 22206 50618
rect 22206 50566 22252 50618
rect 21956 50564 22012 50566
rect 22036 50564 22092 50566
rect 22116 50564 22172 50566
rect 22196 50564 22252 50566
rect 26956 50618 27012 50620
rect 27036 50618 27092 50620
rect 27116 50618 27172 50620
rect 27196 50618 27252 50620
rect 26956 50566 27002 50618
rect 27002 50566 27012 50618
rect 27036 50566 27066 50618
rect 27066 50566 27078 50618
rect 27078 50566 27092 50618
rect 27116 50566 27130 50618
rect 27130 50566 27142 50618
rect 27142 50566 27172 50618
rect 27196 50566 27206 50618
rect 27206 50566 27252 50618
rect 26956 50564 27012 50566
rect 27036 50564 27092 50566
rect 27116 50564 27172 50566
rect 27196 50564 27252 50566
rect 31956 50618 32012 50620
rect 32036 50618 32092 50620
rect 32116 50618 32172 50620
rect 32196 50618 32252 50620
rect 31956 50566 32002 50618
rect 32002 50566 32012 50618
rect 32036 50566 32066 50618
rect 32066 50566 32078 50618
rect 32078 50566 32092 50618
rect 32116 50566 32130 50618
rect 32130 50566 32142 50618
rect 32142 50566 32172 50618
rect 32196 50566 32206 50618
rect 32206 50566 32252 50618
rect 31956 50564 32012 50566
rect 32036 50564 32092 50566
rect 32116 50564 32172 50566
rect 32196 50564 32252 50566
rect 36956 50618 37012 50620
rect 37036 50618 37092 50620
rect 37116 50618 37172 50620
rect 37196 50618 37252 50620
rect 36956 50566 37002 50618
rect 37002 50566 37012 50618
rect 37036 50566 37066 50618
rect 37066 50566 37078 50618
rect 37078 50566 37092 50618
rect 37116 50566 37130 50618
rect 37130 50566 37142 50618
rect 37142 50566 37172 50618
rect 37196 50566 37206 50618
rect 37206 50566 37252 50618
rect 36956 50564 37012 50566
rect 37036 50564 37092 50566
rect 37116 50564 37172 50566
rect 37196 50564 37252 50566
rect 41956 50618 42012 50620
rect 42036 50618 42092 50620
rect 42116 50618 42172 50620
rect 42196 50618 42252 50620
rect 41956 50566 42002 50618
rect 42002 50566 42012 50618
rect 42036 50566 42066 50618
rect 42066 50566 42078 50618
rect 42078 50566 42092 50618
rect 42116 50566 42130 50618
rect 42130 50566 42142 50618
rect 42142 50566 42172 50618
rect 42196 50566 42206 50618
rect 42206 50566 42252 50618
rect 41956 50564 42012 50566
rect 42036 50564 42092 50566
rect 42116 50564 42172 50566
rect 42196 50564 42252 50566
rect 46956 50618 47012 50620
rect 47036 50618 47092 50620
rect 47116 50618 47172 50620
rect 47196 50618 47252 50620
rect 46956 50566 47002 50618
rect 47002 50566 47012 50618
rect 47036 50566 47066 50618
rect 47066 50566 47078 50618
rect 47078 50566 47092 50618
rect 47116 50566 47130 50618
rect 47130 50566 47142 50618
rect 47142 50566 47172 50618
rect 47196 50566 47206 50618
rect 47206 50566 47252 50618
rect 46956 50564 47012 50566
rect 47036 50564 47092 50566
rect 47116 50564 47172 50566
rect 47196 50564 47252 50566
rect 51956 50618 52012 50620
rect 52036 50618 52092 50620
rect 52116 50618 52172 50620
rect 52196 50618 52252 50620
rect 51956 50566 52002 50618
rect 52002 50566 52012 50618
rect 52036 50566 52066 50618
rect 52066 50566 52078 50618
rect 52078 50566 52092 50618
rect 52116 50566 52130 50618
rect 52130 50566 52142 50618
rect 52142 50566 52172 50618
rect 52196 50566 52206 50618
rect 52206 50566 52252 50618
rect 51956 50564 52012 50566
rect 52036 50564 52092 50566
rect 52116 50564 52172 50566
rect 52196 50564 52252 50566
rect 56956 50618 57012 50620
rect 57036 50618 57092 50620
rect 57116 50618 57172 50620
rect 57196 50618 57252 50620
rect 56956 50566 57002 50618
rect 57002 50566 57012 50618
rect 57036 50566 57066 50618
rect 57066 50566 57078 50618
rect 57078 50566 57092 50618
rect 57116 50566 57130 50618
rect 57130 50566 57142 50618
rect 57142 50566 57172 50618
rect 57196 50566 57206 50618
rect 57206 50566 57252 50618
rect 56956 50564 57012 50566
rect 57036 50564 57092 50566
rect 57116 50564 57172 50566
rect 57196 50564 57252 50566
rect 2616 50074 2672 50076
rect 2696 50074 2752 50076
rect 2776 50074 2832 50076
rect 2856 50074 2912 50076
rect 2616 50022 2662 50074
rect 2662 50022 2672 50074
rect 2696 50022 2726 50074
rect 2726 50022 2738 50074
rect 2738 50022 2752 50074
rect 2776 50022 2790 50074
rect 2790 50022 2802 50074
rect 2802 50022 2832 50074
rect 2856 50022 2866 50074
rect 2866 50022 2912 50074
rect 2616 50020 2672 50022
rect 2696 50020 2752 50022
rect 2776 50020 2832 50022
rect 2856 50020 2912 50022
rect 7616 50074 7672 50076
rect 7696 50074 7752 50076
rect 7776 50074 7832 50076
rect 7856 50074 7912 50076
rect 7616 50022 7662 50074
rect 7662 50022 7672 50074
rect 7696 50022 7726 50074
rect 7726 50022 7738 50074
rect 7738 50022 7752 50074
rect 7776 50022 7790 50074
rect 7790 50022 7802 50074
rect 7802 50022 7832 50074
rect 7856 50022 7866 50074
rect 7866 50022 7912 50074
rect 7616 50020 7672 50022
rect 7696 50020 7752 50022
rect 7776 50020 7832 50022
rect 7856 50020 7912 50022
rect 12616 50074 12672 50076
rect 12696 50074 12752 50076
rect 12776 50074 12832 50076
rect 12856 50074 12912 50076
rect 12616 50022 12662 50074
rect 12662 50022 12672 50074
rect 12696 50022 12726 50074
rect 12726 50022 12738 50074
rect 12738 50022 12752 50074
rect 12776 50022 12790 50074
rect 12790 50022 12802 50074
rect 12802 50022 12832 50074
rect 12856 50022 12866 50074
rect 12866 50022 12912 50074
rect 12616 50020 12672 50022
rect 12696 50020 12752 50022
rect 12776 50020 12832 50022
rect 12856 50020 12912 50022
rect 17616 50074 17672 50076
rect 17696 50074 17752 50076
rect 17776 50074 17832 50076
rect 17856 50074 17912 50076
rect 17616 50022 17662 50074
rect 17662 50022 17672 50074
rect 17696 50022 17726 50074
rect 17726 50022 17738 50074
rect 17738 50022 17752 50074
rect 17776 50022 17790 50074
rect 17790 50022 17802 50074
rect 17802 50022 17832 50074
rect 17856 50022 17866 50074
rect 17866 50022 17912 50074
rect 17616 50020 17672 50022
rect 17696 50020 17752 50022
rect 17776 50020 17832 50022
rect 17856 50020 17912 50022
rect 22616 50074 22672 50076
rect 22696 50074 22752 50076
rect 22776 50074 22832 50076
rect 22856 50074 22912 50076
rect 22616 50022 22662 50074
rect 22662 50022 22672 50074
rect 22696 50022 22726 50074
rect 22726 50022 22738 50074
rect 22738 50022 22752 50074
rect 22776 50022 22790 50074
rect 22790 50022 22802 50074
rect 22802 50022 22832 50074
rect 22856 50022 22866 50074
rect 22866 50022 22912 50074
rect 22616 50020 22672 50022
rect 22696 50020 22752 50022
rect 22776 50020 22832 50022
rect 22856 50020 22912 50022
rect 27616 50074 27672 50076
rect 27696 50074 27752 50076
rect 27776 50074 27832 50076
rect 27856 50074 27912 50076
rect 27616 50022 27662 50074
rect 27662 50022 27672 50074
rect 27696 50022 27726 50074
rect 27726 50022 27738 50074
rect 27738 50022 27752 50074
rect 27776 50022 27790 50074
rect 27790 50022 27802 50074
rect 27802 50022 27832 50074
rect 27856 50022 27866 50074
rect 27866 50022 27912 50074
rect 27616 50020 27672 50022
rect 27696 50020 27752 50022
rect 27776 50020 27832 50022
rect 27856 50020 27912 50022
rect 32616 50074 32672 50076
rect 32696 50074 32752 50076
rect 32776 50074 32832 50076
rect 32856 50074 32912 50076
rect 32616 50022 32662 50074
rect 32662 50022 32672 50074
rect 32696 50022 32726 50074
rect 32726 50022 32738 50074
rect 32738 50022 32752 50074
rect 32776 50022 32790 50074
rect 32790 50022 32802 50074
rect 32802 50022 32832 50074
rect 32856 50022 32866 50074
rect 32866 50022 32912 50074
rect 32616 50020 32672 50022
rect 32696 50020 32752 50022
rect 32776 50020 32832 50022
rect 32856 50020 32912 50022
rect 37616 50074 37672 50076
rect 37696 50074 37752 50076
rect 37776 50074 37832 50076
rect 37856 50074 37912 50076
rect 37616 50022 37662 50074
rect 37662 50022 37672 50074
rect 37696 50022 37726 50074
rect 37726 50022 37738 50074
rect 37738 50022 37752 50074
rect 37776 50022 37790 50074
rect 37790 50022 37802 50074
rect 37802 50022 37832 50074
rect 37856 50022 37866 50074
rect 37866 50022 37912 50074
rect 37616 50020 37672 50022
rect 37696 50020 37752 50022
rect 37776 50020 37832 50022
rect 37856 50020 37912 50022
rect 42616 50074 42672 50076
rect 42696 50074 42752 50076
rect 42776 50074 42832 50076
rect 42856 50074 42912 50076
rect 42616 50022 42662 50074
rect 42662 50022 42672 50074
rect 42696 50022 42726 50074
rect 42726 50022 42738 50074
rect 42738 50022 42752 50074
rect 42776 50022 42790 50074
rect 42790 50022 42802 50074
rect 42802 50022 42832 50074
rect 42856 50022 42866 50074
rect 42866 50022 42912 50074
rect 42616 50020 42672 50022
rect 42696 50020 42752 50022
rect 42776 50020 42832 50022
rect 42856 50020 42912 50022
rect 47616 50074 47672 50076
rect 47696 50074 47752 50076
rect 47776 50074 47832 50076
rect 47856 50074 47912 50076
rect 47616 50022 47662 50074
rect 47662 50022 47672 50074
rect 47696 50022 47726 50074
rect 47726 50022 47738 50074
rect 47738 50022 47752 50074
rect 47776 50022 47790 50074
rect 47790 50022 47802 50074
rect 47802 50022 47832 50074
rect 47856 50022 47866 50074
rect 47866 50022 47912 50074
rect 47616 50020 47672 50022
rect 47696 50020 47752 50022
rect 47776 50020 47832 50022
rect 47856 50020 47912 50022
rect 52616 50074 52672 50076
rect 52696 50074 52752 50076
rect 52776 50074 52832 50076
rect 52856 50074 52912 50076
rect 52616 50022 52662 50074
rect 52662 50022 52672 50074
rect 52696 50022 52726 50074
rect 52726 50022 52738 50074
rect 52738 50022 52752 50074
rect 52776 50022 52790 50074
rect 52790 50022 52802 50074
rect 52802 50022 52832 50074
rect 52856 50022 52866 50074
rect 52866 50022 52912 50074
rect 52616 50020 52672 50022
rect 52696 50020 52752 50022
rect 52776 50020 52832 50022
rect 52856 50020 52912 50022
rect 57616 50074 57672 50076
rect 57696 50074 57752 50076
rect 57776 50074 57832 50076
rect 57856 50074 57912 50076
rect 57616 50022 57662 50074
rect 57662 50022 57672 50074
rect 57696 50022 57726 50074
rect 57726 50022 57738 50074
rect 57738 50022 57752 50074
rect 57776 50022 57790 50074
rect 57790 50022 57802 50074
rect 57802 50022 57832 50074
rect 57856 50022 57866 50074
rect 57866 50022 57912 50074
rect 57616 50020 57672 50022
rect 57696 50020 57752 50022
rect 57776 50020 57832 50022
rect 57856 50020 57912 50022
rect 58530 49816 58586 49872
rect 1956 49530 2012 49532
rect 2036 49530 2092 49532
rect 2116 49530 2172 49532
rect 2196 49530 2252 49532
rect 1956 49478 2002 49530
rect 2002 49478 2012 49530
rect 2036 49478 2066 49530
rect 2066 49478 2078 49530
rect 2078 49478 2092 49530
rect 2116 49478 2130 49530
rect 2130 49478 2142 49530
rect 2142 49478 2172 49530
rect 2196 49478 2206 49530
rect 2206 49478 2252 49530
rect 1956 49476 2012 49478
rect 2036 49476 2092 49478
rect 2116 49476 2172 49478
rect 2196 49476 2252 49478
rect 6956 49530 7012 49532
rect 7036 49530 7092 49532
rect 7116 49530 7172 49532
rect 7196 49530 7252 49532
rect 6956 49478 7002 49530
rect 7002 49478 7012 49530
rect 7036 49478 7066 49530
rect 7066 49478 7078 49530
rect 7078 49478 7092 49530
rect 7116 49478 7130 49530
rect 7130 49478 7142 49530
rect 7142 49478 7172 49530
rect 7196 49478 7206 49530
rect 7206 49478 7252 49530
rect 6956 49476 7012 49478
rect 7036 49476 7092 49478
rect 7116 49476 7172 49478
rect 7196 49476 7252 49478
rect 11956 49530 12012 49532
rect 12036 49530 12092 49532
rect 12116 49530 12172 49532
rect 12196 49530 12252 49532
rect 11956 49478 12002 49530
rect 12002 49478 12012 49530
rect 12036 49478 12066 49530
rect 12066 49478 12078 49530
rect 12078 49478 12092 49530
rect 12116 49478 12130 49530
rect 12130 49478 12142 49530
rect 12142 49478 12172 49530
rect 12196 49478 12206 49530
rect 12206 49478 12252 49530
rect 11956 49476 12012 49478
rect 12036 49476 12092 49478
rect 12116 49476 12172 49478
rect 12196 49476 12252 49478
rect 16956 49530 17012 49532
rect 17036 49530 17092 49532
rect 17116 49530 17172 49532
rect 17196 49530 17252 49532
rect 16956 49478 17002 49530
rect 17002 49478 17012 49530
rect 17036 49478 17066 49530
rect 17066 49478 17078 49530
rect 17078 49478 17092 49530
rect 17116 49478 17130 49530
rect 17130 49478 17142 49530
rect 17142 49478 17172 49530
rect 17196 49478 17206 49530
rect 17206 49478 17252 49530
rect 16956 49476 17012 49478
rect 17036 49476 17092 49478
rect 17116 49476 17172 49478
rect 17196 49476 17252 49478
rect 21956 49530 22012 49532
rect 22036 49530 22092 49532
rect 22116 49530 22172 49532
rect 22196 49530 22252 49532
rect 21956 49478 22002 49530
rect 22002 49478 22012 49530
rect 22036 49478 22066 49530
rect 22066 49478 22078 49530
rect 22078 49478 22092 49530
rect 22116 49478 22130 49530
rect 22130 49478 22142 49530
rect 22142 49478 22172 49530
rect 22196 49478 22206 49530
rect 22206 49478 22252 49530
rect 21956 49476 22012 49478
rect 22036 49476 22092 49478
rect 22116 49476 22172 49478
rect 22196 49476 22252 49478
rect 26956 49530 27012 49532
rect 27036 49530 27092 49532
rect 27116 49530 27172 49532
rect 27196 49530 27252 49532
rect 26956 49478 27002 49530
rect 27002 49478 27012 49530
rect 27036 49478 27066 49530
rect 27066 49478 27078 49530
rect 27078 49478 27092 49530
rect 27116 49478 27130 49530
rect 27130 49478 27142 49530
rect 27142 49478 27172 49530
rect 27196 49478 27206 49530
rect 27206 49478 27252 49530
rect 26956 49476 27012 49478
rect 27036 49476 27092 49478
rect 27116 49476 27172 49478
rect 27196 49476 27252 49478
rect 31956 49530 32012 49532
rect 32036 49530 32092 49532
rect 32116 49530 32172 49532
rect 32196 49530 32252 49532
rect 31956 49478 32002 49530
rect 32002 49478 32012 49530
rect 32036 49478 32066 49530
rect 32066 49478 32078 49530
rect 32078 49478 32092 49530
rect 32116 49478 32130 49530
rect 32130 49478 32142 49530
rect 32142 49478 32172 49530
rect 32196 49478 32206 49530
rect 32206 49478 32252 49530
rect 31956 49476 32012 49478
rect 32036 49476 32092 49478
rect 32116 49476 32172 49478
rect 32196 49476 32252 49478
rect 36956 49530 37012 49532
rect 37036 49530 37092 49532
rect 37116 49530 37172 49532
rect 37196 49530 37252 49532
rect 36956 49478 37002 49530
rect 37002 49478 37012 49530
rect 37036 49478 37066 49530
rect 37066 49478 37078 49530
rect 37078 49478 37092 49530
rect 37116 49478 37130 49530
rect 37130 49478 37142 49530
rect 37142 49478 37172 49530
rect 37196 49478 37206 49530
rect 37206 49478 37252 49530
rect 36956 49476 37012 49478
rect 37036 49476 37092 49478
rect 37116 49476 37172 49478
rect 37196 49476 37252 49478
rect 41956 49530 42012 49532
rect 42036 49530 42092 49532
rect 42116 49530 42172 49532
rect 42196 49530 42252 49532
rect 41956 49478 42002 49530
rect 42002 49478 42012 49530
rect 42036 49478 42066 49530
rect 42066 49478 42078 49530
rect 42078 49478 42092 49530
rect 42116 49478 42130 49530
rect 42130 49478 42142 49530
rect 42142 49478 42172 49530
rect 42196 49478 42206 49530
rect 42206 49478 42252 49530
rect 41956 49476 42012 49478
rect 42036 49476 42092 49478
rect 42116 49476 42172 49478
rect 42196 49476 42252 49478
rect 46956 49530 47012 49532
rect 47036 49530 47092 49532
rect 47116 49530 47172 49532
rect 47196 49530 47252 49532
rect 46956 49478 47002 49530
rect 47002 49478 47012 49530
rect 47036 49478 47066 49530
rect 47066 49478 47078 49530
rect 47078 49478 47092 49530
rect 47116 49478 47130 49530
rect 47130 49478 47142 49530
rect 47142 49478 47172 49530
rect 47196 49478 47206 49530
rect 47206 49478 47252 49530
rect 46956 49476 47012 49478
rect 47036 49476 47092 49478
rect 47116 49476 47172 49478
rect 47196 49476 47252 49478
rect 51956 49530 52012 49532
rect 52036 49530 52092 49532
rect 52116 49530 52172 49532
rect 52196 49530 52252 49532
rect 51956 49478 52002 49530
rect 52002 49478 52012 49530
rect 52036 49478 52066 49530
rect 52066 49478 52078 49530
rect 52078 49478 52092 49530
rect 52116 49478 52130 49530
rect 52130 49478 52142 49530
rect 52142 49478 52172 49530
rect 52196 49478 52206 49530
rect 52206 49478 52252 49530
rect 51956 49476 52012 49478
rect 52036 49476 52092 49478
rect 52116 49476 52172 49478
rect 52196 49476 52252 49478
rect 56956 49530 57012 49532
rect 57036 49530 57092 49532
rect 57116 49530 57172 49532
rect 57196 49530 57252 49532
rect 56956 49478 57002 49530
rect 57002 49478 57012 49530
rect 57036 49478 57066 49530
rect 57066 49478 57078 49530
rect 57078 49478 57092 49530
rect 57116 49478 57130 49530
rect 57130 49478 57142 49530
rect 57142 49478 57172 49530
rect 57196 49478 57206 49530
rect 57206 49478 57252 49530
rect 56956 49476 57012 49478
rect 57036 49476 57092 49478
rect 57116 49476 57172 49478
rect 57196 49476 57252 49478
rect 58530 49000 58586 49056
rect 2616 48986 2672 48988
rect 2696 48986 2752 48988
rect 2776 48986 2832 48988
rect 2856 48986 2912 48988
rect 2616 48934 2662 48986
rect 2662 48934 2672 48986
rect 2696 48934 2726 48986
rect 2726 48934 2738 48986
rect 2738 48934 2752 48986
rect 2776 48934 2790 48986
rect 2790 48934 2802 48986
rect 2802 48934 2832 48986
rect 2856 48934 2866 48986
rect 2866 48934 2912 48986
rect 2616 48932 2672 48934
rect 2696 48932 2752 48934
rect 2776 48932 2832 48934
rect 2856 48932 2912 48934
rect 7616 48986 7672 48988
rect 7696 48986 7752 48988
rect 7776 48986 7832 48988
rect 7856 48986 7912 48988
rect 7616 48934 7662 48986
rect 7662 48934 7672 48986
rect 7696 48934 7726 48986
rect 7726 48934 7738 48986
rect 7738 48934 7752 48986
rect 7776 48934 7790 48986
rect 7790 48934 7802 48986
rect 7802 48934 7832 48986
rect 7856 48934 7866 48986
rect 7866 48934 7912 48986
rect 7616 48932 7672 48934
rect 7696 48932 7752 48934
rect 7776 48932 7832 48934
rect 7856 48932 7912 48934
rect 12616 48986 12672 48988
rect 12696 48986 12752 48988
rect 12776 48986 12832 48988
rect 12856 48986 12912 48988
rect 12616 48934 12662 48986
rect 12662 48934 12672 48986
rect 12696 48934 12726 48986
rect 12726 48934 12738 48986
rect 12738 48934 12752 48986
rect 12776 48934 12790 48986
rect 12790 48934 12802 48986
rect 12802 48934 12832 48986
rect 12856 48934 12866 48986
rect 12866 48934 12912 48986
rect 12616 48932 12672 48934
rect 12696 48932 12752 48934
rect 12776 48932 12832 48934
rect 12856 48932 12912 48934
rect 17616 48986 17672 48988
rect 17696 48986 17752 48988
rect 17776 48986 17832 48988
rect 17856 48986 17912 48988
rect 17616 48934 17662 48986
rect 17662 48934 17672 48986
rect 17696 48934 17726 48986
rect 17726 48934 17738 48986
rect 17738 48934 17752 48986
rect 17776 48934 17790 48986
rect 17790 48934 17802 48986
rect 17802 48934 17832 48986
rect 17856 48934 17866 48986
rect 17866 48934 17912 48986
rect 17616 48932 17672 48934
rect 17696 48932 17752 48934
rect 17776 48932 17832 48934
rect 17856 48932 17912 48934
rect 22616 48986 22672 48988
rect 22696 48986 22752 48988
rect 22776 48986 22832 48988
rect 22856 48986 22912 48988
rect 22616 48934 22662 48986
rect 22662 48934 22672 48986
rect 22696 48934 22726 48986
rect 22726 48934 22738 48986
rect 22738 48934 22752 48986
rect 22776 48934 22790 48986
rect 22790 48934 22802 48986
rect 22802 48934 22832 48986
rect 22856 48934 22866 48986
rect 22866 48934 22912 48986
rect 22616 48932 22672 48934
rect 22696 48932 22752 48934
rect 22776 48932 22832 48934
rect 22856 48932 22912 48934
rect 27616 48986 27672 48988
rect 27696 48986 27752 48988
rect 27776 48986 27832 48988
rect 27856 48986 27912 48988
rect 27616 48934 27662 48986
rect 27662 48934 27672 48986
rect 27696 48934 27726 48986
rect 27726 48934 27738 48986
rect 27738 48934 27752 48986
rect 27776 48934 27790 48986
rect 27790 48934 27802 48986
rect 27802 48934 27832 48986
rect 27856 48934 27866 48986
rect 27866 48934 27912 48986
rect 27616 48932 27672 48934
rect 27696 48932 27752 48934
rect 27776 48932 27832 48934
rect 27856 48932 27912 48934
rect 32616 48986 32672 48988
rect 32696 48986 32752 48988
rect 32776 48986 32832 48988
rect 32856 48986 32912 48988
rect 32616 48934 32662 48986
rect 32662 48934 32672 48986
rect 32696 48934 32726 48986
rect 32726 48934 32738 48986
rect 32738 48934 32752 48986
rect 32776 48934 32790 48986
rect 32790 48934 32802 48986
rect 32802 48934 32832 48986
rect 32856 48934 32866 48986
rect 32866 48934 32912 48986
rect 32616 48932 32672 48934
rect 32696 48932 32752 48934
rect 32776 48932 32832 48934
rect 32856 48932 32912 48934
rect 37616 48986 37672 48988
rect 37696 48986 37752 48988
rect 37776 48986 37832 48988
rect 37856 48986 37912 48988
rect 37616 48934 37662 48986
rect 37662 48934 37672 48986
rect 37696 48934 37726 48986
rect 37726 48934 37738 48986
rect 37738 48934 37752 48986
rect 37776 48934 37790 48986
rect 37790 48934 37802 48986
rect 37802 48934 37832 48986
rect 37856 48934 37866 48986
rect 37866 48934 37912 48986
rect 37616 48932 37672 48934
rect 37696 48932 37752 48934
rect 37776 48932 37832 48934
rect 37856 48932 37912 48934
rect 42616 48986 42672 48988
rect 42696 48986 42752 48988
rect 42776 48986 42832 48988
rect 42856 48986 42912 48988
rect 42616 48934 42662 48986
rect 42662 48934 42672 48986
rect 42696 48934 42726 48986
rect 42726 48934 42738 48986
rect 42738 48934 42752 48986
rect 42776 48934 42790 48986
rect 42790 48934 42802 48986
rect 42802 48934 42832 48986
rect 42856 48934 42866 48986
rect 42866 48934 42912 48986
rect 42616 48932 42672 48934
rect 42696 48932 42752 48934
rect 42776 48932 42832 48934
rect 42856 48932 42912 48934
rect 47616 48986 47672 48988
rect 47696 48986 47752 48988
rect 47776 48986 47832 48988
rect 47856 48986 47912 48988
rect 47616 48934 47662 48986
rect 47662 48934 47672 48986
rect 47696 48934 47726 48986
rect 47726 48934 47738 48986
rect 47738 48934 47752 48986
rect 47776 48934 47790 48986
rect 47790 48934 47802 48986
rect 47802 48934 47832 48986
rect 47856 48934 47866 48986
rect 47866 48934 47912 48986
rect 47616 48932 47672 48934
rect 47696 48932 47752 48934
rect 47776 48932 47832 48934
rect 47856 48932 47912 48934
rect 52616 48986 52672 48988
rect 52696 48986 52752 48988
rect 52776 48986 52832 48988
rect 52856 48986 52912 48988
rect 52616 48934 52662 48986
rect 52662 48934 52672 48986
rect 52696 48934 52726 48986
rect 52726 48934 52738 48986
rect 52738 48934 52752 48986
rect 52776 48934 52790 48986
rect 52790 48934 52802 48986
rect 52802 48934 52832 48986
rect 52856 48934 52866 48986
rect 52866 48934 52912 48986
rect 52616 48932 52672 48934
rect 52696 48932 52752 48934
rect 52776 48932 52832 48934
rect 52856 48932 52912 48934
rect 57616 48986 57672 48988
rect 57696 48986 57752 48988
rect 57776 48986 57832 48988
rect 57856 48986 57912 48988
rect 57616 48934 57662 48986
rect 57662 48934 57672 48986
rect 57696 48934 57726 48986
rect 57726 48934 57738 48986
rect 57738 48934 57752 48986
rect 57776 48934 57790 48986
rect 57790 48934 57802 48986
rect 57802 48934 57832 48986
rect 57856 48934 57866 48986
rect 57866 48934 57912 48986
rect 57616 48932 57672 48934
rect 57696 48932 57752 48934
rect 57776 48932 57832 48934
rect 57856 48932 57912 48934
rect 1956 48442 2012 48444
rect 2036 48442 2092 48444
rect 2116 48442 2172 48444
rect 2196 48442 2252 48444
rect 1956 48390 2002 48442
rect 2002 48390 2012 48442
rect 2036 48390 2066 48442
rect 2066 48390 2078 48442
rect 2078 48390 2092 48442
rect 2116 48390 2130 48442
rect 2130 48390 2142 48442
rect 2142 48390 2172 48442
rect 2196 48390 2206 48442
rect 2206 48390 2252 48442
rect 1956 48388 2012 48390
rect 2036 48388 2092 48390
rect 2116 48388 2172 48390
rect 2196 48388 2252 48390
rect 6956 48442 7012 48444
rect 7036 48442 7092 48444
rect 7116 48442 7172 48444
rect 7196 48442 7252 48444
rect 6956 48390 7002 48442
rect 7002 48390 7012 48442
rect 7036 48390 7066 48442
rect 7066 48390 7078 48442
rect 7078 48390 7092 48442
rect 7116 48390 7130 48442
rect 7130 48390 7142 48442
rect 7142 48390 7172 48442
rect 7196 48390 7206 48442
rect 7206 48390 7252 48442
rect 6956 48388 7012 48390
rect 7036 48388 7092 48390
rect 7116 48388 7172 48390
rect 7196 48388 7252 48390
rect 11956 48442 12012 48444
rect 12036 48442 12092 48444
rect 12116 48442 12172 48444
rect 12196 48442 12252 48444
rect 11956 48390 12002 48442
rect 12002 48390 12012 48442
rect 12036 48390 12066 48442
rect 12066 48390 12078 48442
rect 12078 48390 12092 48442
rect 12116 48390 12130 48442
rect 12130 48390 12142 48442
rect 12142 48390 12172 48442
rect 12196 48390 12206 48442
rect 12206 48390 12252 48442
rect 11956 48388 12012 48390
rect 12036 48388 12092 48390
rect 12116 48388 12172 48390
rect 12196 48388 12252 48390
rect 16956 48442 17012 48444
rect 17036 48442 17092 48444
rect 17116 48442 17172 48444
rect 17196 48442 17252 48444
rect 16956 48390 17002 48442
rect 17002 48390 17012 48442
rect 17036 48390 17066 48442
rect 17066 48390 17078 48442
rect 17078 48390 17092 48442
rect 17116 48390 17130 48442
rect 17130 48390 17142 48442
rect 17142 48390 17172 48442
rect 17196 48390 17206 48442
rect 17206 48390 17252 48442
rect 16956 48388 17012 48390
rect 17036 48388 17092 48390
rect 17116 48388 17172 48390
rect 17196 48388 17252 48390
rect 21956 48442 22012 48444
rect 22036 48442 22092 48444
rect 22116 48442 22172 48444
rect 22196 48442 22252 48444
rect 21956 48390 22002 48442
rect 22002 48390 22012 48442
rect 22036 48390 22066 48442
rect 22066 48390 22078 48442
rect 22078 48390 22092 48442
rect 22116 48390 22130 48442
rect 22130 48390 22142 48442
rect 22142 48390 22172 48442
rect 22196 48390 22206 48442
rect 22206 48390 22252 48442
rect 21956 48388 22012 48390
rect 22036 48388 22092 48390
rect 22116 48388 22172 48390
rect 22196 48388 22252 48390
rect 26956 48442 27012 48444
rect 27036 48442 27092 48444
rect 27116 48442 27172 48444
rect 27196 48442 27252 48444
rect 26956 48390 27002 48442
rect 27002 48390 27012 48442
rect 27036 48390 27066 48442
rect 27066 48390 27078 48442
rect 27078 48390 27092 48442
rect 27116 48390 27130 48442
rect 27130 48390 27142 48442
rect 27142 48390 27172 48442
rect 27196 48390 27206 48442
rect 27206 48390 27252 48442
rect 26956 48388 27012 48390
rect 27036 48388 27092 48390
rect 27116 48388 27172 48390
rect 27196 48388 27252 48390
rect 31956 48442 32012 48444
rect 32036 48442 32092 48444
rect 32116 48442 32172 48444
rect 32196 48442 32252 48444
rect 31956 48390 32002 48442
rect 32002 48390 32012 48442
rect 32036 48390 32066 48442
rect 32066 48390 32078 48442
rect 32078 48390 32092 48442
rect 32116 48390 32130 48442
rect 32130 48390 32142 48442
rect 32142 48390 32172 48442
rect 32196 48390 32206 48442
rect 32206 48390 32252 48442
rect 31956 48388 32012 48390
rect 32036 48388 32092 48390
rect 32116 48388 32172 48390
rect 32196 48388 32252 48390
rect 36956 48442 37012 48444
rect 37036 48442 37092 48444
rect 37116 48442 37172 48444
rect 37196 48442 37252 48444
rect 36956 48390 37002 48442
rect 37002 48390 37012 48442
rect 37036 48390 37066 48442
rect 37066 48390 37078 48442
rect 37078 48390 37092 48442
rect 37116 48390 37130 48442
rect 37130 48390 37142 48442
rect 37142 48390 37172 48442
rect 37196 48390 37206 48442
rect 37206 48390 37252 48442
rect 36956 48388 37012 48390
rect 37036 48388 37092 48390
rect 37116 48388 37172 48390
rect 37196 48388 37252 48390
rect 41956 48442 42012 48444
rect 42036 48442 42092 48444
rect 42116 48442 42172 48444
rect 42196 48442 42252 48444
rect 41956 48390 42002 48442
rect 42002 48390 42012 48442
rect 42036 48390 42066 48442
rect 42066 48390 42078 48442
rect 42078 48390 42092 48442
rect 42116 48390 42130 48442
rect 42130 48390 42142 48442
rect 42142 48390 42172 48442
rect 42196 48390 42206 48442
rect 42206 48390 42252 48442
rect 41956 48388 42012 48390
rect 42036 48388 42092 48390
rect 42116 48388 42172 48390
rect 42196 48388 42252 48390
rect 46956 48442 47012 48444
rect 47036 48442 47092 48444
rect 47116 48442 47172 48444
rect 47196 48442 47252 48444
rect 46956 48390 47002 48442
rect 47002 48390 47012 48442
rect 47036 48390 47066 48442
rect 47066 48390 47078 48442
rect 47078 48390 47092 48442
rect 47116 48390 47130 48442
rect 47130 48390 47142 48442
rect 47142 48390 47172 48442
rect 47196 48390 47206 48442
rect 47206 48390 47252 48442
rect 46956 48388 47012 48390
rect 47036 48388 47092 48390
rect 47116 48388 47172 48390
rect 47196 48388 47252 48390
rect 51956 48442 52012 48444
rect 52036 48442 52092 48444
rect 52116 48442 52172 48444
rect 52196 48442 52252 48444
rect 51956 48390 52002 48442
rect 52002 48390 52012 48442
rect 52036 48390 52066 48442
rect 52066 48390 52078 48442
rect 52078 48390 52092 48442
rect 52116 48390 52130 48442
rect 52130 48390 52142 48442
rect 52142 48390 52172 48442
rect 52196 48390 52206 48442
rect 52206 48390 52252 48442
rect 51956 48388 52012 48390
rect 52036 48388 52092 48390
rect 52116 48388 52172 48390
rect 52196 48388 52252 48390
rect 56956 48442 57012 48444
rect 57036 48442 57092 48444
rect 57116 48442 57172 48444
rect 57196 48442 57252 48444
rect 56956 48390 57002 48442
rect 57002 48390 57012 48442
rect 57036 48390 57066 48442
rect 57066 48390 57078 48442
rect 57078 48390 57092 48442
rect 57116 48390 57130 48442
rect 57130 48390 57142 48442
rect 57142 48390 57172 48442
rect 57196 48390 57206 48442
rect 57206 48390 57252 48442
rect 56956 48388 57012 48390
rect 57036 48388 57092 48390
rect 57116 48388 57172 48390
rect 57196 48388 57252 48390
rect 58530 48184 58586 48240
rect 2616 47898 2672 47900
rect 2696 47898 2752 47900
rect 2776 47898 2832 47900
rect 2856 47898 2912 47900
rect 2616 47846 2662 47898
rect 2662 47846 2672 47898
rect 2696 47846 2726 47898
rect 2726 47846 2738 47898
rect 2738 47846 2752 47898
rect 2776 47846 2790 47898
rect 2790 47846 2802 47898
rect 2802 47846 2832 47898
rect 2856 47846 2866 47898
rect 2866 47846 2912 47898
rect 2616 47844 2672 47846
rect 2696 47844 2752 47846
rect 2776 47844 2832 47846
rect 2856 47844 2912 47846
rect 7616 47898 7672 47900
rect 7696 47898 7752 47900
rect 7776 47898 7832 47900
rect 7856 47898 7912 47900
rect 7616 47846 7662 47898
rect 7662 47846 7672 47898
rect 7696 47846 7726 47898
rect 7726 47846 7738 47898
rect 7738 47846 7752 47898
rect 7776 47846 7790 47898
rect 7790 47846 7802 47898
rect 7802 47846 7832 47898
rect 7856 47846 7866 47898
rect 7866 47846 7912 47898
rect 7616 47844 7672 47846
rect 7696 47844 7752 47846
rect 7776 47844 7832 47846
rect 7856 47844 7912 47846
rect 12616 47898 12672 47900
rect 12696 47898 12752 47900
rect 12776 47898 12832 47900
rect 12856 47898 12912 47900
rect 12616 47846 12662 47898
rect 12662 47846 12672 47898
rect 12696 47846 12726 47898
rect 12726 47846 12738 47898
rect 12738 47846 12752 47898
rect 12776 47846 12790 47898
rect 12790 47846 12802 47898
rect 12802 47846 12832 47898
rect 12856 47846 12866 47898
rect 12866 47846 12912 47898
rect 12616 47844 12672 47846
rect 12696 47844 12752 47846
rect 12776 47844 12832 47846
rect 12856 47844 12912 47846
rect 17616 47898 17672 47900
rect 17696 47898 17752 47900
rect 17776 47898 17832 47900
rect 17856 47898 17912 47900
rect 17616 47846 17662 47898
rect 17662 47846 17672 47898
rect 17696 47846 17726 47898
rect 17726 47846 17738 47898
rect 17738 47846 17752 47898
rect 17776 47846 17790 47898
rect 17790 47846 17802 47898
rect 17802 47846 17832 47898
rect 17856 47846 17866 47898
rect 17866 47846 17912 47898
rect 17616 47844 17672 47846
rect 17696 47844 17752 47846
rect 17776 47844 17832 47846
rect 17856 47844 17912 47846
rect 22616 47898 22672 47900
rect 22696 47898 22752 47900
rect 22776 47898 22832 47900
rect 22856 47898 22912 47900
rect 22616 47846 22662 47898
rect 22662 47846 22672 47898
rect 22696 47846 22726 47898
rect 22726 47846 22738 47898
rect 22738 47846 22752 47898
rect 22776 47846 22790 47898
rect 22790 47846 22802 47898
rect 22802 47846 22832 47898
rect 22856 47846 22866 47898
rect 22866 47846 22912 47898
rect 22616 47844 22672 47846
rect 22696 47844 22752 47846
rect 22776 47844 22832 47846
rect 22856 47844 22912 47846
rect 27616 47898 27672 47900
rect 27696 47898 27752 47900
rect 27776 47898 27832 47900
rect 27856 47898 27912 47900
rect 27616 47846 27662 47898
rect 27662 47846 27672 47898
rect 27696 47846 27726 47898
rect 27726 47846 27738 47898
rect 27738 47846 27752 47898
rect 27776 47846 27790 47898
rect 27790 47846 27802 47898
rect 27802 47846 27832 47898
rect 27856 47846 27866 47898
rect 27866 47846 27912 47898
rect 27616 47844 27672 47846
rect 27696 47844 27752 47846
rect 27776 47844 27832 47846
rect 27856 47844 27912 47846
rect 32616 47898 32672 47900
rect 32696 47898 32752 47900
rect 32776 47898 32832 47900
rect 32856 47898 32912 47900
rect 32616 47846 32662 47898
rect 32662 47846 32672 47898
rect 32696 47846 32726 47898
rect 32726 47846 32738 47898
rect 32738 47846 32752 47898
rect 32776 47846 32790 47898
rect 32790 47846 32802 47898
rect 32802 47846 32832 47898
rect 32856 47846 32866 47898
rect 32866 47846 32912 47898
rect 32616 47844 32672 47846
rect 32696 47844 32752 47846
rect 32776 47844 32832 47846
rect 32856 47844 32912 47846
rect 37616 47898 37672 47900
rect 37696 47898 37752 47900
rect 37776 47898 37832 47900
rect 37856 47898 37912 47900
rect 37616 47846 37662 47898
rect 37662 47846 37672 47898
rect 37696 47846 37726 47898
rect 37726 47846 37738 47898
rect 37738 47846 37752 47898
rect 37776 47846 37790 47898
rect 37790 47846 37802 47898
rect 37802 47846 37832 47898
rect 37856 47846 37866 47898
rect 37866 47846 37912 47898
rect 37616 47844 37672 47846
rect 37696 47844 37752 47846
rect 37776 47844 37832 47846
rect 37856 47844 37912 47846
rect 42616 47898 42672 47900
rect 42696 47898 42752 47900
rect 42776 47898 42832 47900
rect 42856 47898 42912 47900
rect 42616 47846 42662 47898
rect 42662 47846 42672 47898
rect 42696 47846 42726 47898
rect 42726 47846 42738 47898
rect 42738 47846 42752 47898
rect 42776 47846 42790 47898
rect 42790 47846 42802 47898
rect 42802 47846 42832 47898
rect 42856 47846 42866 47898
rect 42866 47846 42912 47898
rect 42616 47844 42672 47846
rect 42696 47844 42752 47846
rect 42776 47844 42832 47846
rect 42856 47844 42912 47846
rect 47616 47898 47672 47900
rect 47696 47898 47752 47900
rect 47776 47898 47832 47900
rect 47856 47898 47912 47900
rect 47616 47846 47662 47898
rect 47662 47846 47672 47898
rect 47696 47846 47726 47898
rect 47726 47846 47738 47898
rect 47738 47846 47752 47898
rect 47776 47846 47790 47898
rect 47790 47846 47802 47898
rect 47802 47846 47832 47898
rect 47856 47846 47866 47898
rect 47866 47846 47912 47898
rect 47616 47844 47672 47846
rect 47696 47844 47752 47846
rect 47776 47844 47832 47846
rect 47856 47844 47912 47846
rect 52616 47898 52672 47900
rect 52696 47898 52752 47900
rect 52776 47898 52832 47900
rect 52856 47898 52912 47900
rect 52616 47846 52662 47898
rect 52662 47846 52672 47898
rect 52696 47846 52726 47898
rect 52726 47846 52738 47898
rect 52738 47846 52752 47898
rect 52776 47846 52790 47898
rect 52790 47846 52802 47898
rect 52802 47846 52832 47898
rect 52856 47846 52866 47898
rect 52866 47846 52912 47898
rect 52616 47844 52672 47846
rect 52696 47844 52752 47846
rect 52776 47844 52832 47846
rect 52856 47844 52912 47846
rect 57616 47898 57672 47900
rect 57696 47898 57752 47900
rect 57776 47898 57832 47900
rect 57856 47898 57912 47900
rect 57616 47846 57662 47898
rect 57662 47846 57672 47898
rect 57696 47846 57726 47898
rect 57726 47846 57738 47898
rect 57738 47846 57752 47898
rect 57776 47846 57790 47898
rect 57790 47846 57802 47898
rect 57802 47846 57832 47898
rect 57856 47846 57866 47898
rect 57866 47846 57912 47898
rect 57616 47844 57672 47846
rect 57696 47844 57752 47846
rect 57776 47844 57832 47846
rect 57856 47844 57912 47846
rect 58530 47404 58532 47424
rect 58532 47404 58584 47424
rect 58584 47404 58586 47424
rect 58530 47368 58586 47404
rect 1956 47354 2012 47356
rect 2036 47354 2092 47356
rect 2116 47354 2172 47356
rect 2196 47354 2252 47356
rect 1956 47302 2002 47354
rect 2002 47302 2012 47354
rect 2036 47302 2066 47354
rect 2066 47302 2078 47354
rect 2078 47302 2092 47354
rect 2116 47302 2130 47354
rect 2130 47302 2142 47354
rect 2142 47302 2172 47354
rect 2196 47302 2206 47354
rect 2206 47302 2252 47354
rect 1956 47300 2012 47302
rect 2036 47300 2092 47302
rect 2116 47300 2172 47302
rect 2196 47300 2252 47302
rect 6956 47354 7012 47356
rect 7036 47354 7092 47356
rect 7116 47354 7172 47356
rect 7196 47354 7252 47356
rect 6956 47302 7002 47354
rect 7002 47302 7012 47354
rect 7036 47302 7066 47354
rect 7066 47302 7078 47354
rect 7078 47302 7092 47354
rect 7116 47302 7130 47354
rect 7130 47302 7142 47354
rect 7142 47302 7172 47354
rect 7196 47302 7206 47354
rect 7206 47302 7252 47354
rect 6956 47300 7012 47302
rect 7036 47300 7092 47302
rect 7116 47300 7172 47302
rect 7196 47300 7252 47302
rect 11956 47354 12012 47356
rect 12036 47354 12092 47356
rect 12116 47354 12172 47356
rect 12196 47354 12252 47356
rect 11956 47302 12002 47354
rect 12002 47302 12012 47354
rect 12036 47302 12066 47354
rect 12066 47302 12078 47354
rect 12078 47302 12092 47354
rect 12116 47302 12130 47354
rect 12130 47302 12142 47354
rect 12142 47302 12172 47354
rect 12196 47302 12206 47354
rect 12206 47302 12252 47354
rect 11956 47300 12012 47302
rect 12036 47300 12092 47302
rect 12116 47300 12172 47302
rect 12196 47300 12252 47302
rect 16956 47354 17012 47356
rect 17036 47354 17092 47356
rect 17116 47354 17172 47356
rect 17196 47354 17252 47356
rect 16956 47302 17002 47354
rect 17002 47302 17012 47354
rect 17036 47302 17066 47354
rect 17066 47302 17078 47354
rect 17078 47302 17092 47354
rect 17116 47302 17130 47354
rect 17130 47302 17142 47354
rect 17142 47302 17172 47354
rect 17196 47302 17206 47354
rect 17206 47302 17252 47354
rect 16956 47300 17012 47302
rect 17036 47300 17092 47302
rect 17116 47300 17172 47302
rect 17196 47300 17252 47302
rect 21956 47354 22012 47356
rect 22036 47354 22092 47356
rect 22116 47354 22172 47356
rect 22196 47354 22252 47356
rect 21956 47302 22002 47354
rect 22002 47302 22012 47354
rect 22036 47302 22066 47354
rect 22066 47302 22078 47354
rect 22078 47302 22092 47354
rect 22116 47302 22130 47354
rect 22130 47302 22142 47354
rect 22142 47302 22172 47354
rect 22196 47302 22206 47354
rect 22206 47302 22252 47354
rect 21956 47300 22012 47302
rect 22036 47300 22092 47302
rect 22116 47300 22172 47302
rect 22196 47300 22252 47302
rect 26956 47354 27012 47356
rect 27036 47354 27092 47356
rect 27116 47354 27172 47356
rect 27196 47354 27252 47356
rect 26956 47302 27002 47354
rect 27002 47302 27012 47354
rect 27036 47302 27066 47354
rect 27066 47302 27078 47354
rect 27078 47302 27092 47354
rect 27116 47302 27130 47354
rect 27130 47302 27142 47354
rect 27142 47302 27172 47354
rect 27196 47302 27206 47354
rect 27206 47302 27252 47354
rect 26956 47300 27012 47302
rect 27036 47300 27092 47302
rect 27116 47300 27172 47302
rect 27196 47300 27252 47302
rect 31956 47354 32012 47356
rect 32036 47354 32092 47356
rect 32116 47354 32172 47356
rect 32196 47354 32252 47356
rect 31956 47302 32002 47354
rect 32002 47302 32012 47354
rect 32036 47302 32066 47354
rect 32066 47302 32078 47354
rect 32078 47302 32092 47354
rect 32116 47302 32130 47354
rect 32130 47302 32142 47354
rect 32142 47302 32172 47354
rect 32196 47302 32206 47354
rect 32206 47302 32252 47354
rect 31956 47300 32012 47302
rect 32036 47300 32092 47302
rect 32116 47300 32172 47302
rect 32196 47300 32252 47302
rect 36956 47354 37012 47356
rect 37036 47354 37092 47356
rect 37116 47354 37172 47356
rect 37196 47354 37252 47356
rect 36956 47302 37002 47354
rect 37002 47302 37012 47354
rect 37036 47302 37066 47354
rect 37066 47302 37078 47354
rect 37078 47302 37092 47354
rect 37116 47302 37130 47354
rect 37130 47302 37142 47354
rect 37142 47302 37172 47354
rect 37196 47302 37206 47354
rect 37206 47302 37252 47354
rect 36956 47300 37012 47302
rect 37036 47300 37092 47302
rect 37116 47300 37172 47302
rect 37196 47300 37252 47302
rect 41956 47354 42012 47356
rect 42036 47354 42092 47356
rect 42116 47354 42172 47356
rect 42196 47354 42252 47356
rect 41956 47302 42002 47354
rect 42002 47302 42012 47354
rect 42036 47302 42066 47354
rect 42066 47302 42078 47354
rect 42078 47302 42092 47354
rect 42116 47302 42130 47354
rect 42130 47302 42142 47354
rect 42142 47302 42172 47354
rect 42196 47302 42206 47354
rect 42206 47302 42252 47354
rect 41956 47300 42012 47302
rect 42036 47300 42092 47302
rect 42116 47300 42172 47302
rect 42196 47300 42252 47302
rect 46956 47354 47012 47356
rect 47036 47354 47092 47356
rect 47116 47354 47172 47356
rect 47196 47354 47252 47356
rect 46956 47302 47002 47354
rect 47002 47302 47012 47354
rect 47036 47302 47066 47354
rect 47066 47302 47078 47354
rect 47078 47302 47092 47354
rect 47116 47302 47130 47354
rect 47130 47302 47142 47354
rect 47142 47302 47172 47354
rect 47196 47302 47206 47354
rect 47206 47302 47252 47354
rect 46956 47300 47012 47302
rect 47036 47300 47092 47302
rect 47116 47300 47172 47302
rect 47196 47300 47252 47302
rect 51956 47354 52012 47356
rect 52036 47354 52092 47356
rect 52116 47354 52172 47356
rect 52196 47354 52252 47356
rect 51956 47302 52002 47354
rect 52002 47302 52012 47354
rect 52036 47302 52066 47354
rect 52066 47302 52078 47354
rect 52078 47302 52092 47354
rect 52116 47302 52130 47354
rect 52130 47302 52142 47354
rect 52142 47302 52172 47354
rect 52196 47302 52206 47354
rect 52206 47302 52252 47354
rect 51956 47300 52012 47302
rect 52036 47300 52092 47302
rect 52116 47300 52172 47302
rect 52196 47300 52252 47302
rect 56956 47354 57012 47356
rect 57036 47354 57092 47356
rect 57116 47354 57172 47356
rect 57196 47354 57252 47356
rect 56956 47302 57002 47354
rect 57002 47302 57012 47354
rect 57036 47302 57066 47354
rect 57066 47302 57078 47354
rect 57078 47302 57092 47354
rect 57116 47302 57130 47354
rect 57130 47302 57142 47354
rect 57142 47302 57172 47354
rect 57196 47302 57206 47354
rect 57206 47302 57252 47354
rect 56956 47300 57012 47302
rect 57036 47300 57092 47302
rect 57116 47300 57172 47302
rect 57196 47300 57252 47302
rect 2616 46810 2672 46812
rect 2696 46810 2752 46812
rect 2776 46810 2832 46812
rect 2856 46810 2912 46812
rect 2616 46758 2662 46810
rect 2662 46758 2672 46810
rect 2696 46758 2726 46810
rect 2726 46758 2738 46810
rect 2738 46758 2752 46810
rect 2776 46758 2790 46810
rect 2790 46758 2802 46810
rect 2802 46758 2832 46810
rect 2856 46758 2866 46810
rect 2866 46758 2912 46810
rect 2616 46756 2672 46758
rect 2696 46756 2752 46758
rect 2776 46756 2832 46758
rect 2856 46756 2912 46758
rect 7616 46810 7672 46812
rect 7696 46810 7752 46812
rect 7776 46810 7832 46812
rect 7856 46810 7912 46812
rect 7616 46758 7662 46810
rect 7662 46758 7672 46810
rect 7696 46758 7726 46810
rect 7726 46758 7738 46810
rect 7738 46758 7752 46810
rect 7776 46758 7790 46810
rect 7790 46758 7802 46810
rect 7802 46758 7832 46810
rect 7856 46758 7866 46810
rect 7866 46758 7912 46810
rect 7616 46756 7672 46758
rect 7696 46756 7752 46758
rect 7776 46756 7832 46758
rect 7856 46756 7912 46758
rect 12616 46810 12672 46812
rect 12696 46810 12752 46812
rect 12776 46810 12832 46812
rect 12856 46810 12912 46812
rect 12616 46758 12662 46810
rect 12662 46758 12672 46810
rect 12696 46758 12726 46810
rect 12726 46758 12738 46810
rect 12738 46758 12752 46810
rect 12776 46758 12790 46810
rect 12790 46758 12802 46810
rect 12802 46758 12832 46810
rect 12856 46758 12866 46810
rect 12866 46758 12912 46810
rect 12616 46756 12672 46758
rect 12696 46756 12752 46758
rect 12776 46756 12832 46758
rect 12856 46756 12912 46758
rect 17616 46810 17672 46812
rect 17696 46810 17752 46812
rect 17776 46810 17832 46812
rect 17856 46810 17912 46812
rect 17616 46758 17662 46810
rect 17662 46758 17672 46810
rect 17696 46758 17726 46810
rect 17726 46758 17738 46810
rect 17738 46758 17752 46810
rect 17776 46758 17790 46810
rect 17790 46758 17802 46810
rect 17802 46758 17832 46810
rect 17856 46758 17866 46810
rect 17866 46758 17912 46810
rect 17616 46756 17672 46758
rect 17696 46756 17752 46758
rect 17776 46756 17832 46758
rect 17856 46756 17912 46758
rect 22616 46810 22672 46812
rect 22696 46810 22752 46812
rect 22776 46810 22832 46812
rect 22856 46810 22912 46812
rect 22616 46758 22662 46810
rect 22662 46758 22672 46810
rect 22696 46758 22726 46810
rect 22726 46758 22738 46810
rect 22738 46758 22752 46810
rect 22776 46758 22790 46810
rect 22790 46758 22802 46810
rect 22802 46758 22832 46810
rect 22856 46758 22866 46810
rect 22866 46758 22912 46810
rect 22616 46756 22672 46758
rect 22696 46756 22752 46758
rect 22776 46756 22832 46758
rect 22856 46756 22912 46758
rect 27616 46810 27672 46812
rect 27696 46810 27752 46812
rect 27776 46810 27832 46812
rect 27856 46810 27912 46812
rect 27616 46758 27662 46810
rect 27662 46758 27672 46810
rect 27696 46758 27726 46810
rect 27726 46758 27738 46810
rect 27738 46758 27752 46810
rect 27776 46758 27790 46810
rect 27790 46758 27802 46810
rect 27802 46758 27832 46810
rect 27856 46758 27866 46810
rect 27866 46758 27912 46810
rect 27616 46756 27672 46758
rect 27696 46756 27752 46758
rect 27776 46756 27832 46758
rect 27856 46756 27912 46758
rect 32616 46810 32672 46812
rect 32696 46810 32752 46812
rect 32776 46810 32832 46812
rect 32856 46810 32912 46812
rect 32616 46758 32662 46810
rect 32662 46758 32672 46810
rect 32696 46758 32726 46810
rect 32726 46758 32738 46810
rect 32738 46758 32752 46810
rect 32776 46758 32790 46810
rect 32790 46758 32802 46810
rect 32802 46758 32832 46810
rect 32856 46758 32866 46810
rect 32866 46758 32912 46810
rect 32616 46756 32672 46758
rect 32696 46756 32752 46758
rect 32776 46756 32832 46758
rect 32856 46756 32912 46758
rect 37616 46810 37672 46812
rect 37696 46810 37752 46812
rect 37776 46810 37832 46812
rect 37856 46810 37912 46812
rect 37616 46758 37662 46810
rect 37662 46758 37672 46810
rect 37696 46758 37726 46810
rect 37726 46758 37738 46810
rect 37738 46758 37752 46810
rect 37776 46758 37790 46810
rect 37790 46758 37802 46810
rect 37802 46758 37832 46810
rect 37856 46758 37866 46810
rect 37866 46758 37912 46810
rect 37616 46756 37672 46758
rect 37696 46756 37752 46758
rect 37776 46756 37832 46758
rect 37856 46756 37912 46758
rect 42616 46810 42672 46812
rect 42696 46810 42752 46812
rect 42776 46810 42832 46812
rect 42856 46810 42912 46812
rect 42616 46758 42662 46810
rect 42662 46758 42672 46810
rect 42696 46758 42726 46810
rect 42726 46758 42738 46810
rect 42738 46758 42752 46810
rect 42776 46758 42790 46810
rect 42790 46758 42802 46810
rect 42802 46758 42832 46810
rect 42856 46758 42866 46810
rect 42866 46758 42912 46810
rect 42616 46756 42672 46758
rect 42696 46756 42752 46758
rect 42776 46756 42832 46758
rect 42856 46756 42912 46758
rect 47616 46810 47672 46812
rect 47696 46810 47752 46812
rect 47776 46810 47832 46812
rect 47856 46810 47912 46812
rect 47616 46758 47662 46810
rect 47662 46758 47672 46810
rect 47696 46758 47726 46810
rect 47726 46758 47738 46810
rect 47738 46758 47752 46810
rect 47776 46758 47790 46810
rect 47790 46758 47802 46810
rect 47802 46758 47832 46810
rect 47856 46758 47866 46810
rect 47866 46758 47912 46810
rect 47616 46756 47672 46758
rect 47696 46756 47752 46758
rect 47776 46756 47832 46758
rect 47856 46756 47912 46758
rect 52616 46810 52672 46812
rect 52696 46810 52752 46812
rect 52776 46810 52832 46812
rect 52856 46810 52912 46812
rect 52616 46758 52662 46810
rect 52662 46758 52672 46810
rect 52696 46758 52726 46810
rect 52726 46758 52738 46810
rect 52738 46758 52752 46810
rect 52776 46758 52790 46810
rect 52790 46758 52802 46810
rect 52802 46758 52832 46810
rect 52856 46758 52866 46810
rect 52866 46758 52912 46810
rect 52616 46756 52672 46758
rect 52696 46756 52752 46758
rect 52776 46756 52832 46758
rect 52856 46756 52912 46758
rect 57616 46810 57672 46812
rect 57696 46810 57752 46812
rect 57776 46810 57832 46812
rect 57856 46810 57912 46812
rect 57616 46758 57662 46810
rect 57662 46758 57672 46810
rect 57696 46758 57726 46810
rect 57726 46758 57738 46810
rect 57738 46758 57752 46810
rect 57776 46758 57790 46810
rect 57790 46758 57802 46810
rect 57802 46758 57832 46810
rect 57856 46758 57866 46810
rect 57866 46758 57912 46810
rect 57616 46756 57672 46758
rect 57696 46756 57752 46758
rect 57776 46756 57832 46758
rect 57856 46756 57912 46758
rect 58530 46552 58586 46608
rect 1956 46266 2012 46268
rect 2036 46266 2092 46268
rect 2116 46266 2172 46268
rect 2196 46266 2252 46268
rect 1956 46214 2002 46266
rect 2002 46214 2012 46266
rect 2036 46214 2066 46266
rect 2066 46214 2078 46266
rect 2078 46214 2092 46266
rect 2116 46214 2130 46266
rect 2130 46214 2142 46266
rect 2142 46214 2172 46266
rect 2196 46214 2206 46266
rect 2206 46214 2252 46266
rect 1956 46212 2012 46214
rect 2036 46212 2092 46214
rect 2116 46212 2172 46214
rect 2196 46212 2252 46214
rect 6956 46266 7012 46268
rect 7036 46266 7092 46268
rect 7116 46266 7172 46268
rect 7196 46266 7252 46268
rect 6956 46214 7002 46266
rect 7002 46214 7012 46266
rect 7036 46214 7066 46266
rect 7066 46214 7078 46266
rect 7078 46214 7092 46266
rect 7116 46214 7130 46266
rect 7130 46214 7142 46266
rect 7142 46214 7172 46266
rect 7196 46214 7206 46266
rect 7206 46214 7252 46266
rect 6956 46212 7012 46214
rect 7036 46212 7092 46214
rect 7116 46212 7172 46214
rect 7196 46212 7252 46214
rect 11956 46266 12012 46268
rect 12036 46266 12092 46268
rect 12116 46266 12172 46268
rect 12196 46266 12252 46268
rect 11956 46214 12002 46266
rect 12002 46214 12012 46266
rect 12036 46214 12066 46266
rect 12066 46214 12078 46266
rect 12078 46214 12092 46266
rect 12116 46214 12130 46266
rect 12130 46214 12142 46266
rect 12142 46214 12172 46266
rect 12196 46214 12206 46266
rect 12206 46214 12252 46266
rect 11956 46212 12012 46214
rect 12036 46212 12092 46214
rect 12116 46212 12172 46214
rect 12196 46212 12252 46214
rect 16956 46266 17012 46268
rect 17036 46266 17092 46268
rect 17116 46266 17172 46268
rect 17196 46266 17252 46268
rect 16956 46214 17002 46266
rect 17002 46214 17012 46266
rect 17036 46214 17066 46266
rect 17066 46214 17078 46266
rect 17078 46214 17092 46266
rect 17116 46214 17130 46266
rect 17130 46214 17142 46266
rect 17142 46214 17172 46266
rect 17196 46214 17206 46266
rect 17206 46214 17252 46266
rect 16956 46212 17012 46214
rect 17036 46212 17092 46214
rect 17116 46212 17172 46214
rect 17196 46212 17252 46214
rect 21956 46266 22012 46268
rect 22036 46266 22092 46268
rect 22116 46266 22172 46268
rect 22196 46266 22252 46268
rect 21956 46214 22002 46266
rect 22002 46214 22012 46266
rect 22036 46214 22066 46266
rect 22066 46214 22078 46266
rect 22078 46214 22092 46266
rect 22116 46214 22130 46266
rect 22130 46214 22142 46266
rect 22142 46214 22172 46266
rect 22196 46214 22206 46266
rect 22206 46214 22252 46266
rect 21956 46212 22012 46214
rect 22036 46212 22092 46214
rect 22116 46212 22172 46214
rect 22196 46212 22252 46214
rect 26956 46266 27012 46268
rect 27036 46266 27092 46268
rect 27116 46266 27172 46268
rect 27196 46266 27252 46268
rect 26956 46214 27002 46266
rect 27002 46214 27012 46266
rect 27036 46214 27066 46266
rect 27066 46214 27078 46266
rect 27078 46214 27092 46266
rect 27116 46214 27130 46266
rect 27130 46214 27142 46266
rect 27142 46214 27172 46266
rect 27196 46214 27206 46266
rect 27206 46214 27252 46266
rect 26956 46212 27012 46214
rect 27036 46212 27092 46214
rect 27116 46212 27172 46214
rect 27196 46212 27252 46214
rect 31956 46266 32012 46268
rect 32036 46266 32092 46268
rect 32116 46266 32172 46268
rect 32196 46266 32252 46268
rect 31956 46214 32002 46266
rect 32002 46214 32012 46266
rect 32036 46214 32066 46266
rect 32066 46214 32078 46266
rect 32078 46214 32092 46266
rect 32116 46214 32130 46266
rect 32130 46214 32142 46266
rect 32142 46214 32172 46266
rect 32196 46214 32206 46266
rect 32206 46214 32252 46266
rect 31956 46212 32012 46214
rect 32036 46212 32092 46214
rect 32116 46212 32172 46214
rect 32196 46212 32252 46214
rect 36956 46266 37012 46268
rect 37036 46266 37092 46268
rect 37116 46266 37172 46268
rect 37196 46266 37252 46268
rect 36956 46214 37002 46266
rect 37002 46214 37012 46266
rect 37036 46214 37066 46266
rect 37066 46214 37078 46266
rect 37078 46214 37092 46266
rect 37116 46214 37130 46266
rect 37130 46214 37142 46266
rect 37142 46214 37172 46266
rect 37196 46214 37206 46266
rect 37206 46214 37252 46266
rect 36956 46212 37012 46214
rect 37036 46212 37092 46214
rect 37116 46212 37172 46214
rect 37196 46212 37252 46214
rect 41956 46266 42012 46268
rect 42036 46266 42092 46268
rect 42116 46266 42172 46268
rect 42196 46266 42252 46268
rect 41956 46214 42002 46266
rect 42002 46214 42012 46266
rect 42036 46214 42066 46266
rect 42066 46214 42078 46266
rect 42078 46214 42092 46266
rect 42116 46214 42130 46266
rect 42130 46214 42142 46266
rect 42142 46214 42172 46266
rect 42196 46214 42206 46266
rect 42206 46214 42252 46266
rect 41956 46212 42012 46214
rect 42036 46212 42092 46214
rect 42116 46212 42172 46214
rect 42196 46212 42252 46214
rect 46956 46266 47012 46268
rect 47036 46266 47092 46268
rect 47116 46266 47172 46268
rect 47196 46266 47252 46268
rect 46956 46214 47002 46266
rect 47002 46214 47012 46266
rect 47036 46214 47066 46266
rect 47066 46214 47078 46266
rect 47078 46214 47092 46266
rect 47116 46214 47130 46266
rect 47130 46214 47142 46266
rect 47142 46214 47172 46266
rect 47196 46214 47206 46266
rect 47206 46214 47252 46266
rect 46956 46212 47012 46214
rect 47036 46212 47092 46214
rect 47116 46212 47172 46214
rect 47196 46212 47252 46214
rect 51956 46266 52012 46268
rect 52036 46266 52092 46268
rect 52116 46266 52172 46268
rect 52196 46266 52252 46268
rect 51956 46214 52002 46266
rect 52002 46214 52012 46266
rect 52036 46214 52066 46266
rect 52066 46214 52078 46266
rect 52078 46214 52092 46266
rect 52116 46214 52130 46266
rect 52130 46214 52142 46266
rect 52142 46214 52172 46266
rect 52196 46214 52206 46266
rect 52206 46214 52252 46266
rect 51956 46212 52012 46214
rect 52036 46212 52092 46214
rect 52116 46212 52172 46214
rect 52196 46212 52252 46214
rect 56956 46266 57012 46268
rect 57036 46266 57092 46268
rect 57116 46266 57172 46268
rect 57196 46266 57252 46268
rect 56956 46214 57002 46266
rect 57002 46214 57012 46266
rect 57036 46214 57066 46266
rect 57066 46214 57078 46266
rect 57078 46214 57092 46266
rect 57116 46214 57130 46266
rect 57130 46214 57142 46266
rect 57142 46214 57172 46266
rect 57196 46214 57206 46266
rect 57206 46214 57252 46266
rect 56956 46212 57012 46214
rect 57036 46212 57092 46214
rect 57116 46212 57172 46214
rect 57196 46212 57252 46214
rect 58530 45736 58586 45792
rect 2616 45722 2672 45724
rect 2696 45722 2752 45724
rect 2776 45722 2832 45724
rect 2856 45722 2912 45724
rect 2616 45670 2662 45722
rect 2662 45670 2672 45722
rect 2696 45670 2726 45722
rect 2726 45670 2738 45722
rect 2738 45670 2752 45722
rect 2776 45670 2790 45722
rect 2790 45670 2802 45722
rect 2802 45670 2832 45722
rect 2856 45670 2866 45722
rect 2866 45670 2912 45722
rect 2616 45668 2672 45670
rect 2696 45668 2752 45670
rect 2776 45668 2832 45670
rect 2856 45668 2912 45670
rect 7616 45722 7672 45724
rect 7696 45722 7752 45724
rect 7776 45722 7832 45724
rect 7856 45722 7912 45724
rect 7616 45670 7662 45722
rect 7662 45670 7672 45722
rect 7696 45670 7726 45722
rect 7726 45670 7738 45722
rect 7738 45670 7752 45722
rect 7776 45670 7790 45722
rect 7790 45670 7802 45722
rect 7802 45670 7832 45722
rect 7856 45670 7866 45722
rect 7866 45670 7912 45722
rect 7616 45668 7672 45670
rect 7696 45668 7752 45670
rect 7776 45668 7832 45670
rect 7856 45668 7912 45670
rect 12616 45722 12672 45724
rect 12696 45722 12752 45724
rect 12776 45722 12832 45724
rect 12856 45722 12912 45724
rect 12616 45670 12662 45722
rect 12662 45670 12672 45722
rect 12696 45670 12726 45722
rect 12726 45670 12738 45722
rect 12738 45670 12752 45722
rect 12776 45670 12790 45722
rect 12790 45670 12802 45722
rect 12802 45670 12832 45722
rect 12856 45670 12866 45722
rect 12866 45670 12912 45722
rect 12616 45668 12672 45670
rect 12696 45668 12752 45670
rect 12776 45668 12832 45670
rect 12856 45668 12912 45670
rect 17616 45722 17672 45724
rect 17696 45722 17752 45724
rect 17776 45722 17832 45724
rect 17856 45722 17912 45724
rect 17616 45670 17662 45722
rect 17662 45670 17672 45722
rect 17696 45670 17726 45722
rect 17726 45670 17738 45722
rect 17738 45670 17752 45722
rect 17776 45670 17790 45722
rect 17790 45670 17802 45722
rect 17802 45670 17832 45722
rect 17856 45670 17866 45722
rect 17866 45670 17912 45722
rect 17616 45668 17672 45670
rect 17696 45668 17752 45670
rect 17776 45668 17832 45670
rect 17856 45668 17912 45670
rect 22616 45722 22672 45724
rect 22696 45722 22752 45724
rect 22776 45722 22832 45724
rect 22856 45722 22912 45724
rect 22616 45670 22662 45722
rect 22662 45670 22672 45722
rect 22696 45670 22726 45722
rect 22726 45670 22738 45722
rect 22738 45670 22752 45722
rect 22776 45670 22790 45722
rect 22790 45670 22802 45722
rect 22802 45670 22832 45722
rect 22856 45670 22866 45722
rect 22866 45670 22912 45722
rect 22616 45668 22672 45670
rect 22696 45668 22752 45670
rect 22776 45668 22832 45670
rect 22856 45668 22912 45670
rect 27616 45722 27672 45724
rect 27696 45722 27752 45724
rect 27776 45722 27832 45724
rect 27856 45722 27912 45724
rect 27616 45670 27662 45722
rect 27662 45670 27672 45722
rect 27696 45670 27726 45722
rect 27726 45670 27738 45722
rect 27738 45670 27752 45722
rect 27776 45670 27790 45722
rect 27790 45670 27802 45722
rect 27802 45670 27832 45722
rect 27856 45670 27866 45722
rect 27866 45670 27912 45722
rect 27616 45668 27672 45670
rect 27696 45668 27752 45670
rect 27776 45668 27832 45670
rect 27856 45668 27912 45670
rect 32616 45722 32672 45724
rect 32696 45722 32752 45724
rect 32776 45722 32832 45724
rect 32856 45722 32912 45724
rect 32616 45670 32662 45722
rect 32662 45670 32672 45722
rect 32696 45670 32726 45722
rect 32726 45670 32738 45722
rect 32738 45670 32752 45722
rect 32776 45670 32790 45722
rect 32790 45670 32802 45722
rect 32802 45670 32832 45722
rect 32856 45670 32866 45722
rect 32866 45670 32912 45722
rect 32616 45668 32672 45670
rect 32696 45668 32752 45670
rect 32776 45668 32832 45670
rect 32856 45668 32912 45670
rect 37616 45722 37672 45724
rect 37696 45722 37752 45724
rect 37776 45722 37832 45724
rect 37856 45722 37912 45724
rect 37616 45670 37662 45722
rect 37662 45670 37672 45722
rect 37696 45670 37726 45722
rect 37726 45670 37738 45722
rect 37738 45670 37752 45722
rect 37776 45670 37790 45722
rect 37790 45670 37802 45722
rect 37802 45670 37832 45722
rect 37856 45670 37866 45722
rect 37866 45670 37912 45722
rect 37616 45668 37672 45670
rect 37696 45668 37752 45670
rect 37776 45668 37832 45670
rect 37856 45668 37912 45670
rect 42616 45722 42672 45724
rect 42696 45722 42752 45724
rect 42776 45722 42832 45724
rect 42856 45722 42912 45724
rect 42616 45670 42662 45722
rect 42662 45670 42672 45722
rect 42696 45670 42726 45722
rect 42726 45670 42738 45722
rect 42738 45670 42752 45722
rect 42776 45670 42790 45722
rect 42790 45670 42802 45722
rect 42802 45670 42832 45722
rect 42856 45670 42866 45722
rect 42866 45670 42912 45722
rect 42616 45668 42672 45670
rect 42696 45668 42752 45670
rect 42776 45668 42832 45670
rect 42856 45668 42912 45670
rect 47616 45722 47672 45724
rect 47696 45722 47752 45724
rect 47776 45722 47832 45724
rect 47856 45722 47912 45724
rect 47616 45670 47662 45722
rect 47662 45670 47672 45722
rect 47696 45670 47726 45722
rect 47726 45670 47738 45722
rect 47738 45670 47752 45722
rect 47776 45670 47790 45722
rect 47790 45670 47802 45722
rect 47802 45670 47832 45722
rect 47856 45670 47866 45722
rect 47866 45670 47912 45722
rect 47616 45668 47672 45670
rect 47696 45668 47752 45670
rect 47776 45668 47832 45670
rect 47856 45668 47912 45670
rect 52616 45722 52672 45724
rect 52696 45722 52752 45724
rect 52776 45722 52832 45724
rect 52856 45722 52912 45724
rect 52616 45670 52662 45722
rect 52662 45670 52672 45722
rect 52696 45670 52726 45722
rect 52726 45670 52738 45722
rect 52738 45670 52752 45722
rect 52776 45670 52790 45722
rect 52790 45670 52802 45722
rect 52802 45670 52832 45722
rect 52856 45670 52866 45722
rect 52866 45670 52912 45722
rect 52616 45668 52672 45670
rect 52696 45668 52752 45670
rect 52776 45668 52832 45670
rect 52856 45668 52912 45670
rect 57616 45722 57672 45724
rect 57696 45722 57752 45724
rect 57776 45722 57832 45724
rect 57856 45722 57912 45724
rect 57616 45670 57662 45722
rect 57662 45670 57672 45722
rect 57696 45670 57726 45722
rect 57726 45670 57738 45722
rect 57738 45670 57752 45722
rect 57776 45670 57790 45722
rect 57790 45670 57802 45722
rect 57802 45670 57832 45722
rect 57856 45670 57866 45722
rect 57866 45670 57912 45722
rect 57616 45668 57672 45670
rect 57696 45668 57752 45670
rect 57776 45668 57832 45670
rect 57856 45668 57912 45670
rect 1956 45178 2012 45180
rect 2036 45178 2092 45180
rect 2116 45178 2172 45180
rect 2196 45178 2252 45180
rect 1956 45126 2002 45178
rect 2002 45126 2012 45178
rect 2036 45126 2066 45178
rect 2066 45126 2078 45178
rect 2078 45126 2092 45178
rect 2116 45126 2130 45178
rect 2130 45126 2142 45178
rect 2142 45126 2172 45178
rect 2196 45126 2206 45178
rect 2206 45126 2252 45178
rect 1956 45124 2012 45126
rect 2036 45124 2092 45126
rect 2116 45124 2172 45126
rect 2196 45124 2252 45126
rect 6956 45178 7012 45180
rect 7036 45178 7092 45180
rect 7116 45178 7172 45180
rect 7196 45178 7252 45180
rect 6956 45126 7002 45178
rect 7002 45126 7012 45178
rect 7036 45126 7066 45178
rect 7066 45126 7078 45178
rect 7078 45126 7092 45178
rect 7116 45126 7130 45178
rect 7130 45126 7142 45178
rect 7142 45126 7172 45178
rect 7196 45126 7206 45178
rect 7206 45126 7252 45178
rect 6956 45124 7012 45126
rect 7036 45124 7092 45126
rect 7116 45124 7172 45126
rect 7196 45124 7252 45126
rect 11956 45178 12012 45180
rect 12036 45178 12092 45180
rect 12116 45178 12172 45180
rect 12196 45178 12252 45180
rect 11956 45126 12002 45178
rect 12002 45126 12012 45178
rect 12036 45126 12066 45178
rect 12066 45126 12078 45178
rect 12078 45126 12092 45178
rect 12116 45126 12130 45178
rect 12130 45126 12142 45178
rect 12142 45126 12172 45178
rect 12196 45126 12206 45178
rect 12206 45126 12252 45178
rect 11956 45124 12012 45126
rect 12036 45124 12092 45126
rect 12116 45124 12172 45126
rect 12196 45124 12252 45126
rect 16956 45178 17012 45180
rect 17036 45178 17092 45180
rect 17116 45178 17172 45180
rect 17196 45178 17252 45180
rect 16956 45126 17002 45178
rect 17002 45126 17012 45178
rect 17036 45126 17066 45178
rect 17066 45126 17078 45178
rect 17078 45126 17092 45178
rect 17116 45126 17130 45178
rect 17130 45126 17142 45178
rect 17142 45126 17172 45178
rect 17196 45126 17206 45178
rect 17206 45126 17252 45178
rect 16956 45124 17012 45126
rect 17036 45124 17092 45126
rect 17116 45124 17172 45126
rect 17196 45124 17252 45126
rect 21956 45178 22012 45180
rect 22036 45178 22092 45180
rect 22116 45178 22172 45180
rect 22196 45178 22252 45180
rect 21956 45126 22002 45178
rect 22002 45126 22012 45178
rect 22036 45126 22066 45178
rect 22066 45126 22078 45178
rect 22078 45126 22092 45178
rect 22116 45126 22130 45178
rect 22130 45126 22142 45178
rect 22142 45126 22172 45178
rect 22196 45126 22206 45178
rect 22206 45126 22252 45178
rect 21956 45124 22012 45126
rect 22036 45124 22092 45126
rect 22116 45124 22172 45126
rect 22196 45124 22252 45126
rect 26956 45178 27012 45180
rect 27036 45178 27092 45180
rect 27116 45178 27172 45180
rect 27196 45178 27252 45180
rect 26956 45126 27002 45178
rect 27002 45126 27012 45178
rect 27036 45126 27066 45178
rect 27066 45126 27078 45178
rect 27078 45126 27092 45178
rect 27116 45126 27130 45178
rect 27130 45126 27142 45178
rect 27142 45126 27172 45178
rect 27196 45126 27206 45178
rect 27206 45126 27252 45178
rect 26956 45124 27012 45126
rect 27036 45124 27092 45126
rect 27116 45124 27172 45126
rect 27196 45124 27252 45126
rect 31956 45178 32012 45180
rect 32036 45178 32092 45180
rect 32116 45178 32172 45180
rect 32196 45178 32252 45180
rect 31956 45126 32002 45178
rect 32002 45126 32012 45178
rect 32036 45126 32066 45178
rect 32066 45126 32078 45178
rect 32078 45126 32092 45178
rect 32116 45126 32130 45178
rect 32130 45126 32142 45178
rect 32142 45126 32172 45178
rect 32196 45126 32206 45178
rect 32206 45126 32252 45178
rect 31956 45124 32012 45126
rect 32036 45124 32092 45126
rect 32116 45124 32172 45126
rect 32196 45124 32252 45126
rect 36956 45178 37012 45180
rect 37036 45178 37092 45180
rect 37116 45178 37172 45180
rect 37196 45178 37252 45180
rect 36956 45126 37002 45178
rect 37002 45126 37012 45178
rect 37036 45126 37066 45178
rect 37066 45126 37078 45178
rect 37078 45126 37092 45178
rect 37116 45126 37130 45178
rect 37130 45126 37142 45178
rect 37142 45126 37172 45178
rect 37196 45126 37206 45178
rect 37206 45126 37252 45178
rect 36956 45124 37012 45126
rect 37036 45124 37092 45126
rect 37116 45124 37172 45126
rect 37196 45124 37252 45126
rect 41956 45178 42012 45180
rect 42036 45178 42092 45180
rect 42116 45178 42172 45180
rect 42196 45178 42252 45180
rect 41956 45126 42002 45178
rect 42002 45126 42012 45178
rect 42036 45126 42066 45178
rect 42066 45126 42078 45178
rect 42078 45126 42092 45178
rect 42116 45126 42130 45178
rect 42130 45126 42142 45178
rect 42142 45126 42172 45178
rect 42196 45126 42206 45178
rect 42206 45126 42252 45178
rect 41956 45124 42012 45126
rect 42036 45124 42092 45126
rect 42116 45124 42172 45126
rect 42196 45124 42252 45126
rect 46956 45178 47012 45180
rect 47036 45178 47092 45180
rect 47116 45178 47172 45180
rect 47196 45178 47252 45180
rect 46956 45126 47002 45178
rect 47002 45126 47012 45178
rect 47036 45126 47066 45178
rect 47066 45126 47078 45178
rect 47078 45126 47092 45178
rect 47116 45126 47130 45178
rect 47130 45126 47142 45178
rect 47142 45126 47172 45178
rect 47196 45126 47206 45178
rect 47206 45126 47252 45178
rect 46956 45124 47012 45126
rect 47036 45124 47092 45126
rect 47116 45124 47172 45126
rect 47196 45124 47252 45126
rect 51956 45178 52012 45180
rect 52036 45178 52092 45180
rect 52116 45178 52172 45180
rect 52196 45178 52252 45180
rect 51956 45126 52002 45178
rect 52002 45126 52012 45178
rect 52036 45126 52066 45178
rect 52066 45126 52078 45178
rect 52078 45126 52092 45178
rect 52116 45126 52130 45178
rect 52130 45126 52142 45178
rect 52142 45126 52172 45178
rect 52196 45126 52206 45178
rect 52206 45126 52252 45178
rect 51956 45124 52012 45126
rect 52036 45124 52092 45126
rect 52116 45124 52172 45126
rect 52196 45124 52252 45126
rect 56956 45178 57012 45180
rect 57036 45178 57092 45180
rect 57116 45178 57172 45180
rect 57196 45178 57252 45180
rect 56956 45126 57002 45178
rect 57002 45126 57012 45178
rect 57036 45126 57066 45178
rect 57066 45126 57078 45178
rect 57078 45126 57092 45178
rect 57116 45126 57130 45178
rect 57130 45126 57142 45178
rect 57142 45126 57172 45178
rect 57196 45126 57206 45178
rect 57206 45126 57252 45178
rect 56956 45124 57012 45126
rect 57036 45124 57092 45126
rect 57116 45124 57172 45126
rect 57196 45124 57252 45126
rect 58530 44920 58586 44976
rect 2616 44634 2672 44636
rect 2696 44634 2752 44636
rect 2776 44634 2832 44636
rect 2856 44634 2912 44636
rect 2616 44582 2662 44634
rect 2662 44582 2672 44634
rect 2696 44582 2726 44634
rect 2726 44582 2738 44634
rect 2738 44582 2752 44634
rect 2776 44582 2790 44634
rect 2790 44582 2802 44634
rect 2802 44582 2832 44634
rect 2856 44582 2866 44634
rect 2866 44582 2912 44634
rect 2616 44580 2672 44582
rect 2696 44580 2752 44582
rect 2776 44580 2832 44582
rect 2856 44580 2912 44582
rect 7616 44634 7672 44636
rect 7696 44634 7752 44636
rect 7776 44634 7832 44636
rect 7856 44634 7912 44636
rect 7616 44582 7662 44634
rect 7662 44582 7672 44634
rect 7696 44582 7726 44634
rect 7726 44582 7738 44634
rect 7738 44582 7752 44634
rect 7776 44582 7790 44634
rect 7790 44582 7802 44634
rect 7802 44582 7832 44634
rect 7856 44582 7866 44634
rect 7866 44582 7912 44634
rect 7616 44580 7672 44582
rect 7696 44580 7752 44582
rect 7776 44580 7832 44582
rect 7856 44580 7912 44582
rect 12616 44634 12672 44636
rect 12696 44634 12752 44636
rect 12776 44634 12832 44636
rect 12856 44634 12912 44636
rect 12616 44582 12662 44634
rect 12662 44582 12672 44634
rect 12696 44582 12726 44634
rect 12726 44582 12738 44634
rect 12738 44582 12752 44634
rect 12776 44582 12790 44634
rect 12790 44582 12802 44634
rect 12802 44582 12832 44634
rect 12856 44582 12866 44634
rect 12866 44582 12912 44634
rect 12616 44580 12672 44582
rect 12696 44580 12752 44582
rect 12776 44580 12832 44582
rect 12856 44580 12912 44582
rect 17616 44634 17672 44636
rect 17696 44634 17752 44636
rect 17776 44634 17832 44636
rect 17856 44634 17912 44636
rect 17616 44582 17662 44634
rect 17662 44582 17672 44634
rect 17696 44582 17726 44634
rect 17726 44582 17738 44634
rect 17738 44582 17752 44634
rect 17776 44582 17790 44634
rect 17790 44582 17802 44634
rect 17802 44582 17832 44634
rect 17856 44582 17866 44634
rect 17866 44582 17912 44634
rect 17616 44580 17672 44582
rect 17696 44580 17752 44582
rect 17776 44580 17832 44582
rect 17856 44580 17912 44582
rect 22616 44634 22672 44636
rect 22696 44634 22752 44636
rect 22776 44634 22832 44636
rect 22856 44634 22912 44636
rect 22616 44582 22662 44634
rect 22662 44582 22672 44634
rect 22696 44582 22726 44634
rect 22726 44582 22738 44634
rect 22738 44582 22752 44634
rect 22776 44582 22790 44634
rect 22790 44582 22802 44634
rect 22802 44582 22832 44634
rect 22856 44582 22866 44634
rect 22866 44582 22912 44634
rect 22616 44580 22672 44582
rect 22696 44580 22752 44582
rect 22776 44580 22832 44582
rect 22856 44580 22912 44582
rect 27616 44634 27672 44636
rect 27696 44634 27752 44636
rect 27776 44634 27832 44636
rect 27856 44634 27912 44636
rect 27616 44582 27662 44634
rect 27662 44582 27672 44634
rect 27696 44582 27726 44634
rect 27726 44582 27738 44634
rect 27738 44582 27752 44634
rect 27776 44582 27790 44634
rect 27790 44582 27802 44634
rect 27802 44582 27832 44634
rect 27856 44582 27866 44634
rect 27866 44582 27912 44634
rect 27616 44580 27672 44582
rect 27696 44580 27752 44582
rect 27776 44580 27832 44582
rect 27856 44580 27912 44582
rect 32616 44634 32672 44636
rect 32696 44634 32752 44636
rect 32776 44634 32832 44636
rect 32856 44634 32912 44636
rect 32616 44582 32662 44634
rect 32662 44582 32672 44634
rect 32696 44582 32726 44634
rect 32726 44582 32738 44634
rect 32738 44582 32752 44634
rect 32776 44582 32790 44634
rect 32790 44582 32802 44634
rect 32802 44582 32832 44634
rect 32856 44582 32866 44634
rect 32866 44582 32912 44634
rect 32616 44580 32672 44582
rect 32696 44580 32752 44582
rect 32776 44580 32832 44582
rect 32856 44580 32912 44582
rect 37616 44634 37672 44636
rect 37696 44634 37752 44636
rect 37776 44634 37832 44636
rect 37856 44634 37912 44636
rect 37616 44582 37662 44634
rect 37662 44582 37672 44634
rect 37696 44582 37726 44634
rect 37726 44582 37738 44634
rect 37738 44582 37752 44634
rect 37776 44582 37790 44634
rect 37790 44582 37802 44634
rect 37802 44582 37832 44634
rect 37856 44582 37866 44634
rect 37866 44582 37912 44634
rect 37616 44580 37672 44582
rect 37696 44580 37752 44582
rect 37776 44580 37832 44582
rect 37856 44580 37912 44582
rect 42616 44634 42672 44636
rect 42696 44634 42752 44636
rect 42776 44634 42832 44636
rect 42856 44634 42912 44636
rect 42616 44582 42662 44634
rect 42662 44582 42672 44634
rect 42696 44582 42726 44634
rect 42726 44582 42738 44634
rect 42738 44582 42752 44634
rect 42776 44582 42790 44634
rect 42790 44582 42802 44634
rect 42802 44582 42832 44634
rect 42856 44582 42866 44634
rect 42866 44582 42912 44634
rect 42616 44580 42672 44582
rect 42696 44580 42752 44582
rect 42776 44580 42832 44582
rect 42856 44580 42912 44582
rect 47616 44634 47672 44636
rect 47696 44634 47752 44636
rect 47776 44634 47832 44636
rect 47856 44634 47912 44636
rect 47616 44582 47662 44634
rect 47662 44582 47672 44634
rect 47696 44582 47726 44634
rect 47726 44582 47738 44634
rect 47738 44582 47752 44634
rect 47776 44582 47790 44634
rect 47790 44582 47802 44634
rect 47802 44582 47832 44634
rect 47856 44582 47866 44634
rect 47866 44582 47912 44634
rect 47616 44580 47672 44582
rect 47696 44580 47752 44582
rect 47776 44580 47832 44582
rect 47856 44580 47912 44582
rect 52616 44634 52672 44636
rect 52696 44634 52752 44636
rect 52776 44634 52832 44636
rect 52856 44634 52912 44636
rect 52616 44582 52662 44634
rect 52662 44582 52672 44634
rect 52696 44582 52726 44634
rect 52726 44582 52738 44634
rect 52738 44582 52752 44634
rect 52776 44582 52790 44634
rect 52790 44582 52802 44634
rect 52802 44582 52832 44634
rect 52856 44582 52866 44634
rect 52866 44582 52912 44634
rect 52616 44580 52672 44582
rect 52696 44580 52752 44582
rect 52776 44580 52832 44582
rect 52856 44580 52912 44582
rect 57616 44634 57672 44636
rect 57696 44634 57752 44636
rect 57776 44634 57832 44636
rect 57856 44634 57912 44636
rect 57616 44582 57662 44634
rect 57662 44582 57672 44634
rect 57696 44582 57726 44634
rect 57726 44582 57738 44634
rect 57738 44582 57752 44634
rect 57776 44582 57790 44634
rect 57790 44582 57802 44634
rect 57802 44582 57832 44634
rect 57856 44582 57866 44634
rect 57866 44582 57912 44634
rect 57616 44580 57672 44582
rect 57696 44580 57752 44582
rect 57776 44580 57832 44582
rect 57856 44580 57912 44582
rect 58530 44140 58532 44160
rect 58532 44140 58584 44160
rect 58584 44140 58586 44160
rect 58530 44104 58586 44140
rect 1956 44090 2012 44092
rect 2036 44090 2092 44092
rect 2116 44090 2172 44092
rect 2196 44090 2252 44092
rect 1956 44038 2002 44090
rect 2002 44038 2012 44090
rect 2036 44038 2066 44090
rect 2066 44038 2078 44090
rect 2078 44038 2092 44090
rect 2116 44038 2130 44090
rect 2130 44038 2142 44090
rect 2142 44038 2172 44090
rect 2196 44038 2206 44090
rect 2206 44038 2252 44090
rect 1956 44036 2012 44038
rect 2036 44036 2092 44038
rect 2116 44036 2172 44038
rect 2196 44036 2252 44038
rect 6956 44090 7012 44092
rect 7036 44090 7092 44092
rect 7116 44090 7172 44092
rect 7196 44090 7252 44092
rect 6956 44038 7002 44090
rect 7002 44038 7012 44090
rect 7036 44038 7066 44090
rect 7066 44038 7078 44090
rect 7078 44038 7092 44090
rect 7116 44038 7130 44090
rect 7130 44038 7142 44090
rect 7142 44038 7172 44090
rect 7196 44038 7206 44090
rect 7206 44038 7252 44090
rect 6956 44036 7012 44038
rect 7036 44036 7092 44038
rect 7116 44036 7172 44038
rect 7196 44036 7252 44038
rect 11956 44090 12012 44092
rect 12036 44090 12092 44092
rect 12116 44090 12172 44092
rect 12196 44090 12252 44092
rect 11956 44038 12002 44090
rect 12002 44038 12012 44090
rect 12036 44038 12066 44090
rect 12066 44038 12078 44090
rect 12078 44038 12092 44090
rect 12116 44038 12130 44090
rect 12130 44038 12142 44090
rect 12142 44038 12172 44090
rect 12196 44038 12206 44090
rect 12206 44038 12252 44090
rect 11956 44036 12012 44038
rect 12036 44036 12092 44038
rect 12116 44036 12172 44038
rect 12196 44036 12252 44038
rect 16956 44090 17012 44092
rect 17036 44090 17092 44092
rect 17116 44090 17172 44092
rect 17196 44090 17252 44092
rect 16956 44038 17002 44090
rect 17002 44038 17012 44090
rect 17036 44038 17066 44090
rect 17066 44038 17078 44090
rect 17078 44038 17092 44090
rect 17116 44038 17130 44090
rect 17130 44038 17142 44090
rect 17142 44038 17172 44090
rect 17196 44038 17206 44090
rect 17206 44038 17252 44090
rect 16956 44036 17012 44038
rect 17036 44036 17092 44038
rect 17116 44036 17172 44038
rect 17196 44036 17252 44038
rect 21956 44090 22012 44092
rect 22036 44090 22092 44092
rect 22116 44090 22172 44092
rect 22196 44090 22252 44092
rect 21956 44038 22002 44090
rect 22002 44038 22012 44090
rect 22036 44038 22066 44090
rect 22066 44038 22078 44090
rect 22078 44038 22092 44090
rect 22116 44038 22130 44090
rect 22130 44038 22142 44090
rect 22142 44038 22172 44090
rect 22196 44038 22206 44090
rect 22206 44038 22252 44090
rect 21956 44036 22012 44038
rect 22036 44036 22092 44038
rect 22116 44036 22172 44038
rect 22196 44036 22252 44038
rect 26956 44090 27012 44092
rect 27036 44090 27092 44092
rect 27116 44090 27172 44092
rect 27196 44090 27252 44092
rect 26956 44038 27002 44090
rect 27002 44038 27012 44090
rect 27036 44038 27066 44090
rect 27066 44038 27078 44090
rect 27078 44038 27092 44090
rect 27116 44038 27130 44090
rect 27130 44038 27142 44090
rect 27142 44038 27172 44090
rect 27196 44038 27206 44090
rect 27206 44038 27252 44090
rect 26956 44036 27012 44038
rect 27036 44036 27092 44038
rect 27116 44036 27172 44038
rect 27196 44036 27252 44038
rect 31956 44090 32012 44092
rect 32036 44090 32092 44092
rect 32116 44090 32172 44092
rect 32196 44090 32252 44092
rect 31956 44038 32002 44090
rect 32002 44038 32012 44090
rect 32036 44038 32066 44090
rect 32066 44038 32078 44090
rect 32078 44038 32092 44090
rect 32116 44038 32130 44090
rect 32130 44038 32142 44090
rect 32142 44038 32172 44090
rect 32196 44038 32206 44090
rect 32206 44038 32252 44090
rect 31956 44036 32012 44038
rect 32036 44036 32092 44038
rect 32116 44036 32172 44038
rect 32196 44036 32252 44038
rect 36956 44090 37012 44092
rect 37036 44090 37092 44092
rect 37116 44090 37172 44092
rect 37196 44090 37252 44092
rect 36956 44038 37002 44090
rect 37002 44038 37012 44090
rect 37036 44038 37066 44090
rect 37066 44038 37078 44090
rect 37078 44038 37092 44090
rect 37116 44038 37130 44090
rect 37130 44038 37142 44090
rect 37142 44038 37172 44090
rect 37196 44038 37206 44090
rect 37206 44038 37252 44090
rect 36956 44036 37012 44038
rect 37036 44036 37092 44038
rect 37116 44036 37172 44038
rect 37196 44036 37252 44038
rect 41956 44090 42012 44092
rect 42036 44090 42092 44092
rect 42116 44090 42172 44092
rect 42196 44090 42252 44092
rect 41956 44038 42002 44090
rect 42002 44038 42012 44090
rect 42036 44038 42066 44090
rect 42066 44038 42078 44090
rect 42078 44038 42092 44090
rect 42116 44038 42130 44090
rect 42130 44038 42142 44090
rect 42142 44038 42172 44090
rect 42196 44038 42206 44090
rect 42206 44038 42252 44090
rect 41956 44036 42012 44038
rect 42036 44036 42092 44038
rect 42116 44036 42172 44038
rect 42196 44036 42252 44038
rect 46956 44090 47012 44092
rect 47036 44090 47092 44092
rect 47116 44090 47172 44092
rect 47196 44090 47252 44092
rect 46956 44038 47002 44090
rect 47002 44038 47012 44090
rect 47036 44038 47066 44090
rect 47066 44038 47078 44090
rect 47078 44038 47092 44090
rect 47116 44038 47130 44090
rect 47130 44038 47142 44090
rect 47142 44038 47172 44090
rect 47196 44038 47206 44090
rect 47206 44038 47252 44090
rect 46956 44036 47012 44038
rect 47036 44036 47092 44038
rect 47116 44036 47172 44038
rect 47196 44036 47252 44038
rect 51956 44090 52012 44092
rect 52036 44090 52092 44092
rect 52116 44090 52172 44092
rect 52196 44090 52252 44092
rect 51956 44038 52002 44090
rect 52002 44038 52012 44090
rect 52036 44038 52066 44090
rect 52066 44038 52078 44090
rect 52078 44038 52092 44090
rect 52116 44038 52130 44090
rect 52130 44038 52142 44090
rect 52142 44038 52172 44090
rect 52196 44038 52206 44090
rect 52206 44038 52252 44090
rect 51956 44036 52012 44038
rect 52036 44036 52092 44038
rect 52116 44036 52172 44038
rect 52196 44036 52252 44038
rect 56956 44090 57012 44092
rect 57036 44090 57092 44092
rect 57116 44090 57172 44092
rect 57196 44090 57252 44092
rect 56956 44038 57002 44090
rect 57002 44038 57012 44090
rect 57036 44038 57066 44090
rect 57066 44038 57078 44090
rect 57078 44038 57092 44090
rect 57116 44038 57130 44090
rect 57130 44038 57142 44090
rect 57142 44038 57172 44090
rect 57196 44038 57206 44090
rect 57206 44038 57252 44090
rect 56956 44036 57012 44038
rect 57036 44036 57092 44038
rect 57116 44036 57172 44038
rect 57196 44036 57252 44038
rect 2616 43546 2672 43548
rect 2696 43546 2752 43548
rect 2776 43546 2832 43548
rect 2856 43546 2912 43548
rect 2616 43494 2662 43546
rect 2662 43494 2672 43546
rect 2696 43494 2726 43546
rect 2726 43494 2738 43546
rect 2738 43494 2752 43546
rect 2776 43494 2790 43546
rect 2790 43494 2802 43546
rect 2802 43494 2832 43546
rect 2856 43494 2866 43546
rect 2866 43494 2912 43546
rect 2616 43492 2672 43494
rect 2696 43492 2752 43494
rect 2776 43492 2832 43494
rect 2856 43492 2912 43494
rect 7616 43546 7672 43548
rect 7696 43546 7752 43548
rect 7776 43546 7832 43548
rect 7856 43546 7912 43548
rect 7616 43494 7662 43546
rect 7662 43494 7672 43546
rect 7696 43494 7726 43546
rect 7726 43494 7738 43546
rect 7738 43494 7752 43546
rect 7776 43494 7790 43546
rect 7790 43494 7802 43546
rect 7802 43494 7832 43546
rect 7856 43494 7866 43546
rect 7866 43494 7912 43546
rect 7616 43492 7672 43494
rect 7696 43492 7752 43494
rect 7776 43492 7832 43494
rect 7856 43492 7912 43494
rect 12616 43546 12672 43548
rect 12696 43546 12752 43548
rect 12776 43546 12832 43548
rect 12856 43546 12912 43548
rect 12616 43494 12662 43546
rect 12662 43494 12672 43546
rect 12696 43494 12726 43546
rect 12726 43494 12738 43546
rect 12738 43494 12752 43546
rect 12776 43494 12790 43546
rect 12790 43494 12802 43546
rect 12802 43494 12832 43546
rect 12856 43494 12866 43546
rect 12866 43494 12912 43546
rect 12616 43492 12672 43494
rect 12696 43492 12752 43494
rect 12776 43492 12832 43494
rect 12856 43492 12912 43494
rect 17616 43546 17672 43548
rect 17696 43546 17752 43548
rect 17776 43546 17832 43548
rect 17856 43546 17912 43548
rect 17616 43494 17662 43546
rect 17662 43494 17672 43546
rect 17696 43494 17726 43546
rect 17726 43494 17738 43546
rect 17738 43494 17752 43546
rect 17776 43494 17790 43546
rect 17790 43494 17802 43546
rect 17802 43494 17832 43546
rect 17856 43494 17866 43546
rect 17866 43494 17912 43546
rect 17616 43492 17672 43494
rect 17696 43492 17752 43494
rect 17776 43492 17832 43494
rect 17856 43492 17912 43494
rect 22616 43546 22672 43548
rect 22696 43546 22752 43548
rect 22776 43546 22832 43548
rect 22856 43546 22912 43548
rect 22616 43494 22662 43546
rect 22662 43494 22672 43546
rect 22696 43494 22726 43546
rect 22726 43494 22738 43546
rect 22738 43494 22752 43546
rect 22776 43494 22790 43546
rect 22790 43494 22802 43546
rect 22802 43494 22832 43546
rect 22856 43494 22866 43546
rect 22866 43494 22912 43546
rect 22616 43492 22672 43494
rect 22696 43492 22752 43494
rect 22776 43492 22832 43494
rect 22856 43492 22912 43494
rect 27616 43546 27672 43548
rect 27696 43546 27752 43548
rect 27776 43546 27832 43548
rect 27856 43546 27912 43548
rect 27616 43494 27662 43546
rect 27662 43494 27672 43546
rect 27696 43494 27726 43546
rect 27726 43494 27738 43546
rect 27738 43494 27752 43546
rect 27776 43494 27790 43546
rect 27790 43494 27802 43546
rect 27802 43494 27832 43546
rect 27856 43494 27866 43546
rect 27866 43494 27912 43546
rect 27616 43492 27672 43494
rect 27696 43492 27752 43494
rect 27776 43492 27832 43494
rect 27856 43492 27912 43494
rect 32616 43546 32672 43548
rect 32696 43546 32752 43548
rect 32776 43546 32832 43548
rect 32856 43546 32912 43548
rect 32616 43494 32662 43546
rect 32662 43494 32672 43546
rect 32696 43494 32726 43546
rect 32726 43494 32738 43546
rect 32738 43494 32752 43546
rect 32776 43494 32790 43546
rect 32790 43494 32802 43546
rect 32802 43494 32832 43546
rect 32856 43494 32866 43546
rect 32866 43494 32912 43546
rect 32616 43492 32672 43494
rect 32696 43492 32752 43494
rect 32776 43492 32832 43494
rect 32856 43492 32912 43494
rect 37616 43546 37672 43548
rect 37696 43546 37752 43548
rect 37776 43546 37832 43548
rect 37856 43546 37912 43548
rect 37616 43494 37662 43546
rect 37662 43494 37672 43546
rect 37696 43494 37726 43546
rect 37726 43494 37738 43546
rect 37738 43494 37752 43546
rect 37776 43494 37790 43546
rect 37790 43494 37802 43546
rect 37802 43494 37832 43546
rect 37856 43494 37866 43546
rect 37866 43494 37912 43546
rect 37616 43492 37672 43494
rect 37696 43492 37752 43494
rect 37776 43492 37832 43494
rect 37856 43492 37912 43494
rect 42616 43546 42672 43548
rect 42696 43546 42752 43548
rect 42776 43546 42832 43548
rect 42856 43546 42912 43548
rect 42616 43494 42662 43546
rect 42662 43494 42672 43546
rect 42696 43494 42726 43546
rect 42726 43494 42738 43546
rect 42738 43494 42752 43546
rect 42776 43494 42790 43546
rect 42790 43494 42802 43546
rect 42802 43494 42832 43546
rect 42856 43494 42866 43546
rect 42866 43494 42912 43546
rect 42616 43492 42672 43494
rect 42696 43492 42752 43494
rect 42776 43492 42832 43494
rect 42856 43492 42912 43494
rect 47616 43546 47672 43548
rect 47696 43546 47752 43548
rect 47776 43546 47832 43548
rect 47856 43546 47912 43548
rect 47616 43494 47662 43546
rect 47662 43494 47672 43546
rect 47696 43494 47726 43546
rect 47726 43494 47738 43546
rect 47738 43494 47752 43546
rect 47776 43494 47790 43546
rect 47790 43494 47802 43546
rect 47802 43494 47832 43546
rect 47856 43494 47866 43546
rect 47866 43494 47912 43546
rect 47616 43492 47672 43494
rect 47696 43492 47752 43494
rect 47776 43492 47832 43494
rect 47856 43492 47912 43494
rect 52616 43546 52672 43548
rect 52696 43546 52752 43548
rect 52776 43546 52832 43548
rect 52856 43546 52912 43548
rect 52616 43494 52662 43546
rect 52662 43494 52672 43546
rect 52696 43494 52726 43546
rect 52726 43494 52738 43546
rect 52738 43494 52752 43546
rect 52776 43494 52790 43546
rect 52790 43494 52802 43546
rect 52802 43494 52832 43546
rect 52856 43494 52866 43546
rect 52866 43494 52912 43546
rect 52616 43492 52672 43494
rect 52696 43492 52752 43494
rect 52776 43492 52832 43494
rect 52856 43492 52912 43494
rect 57616 43546 57672 43548
rect 57696 43546 57752 43548
rect 57776 43546 57832 43548
rect 57856 43546 57912 43548
rect 57616 43494 57662 43546
rect 57662 43494 57672 43546
rect 57696 43494 57726 43546
rect 57726 43494 57738 43546
rect 57738 43494 57752 43546
rect 57776 43494 57790 43546
rect 57790 43494 57802 43546
rect 57802 43494 57832 43546
rect 57856 43494 57866 43546
rect 57866 43494 57912 43546
rect 57616 43492 57672 43494
rect 57696 43492 57752 43494
rect 57776 43492 57832 43494
rect 57856 43492 57912 43494
rect 58530 43288 58586 43344
rect 1956 43002 2012 43004
rect 2036 43002 2092 43004
rect 2116 43002 2172 43004
rect 2196 43002 2252 43004
rect 1956 42950 2002 43002
rect 2002 42950 2012 43002
rect 2036 42950 2066 43002
rect 2066 42950 2078 43002
rect 2078 42950 2092 43002
rect 2116 42950 2130 43002
rect 2130 42950 2142 43002
rect 2142 42950 2172 43002
rect 2196 42950 2206 43002
rect 2206 42950 2252 43002
rect 1956 42948 2012 42950
rect 2036 42948 2092 42950
rect 2116 42948 2172 42950
rect 2196 42948 2252 42950
rect 6956 43002 7012 43004
rect 7036 43002 7092 43004
rect 7116 43002 7172 43004
rect 7196 43002 7252 43004
rect 6956 42950 7002 43002
rect 7002 42950 7012 43002
rect 7036 42950 7066 43002
rect 7066 42950 7078 43002
rect 7078 42950 7092 43002
rect 7116 42950 7130 43002
rect 7130 42950 7142 43002
rect 7142 42950 7172 43002
rect 7196 42950 7206 43002
rect 7206 42950 7252 43002
rect 6956 42948 7012 42950
rect 7036 42948 7092 42950
rect 7116 42948 7172 42950
rect 7196 42948 7252 42950
rect 11956 43002 12012 43004
rect 12036 43002 12092 43004
rect 12116 43002 12172 43004
rect 12196 43002 12252 43004
rect 11956 42950 12002 43002
rect 12002 42950 12012 43002
rect 12036 42950 12066 43002
rect 12066 42950 12078 43002
rect 12078 42950 12092 43002
rect 12116 42950 12130 43002
rect 12130 42950 12142 43002
rect 12142 42950 12172 43002
rect 12196 42950 12206 43002
rect 12206 42950 12252 43002
rect 11956 42948 12012 42950
rect 12036 42948 12092 42950
rect 12116 42948 12172 42950
rect 12196 42948 12252 42950
rect 16956 43002 17012 43004
rect 17036 43002 17092 43004
rect 17116 43002 17172 43004
rect 17196 43002 17252 43004
rect 16956 42950 17002 43002
rect 17002 42950 17012 43002
rect 17036 42950 17066 43002
rect 17066 42950 17078 43002
rect 17078 42950 17092 43002
rect 17116 42950 17130 43002
rect 17130 42950 17142 43002
rect 17142 42950 17172 43002
rect 17196 42950 17206 43002
rect 17206 42950 17252 43002
rect 16956 42948 17012 42950
rect 17036 42948 17092 42950
rect 17116 42948 17172 42950
rect 17196 42948 17252 42950
rect 21956 43002 22012 43004
rect 22036 43002 22092 43004
rect 22116 43002 22172 43004
rect 22196 43002 22252 43004
rect 21956 42950 22002 43002
rect 22002 42950 22012 43002
rect 22036 42950 22066 43002
rect 22066 42950 22078 43002
rect 22078 42950 22092 43002
rect 22116 42950 22130 43002
rect 22130 42950 22142 43002
rect 22142 42950 22172 43002
rect 22196 42950 22206 43002
rect 22206 42950 22252 43002
rect 21956 42948 22012 42950
rect 22036 42948 22092 42950
rect 22116 42948 22172 42950
rect 22196 42948 22252 42950
rect 26956 43002 27012 43004
rect 27036 43002 27092 43004
rect 27116 43002 27172 43004
rect 27196 43002 27252 43004
rect 26956 42950 27002 43002
rect 27002 42950 27012 43002
rect 27036 42950 27066 43002
rect 27066 42950 27078 43002
rect 27078 42950 27092 43002
rect 27116 42950 27130 43002
rect 27130 42950 27142 43002
rect 27142 42950 27172 43002
rect 27196 42950 27206 43002
rect 27206 42950 27252 43002
rect 26956 42948 27012 42950
rect 27036 42948 27092 42950
rect 27116 42948 27172 42950
rect 27196 42948 27252 42950
rect 31956 43002 32012 43004
rect 32036 43002 32092 43004
rect 32116 43002 32172 43004
rect 32196 43002 32252 43004
rect 31956 42950 32002 43002
rect 32002 42950 32012 43002
rect 32036 42950 32066 43002
rect 32066 42950 32078 43002
rect 32078 42950 32092 43002
rect 32116 42950 32130 43002
rect 32130 42950 32142 43002
rect 32142 42950 32172 43002
rect 32196 42950 32206 43002
rect 32206 42950 32252 43002
rect 31956 42948 32012 42950
rect 32036 42948 32092 42950
rect 32116 42948 32172 42950
rect 32196 42948 32252 42950
rect 36956 43002 37012 43004
rect 37036 43002 37092 43004
rect 37116 43002 37172 43004
rect 37196 43002 37252 43004
rect 36956 42950 37002 43002
rect 37002 42950 37012 43002
rect 37036 42950 37066 43002
rect 37066 42950 37078 43002
rect 37078 42950 37092 43002
rect 37116 42950 37130 43002
rect 37130 42950 37142 43002
rect 37142 42950 37172 43002
rect 37196 42950 37206 43002
rect 37206 42950 37252 43002
rect 36956 42948 37012 42950
rect 37036 42948 37092 42950
rect 37116 42948 37172 42950
rect 37196 42948 37252 42950
rect 41956 43002 42012 43004
rect 42036 43002 42092 43004
rect 42116 43002 42172 43004
rect 42196 43002 42252 43004
rect 41956 42950 42002 43002
rect 42002 42950 42012 43002
rect 42036 42950 42066 43002
rect 42066 42950 42078 43002
rect 42078 42950 42092 43002
rect 42116 42950 42130 43002
rect 42130 42950 42142 43002
rect 42142 42950 42172 43002
rect 42196 42950 42206 43002
rect 42206 42950 42252 43002
rect 41956 42948 42012 42950
rect 42036 42948 42092 42950
rect 42116 42948 42172 42950
rect 42196 42948 42252 42950
rect 46956 43002 47012 43004
rect 47036 43002 47092 43004
rect 47116 43002 47172 43004
rect 47196 43002 47252 43004
rect 46956 42950 47002 43002
rect 47002 42950 47012 43002
rect 47036 42950 47066 43002
rect 47066 42950 47078 43002
rect 47078 42950 47092 43002
rect 47116 42950 47130 43002
rect 47130 42950 47142 43002
rect 47142 42950 47172 43002
rect 47196 42950 47206 43002
rect 47206 42950 47252 43002
rect 46956 42948 47012 42950
rect 47036 42948 47092 42950
rect 47116 42948 47172 42950
rect 47196 42948 47252 42950
rect 51956 43002 52012 43004
rect 52036 43002 52092 43004
rect 52116 43002 52172 43004
rect 52196 43002 52252 43004
rect 51956 42950 52002 43002
rect 52002 42950 52012 43002
rect 52036 42950 52066 43002
rect 52066 42950 52078 43002
rect 52078 42950 52092 43002
rect 52116 42950 52130 43002
rect 52130 42950 52142 43002
rect 52142 42950 52172 43002
rect 52196 42950 52206 43002
rect 52206 42950 52252 43002
rect 51956 42948 52012 42950
rect 52036 42948 52092 42950
rect 52116 42948 52172 42950
rect 52196 42948 52252 42950
rect 56956 43002 57012 43004
rect 57036 43002 57092 43004
rect 57116 43002 57172 43004
rect 57196 43002 57252 43004
rect 56956 42950 57002 43002
rect 57002 42950 57012 43002
rect 57036 42950 57066 43002
rect 57066 42950 57078 43002
rect 57078 42950 57092 43002
rect 57116 42950 57130 43002
rect 57130 42950 57142 43002
rect 57142 42950 57172 43002
rect 57196 42950 57206 43002
rect 57206 42950 57252 43002
rect 56956 42948 57012 42950
rect 57036 42948 57092 42950
rect 57116 42948 57172 42950
rect 57196 42948 57252 42950
rect 58530 42472 58586 42528
rect 2616 42458 2672 42460
rect 2696 42458 2752 42460
rect 2776 42458 2832 42460
rect 2856 42458 2912 42460
rect 2616 42406 2662 42458
rect 2662 42406 2672 42458
rect 2696 42406 2726 42458
rect 2726 42406 2738 42458
rect 2738 42406 2752 42458
rect 2776 42406 2790 42458
rect 2790 42406 2802 42458
rect 2802 42406 2832 42458
rect 2856 42406 2866 42458
rect 2866 42406 2912 42458
rect 2616 42404 2672 42406
rect 2696 42404 2752 42406
rect 2776 42404 2832 42406
rect 2856 42404 2912 42406
rect 7616 42458 7672 42460
rect 7696 42458 7752 42460
rect 7776 42458 7832 42460
rect 7856 42458 7912 42460
rect 7616 42406 7662 42458
rect 7662 42406 7672 42458
rect 7696 42406 7726 42458
rect 7726 42406 7738 42458
rect 7738 42406 7752 42458
rect 7776 42406 7790 42458
rect 7790 42406 7802 42458
rect 7802 42406 7832 42458
rect 7856 42406 7866 42458
rect 7866 42406 7912 42458
rect 7616 42404 7672 42406
rect 7696 42404 7752 42406
rect 7776 42404 7832 42406
rect 7856 42404 7912 42406
rect 12616 42458 12672 42460
rect 12696 42458 12752 42460
rect 12776 42458 12832 42460
rect 12856 42458 12912 42460
rect 12616 42406 12662 42458
rect 12662 42406 12672 42458
rect 12696 42406 12726 42458
rect 12726 42406 12738 42458
rect 12738 42406 12752 42458
rect 12776 42406 12790 42458
rect 12790 42406 12802 42458
rect 12802 42406 12832 42458
rect 12856 42406 12866 42458
rect 12866 42406 12912 42458
rect 12616 42404 12672 42406
rect 12696 42404 12752 42406
rect 12776 42404 12832 42406
rect 12856 42404 12912 42406
rect 17616 42458 17672 42460
rect 17696 42458 17752 42460
rect 17776 42458 17832 42460
rect 17856 42458 17912 42460
rect 17616 42406 17662 42458
rect 17662 42406 17672 42458
rect 17696 42406 17726 42458
rect 17726 42406 17738 42458
rect 17738 42406 17752 42458
rect 17776 42406 17790 42458
rect 17790 42406 17802 42458
rect 17802 42406 17832 42458
rect 17856 42406 17866 42458
rect 17866 42406 17912 42458
rect 17616 42404 17672 42406
rect 17696 42404 17752 42406
rect 17776 42404 17832 42406
rect 17856 42404 17912 42406
rect 22616 42458 22672 42460
rect 22696 42458 22752 42460
rect 22776 42458 22832 42460
rect 22856 42458 22912 42460
rect 22616 42406 22662 42458
rect 22662 42406 22672 42458
rect 22696 42406 22726 42458
rect 22726 42406 22738 42458
rect 22738 42406 22752 42458
rect 22776 42406 22790 42458
rect 22790 42406 22802 42458
rect 22802 42406 22832 42458
rect 22856 42406 22866 42458
rect 22866 42406 22912 42458
rect 22616 42404 22672 42406
rect 22696 42404 22752 42406
rect 22776 42404 22832 42406
rect 22856 42404 22912 42406
rect 27616 42458 27672 42460
rect 27696 42458 27752 42460
rect 27776 42458 27832 42460
rect 27856 42458 27912 42460
rect 27616 42406 27662 42458
rect 27662 42406 27672 42458
rect 27696 42406 27726 42458
rect 27726 42406 27738 42458
rect 27738 42406 27752 42458
rect 27776 42406 27790 42458
rect 27790 42406 27802 42458
rect 27802 42406 27832 42458
rect 27856 42406 27866 42458
rect 27866 42406 27912 42458
rect 27616 42404 27672 42406
rect 27696 42404 27752 42406
rect 27776 42404 27832 42406
rect 27856 42404 27912 42406
rect 32616 42458 32672 42460
rect 32696 42458 32752 42460
rect 32776 42458 32832 42460
rect 32856 42458 32912 42460
rect 32616 42406 32662 42458
rect 32662 42406 32672 42458
rect 32696 42406 32726 42458
rect 32726 42406 32738 42458
rect 32738 42406 32752 42458
rect 32776 42406 32790 42458
rect 32790 42406 32802 42458
rect 32802 42406 32832 42458
rect 32856 42406 32866 42458
rect 32866 42406 32912 42458
rect 32616 42404 32672 42406
rect 32696 42404 32752 42406
rect 32776 42404 32832 42406
rect 32856 42404 32912 42406
rect 37616 42458 37672 42460
rect 37696 42458 37752 42460
rect 37776 42458 37832 42460
rect 37856 42458 37912 42460
rect 37616 42406 37662 42458
rect 37662 42406 37672 42458
rect 37696 42406 37726 42458
rect 37726 42406 37738 42458
rect 37738 42406 37752 42458
rect 37776 42406 37790 42458
rect 37790 42406 37802 42458
rect 37802 42406 37832 42458
rect 37856 42406 37866 42458
rect 37866 42406 37912 42458
rect 37616 42404 37672 42406
rect 37696 42404 37752 42406
rect 37776 42404 37832 42406
rect 37856 42404 37912 42406
rect 42616 42458 42672 42460
rect 42696 42458 42752 42460
rect 42776 42458 42832 42460
rect 42856 42458 42912 42460
rect 42616 42406 42662 42458
rect 42662 42406 42672 42458
rect 42696 42406 42726 42458
rect 42726 42406 42738 42458
rect 42738 42406 42752 42458
rect 42776 42406 42790 42458
rect 42790 42406 42802 42458
rect 42802 42406 42832 42458
rect 42856 42406 42866 42458
rect 42866 42406 42912 42458
rect 42616 42404 42672 42406
rect 42696 42404 42752 42406
rect 42776 42404 42832 42406
rect 42856 42404 42912 42406
rect 47616 42458 47672 42460
rect 47696 42458 47752 42460
rect 47776 42458 47832 42460
rect 47856 42458 47912 42460
rect 47616 42406 47662 42458
rect 47662 42406 47672 42458
rect 47696 42406 47726 42458
rect 47726 42406 47738 42458
rect 47738 42406 47752 42458
rect 47776 42406 47790 42458
rect 47790 42406 47802 42458
rect 47802 42406 47832 42458
rect 47856 42406 47866 42458
rect 47866 42406 47912 42458
rect 47616 42404 47672 42406
rect 47696 42404 47752 42406
rect 47776 42404 47832 42406
rect 47856 42404 47912 42406
rect 52616 42458 52672 42460
rect 52696 42458 52752 42460
rect 52776 42458 52832 42460
rect 52856 42458 52912 42460
rect 52616 42406 52662 42458
rect 52662 42406 52672 42458
rect 52696 42406 52726 42458
rect 52726 42406 52738 42458
rect 52738 42406 52752 42458
rect 52776 42406 52790 42458
rect 52790 42406 52802 42458
rect 52802 42406 52832 42458
rect 52856 42406 52866 42458
rect 52866 42406 52912 42458
rect 52616 42404 52672 42406
rect 52696 42404 52752 42406
rect 52776 42404 52832 42406
rect 52856 42404 52912 42406
rect 57616 42458 57672 42460
rect 57696 42458 57752 42460
rect 57776 42458 57832 42460
rect 57856 42458 57912 42460
rect 57616 42406 57662 42458
rect 57662 42406 57672 42458
rect 57696 42406 57726 42458
rect 57726 42406 57738 42458
rect 57738 42406 57752 42458
rect 57776 42406 57790 42458
rect 57790 42406 57802 42458
rect 57802 42406 57832 42458
rect 57856 42406 57866 42458
rect 57866 42406 57912 42458
rect 57616 42404 57672 42406
rect 57696 42404 57752 42406
rect 57776 42404 57832 42406
rect 57856 42404 57912 42406
rect 1956 41914 2012 41916
rect 2036 41914 2092 41916
rect 2116 41914 2172 41916
rect 2196 41914 2252 41916
rect 1956 41862 2002 41914
rect 2002 41862 2012 41914
rect 2036 41862 2066 41914
rect 2066 41862 2078 41914
rect 2078 41862 2092 41914
rect 2116 41862 2130 41914
rect 2130 41862 2142 41914
rect 2142 41862 2172 41914
rect 2196 41862 2206 41914
rect 2206 41862 2252 41914
rect 1956 41860 2012 41862
rect 2036 41860 2092 41862
rect 2116 41860 2172 41862
rect 2196 41860 2252 41862
rect 6956 41914 7012 41916
rect 7036 41914 7092 41916
rect 7116 41914 7172 41916
rect 7196 41914 7252 41916
rect 6956 41862 7002 41914
rect 7002 41862 7012 41914
rect 7036 41862 7066 41914
rect 7066 41862 7078 41914
rect 7078 41862 7092 41914
rect 7116 41862 7130 41914
rect 7130 41862 7142 41914
rect 7142 41862 7172 41914
rect 7196 41862 7206 41914
rect 7206 41862 7252 41914
rect 6956 41860 7012 41862
rect 7036 41860 7092 41862
rect 7116 41860 7172 41862
rect 7196 41860 7252 41862
rect 11956 41914 12012 41916
rect 12036 41914 12092 41916
rect 12116 41914 12172 41916
rect 12196 41914 12252 41916
rect 11956 41862 12002 41914
rect 12002 41862 12012 41914
rect 12036 41862 12066 41914
rect 12066 41862 12078 41914
rect 12078 41862 12092 41914
rect 12116 41862 12130 41914
rect 12130 41862 12142 41914
rect 12142 41862 12172 41914
rect 12196 41862 12206 41914
rect 12206 41862 12252 41914
rect 11956 41860 12012 41862
rect 12036 41860 12092 41862
rect 12116 41860 12172 41862
rect 12196 41860 12252 41862
rect 16956 41914 17012 41916
rect 17036 41914 17092 41916
rect 17116 41914 17172 41916
rect 17196 41914 17252 41916
rect 16956 41862 17002 41914
rect 17002 41862 17012 41914
rect 17036 41862 17066 41914
rect 17066 41862 17078 41914
rect 17078 41862 17092 41914
rect 17116 41862 17130 41914
rect 17130 41862 17142 41914
rect 17142 41862 17172 41914
rect 17196 41862 17206 41914
rect 17206 41862 17252 41914
rect 16956 41860 17012 41862
rect 17036 41860 17092 41862
rect 17116 41860 17172 41862
rect 17196 41860 17252 41862
rect 21956 41914 22012 41916
rect 22036 41914 22092 41916
rect 22116 41914 22172 41916
rect 22196 41914 22252 41916
rect 21956 41862 22002 41914
rect 22002 41862 22012 41914
rect 22036 41862 22066 41914
rect 22066 41862 22078 41914
rect 22078 41862 22092 41914
rect 22116 41862 22130 41914
rect 22130 41862 22142 41914
rect 22142 41862 22172 41914
rect 22196 41862 22206 41914
rect 22206 41862 22252 41914
rect 21956 41860 22012 41862
rect 22036 41860 22092 41862
rect 22116 41860 22172 41862
rect 22196 41860 22252 41862
rect 26956 41914 27012 41916
rect 27036 41914 27092 41916
rect 27116 41914 27172 41916
rect 27196 41914 27252 41916
rect 26956 41862 27002 41914
rect 27002 41862 27012 41914
rect 27036 41862 27066 41914
rect 27066 41862 27078 41914
rect 27078 41862 27092 41914
rect 27116 41862 27130 41914
rect 27130 41862 27142 41914
rect 27142 41862 27172 41914
rect 27196 41862 27206 41914
rect 27206 41862 27252 41914
rect 26956 41860 27012 41862
rect 27036 41860 27092 41862
rect 27116 41860 27172 41862
rect 27196 41860 27252 41862
rect 31956 41914 32012 41916
rect 32036 41914 32092 41916
rect 32116 41914 32172 41916
rect 32196 41914 32252 41916
rect 31956 41862 32002 41914
rect 32002 41862 32012 41914
rect 32036 41862 32066 41914
rect 32066 41862 32078 41914
rect 32078 41862 32092 41914
rect 32116 41862 32130 41914
rect 32130 41862 32142 41914
rect 32142 41862 32172 41914
rect 32196 41862 32206 41914
rect 32206 41862 32252 41914
rect 31956 41860 32012 41862
rect 32036 41860 32092 41862
rect 32116 41860 32172 41862
rect 32196 41860 32252 41862
rect 36956 41914 37012 41916
rect 37036 41914 37092 41916
rect 37116 41914 37172 41916
rect 37196 41914 37252 41916
rect 36956 41862 37002 41914
rect 37002 41862 37012 41914
rect 37036 41862 37066 41914
rect 37066 41862 37078 41914
rect 37078 41862 37092 41914
rect 37116 41862 37130 41914
rect 37130 41862 37142 41914
rect 37142 41862 37172 41914
rect 37196 41862 37206 41914
rect 37206 41862 37252 41914
rect 36956 41860 37012 41862
rect 37036 41860 37092 41862
rect 37116 41860 37172 41862
rect 37196 41860 37252 41862
rect 41956 41914 42012 41916
rect 42036 41914 42092 41916
rect 42116 41914 42172 41916
rect 42196 41914 42252 41916
rect 41956 41862 42002 41914
rect 42002 41862 42012 41914
rect 42036 41862 42066 41914
rect 42066 41862 42078 41914
rect 42078 41862 42092 41914
rect 42116 41862 42130 41914
rect 42130 41862 42142 41914
rect 42142 41862 42172 41914
rect 42196 41862 42206 41914
rect 42206 41862 42252 41914
rect 41956 41860 42012 41862
rect 42036 41860 42092 41862
rect 42116 41860 42172 41862
rect 42196 41860 42252 41862
rect 46956 41914 47012 41916
rect 47036 41914 47092 41916
rect 47116 41914 47172 41916
rect 47196 41914 47252 41916
rect 46956 41862 47002 41914
rect 47002 41862 47012 41914
rect 47036 41862 47066 41914
rect 47066 41862 47078 41914
rect 47078 41862 47092 41914
rect 47116 41862 47130 41914
rect 47130 41862 47142 41914
rect 47142 41862 47172 41914
rect 47196 41862 47206 41914
rect 47206 41862 47252 41914
rect 46956 41860 47012 41862
rect 47036 41860 47092 41862
rect 47116 41860 47172 41862
rect 47196 41860 47252 41862
rect 51956 41914 52012 41916
rect 52036 41914 52092 41916
rect 52116 41914 52172 41916
rect 52196 41914 52252 41916
rect 51956 41862 52002 41914
rect 52002 41862 52012 41914
rect 52036 41862 52066 41914
rect 52066 41862 52078 41914
rect 52078 41862 52092 41914
rect 52116 41862 52130 41914
rect 52130 41862 52142 41914
rect 52142 41862 52172 41914
rect 52196 41862 52206 41914
rect 52206 41862 52252 41914
rect 51956 41860 52012 41862
rect 52036 41860 52092 41862
rect 52116 41860 52172 41862
rect 52196 41860 52252 41862
rect 56956 41914 57012 41916
rect 57036 41914 57092 41916
rect 57116 41914 57172 41916
rect 57196 41914 57252 41916
rect 56956 41862 57002 41914
rect 57002 41862 57012 41914
rect 57036 41862 57066 41914
rect 57066 41862 57078 41914
rect 57078 41862 57092 41914
rect 57116 41862 57130 41914
rect 57130 41862 57142 41914
rect 57142 41862 57172 41914
rect 57196 41862 57206 41914
rect 57206 41862 57252 41914
rect 56956 41860 57012 41862
rect 57036 41860 57092 41862
rect 57116 41860 57172 41862
rect 57196 41860 57252 41862
rect 58530 41656 58586 41712
rect 2616 41370 2672 41372
rect 2696 41370 2752 41372
rect 2776 41370 2832 41372
rect 2856 41370 2912 41372
rect 2616 41318 2662 41370
rect 2662 41318 2672 41370
rect 2696 41318 2726 41370
rect 2726 41318 2738 41370
rect 2738 41318 2752 41370
rect 2776 41318 2790 41370
rect 2790 41318 2802 41370
rect 2802 41318 2832 41370
rect 2856 41318 2866 41370
rect 2866 41318 2912 41370
rect 2616 41316 2672 41318
rect 2696 41316 2752 41318
rect 2776 41316 2832 41318
rect 2856 41316 2912 41318
rect 7616 41370 7672 41372
rect 7696 41370 7752 41372
rect 7776 41370 7832 41372
rect 7856 41370 7912 41372
rect 7616 41318 7662 41370
rect 7662 41318 7672 41370
rect 7696 41318 7726 41370
rect 7726 41318 7738 41370
rect 7738 41318 7752 41370
rect 7776 41318 7790 41370
rect 7790 41318 7802 41370
rect 7802 41318 7832 41370
rect 7856 41318 7866 41370
rect 7866 41318 7912 41370
rect 7616 41316 7672 41318
rect 7696 41316 7752 41318
rect 7776 41316 7832 41318
rect 7856 41316 7912 41318
rect 12616 41370 12672 41372
rect 12696 41370 12752 41372
rect 12776 41370 12832 41372
rect 12856 41370 12912 41372
rect 12616 41318 12662 41370
rect 12662 41318 12672 41370
rect 12696 41318 12726 41370
rect 12726 41318 12738 41370
rect 12738 41318 12752 41370
rect 12776 41318 12790 41370
rect 12790 41318 12802 41370
rect 12802 41318 12832 41370
rect 12856 41318 12866 41370
rect 12866 41318 12912 41370
rect 12616 41316 12672 41318
rect 12696 41316 12752 41318
rect 12776 41316 12832 41318
rect 12856 41316 12912 41318
rect 17616 41370 17672 41372
rect 17696 41370 17752 41372
rect 17776 41370 17832 41372
rect 17856 41370 17912 41372
rect 17616 41318 17662 41370
rect 17662 41318 17672 41370
rect 17696 41318 17726 41370
rect 17726 41318 17738 41370
rect 17738 41318 17752 41370
rect 17776 41318 17790 41370
rect 17790 41318 17802 41370
rect 17802 41318 17832 41370
rect 17856 41318 17866 41370
rect 17866 41318 17912 41370
rect 17616 41316 17672 41318
rect 17696 41316 17752 41318
rect 17776 41316 17832 41318
rect 17856 41316 17912 41318
rect 22616 41370 22672 41372
rect 22696 41370 22752 41372
rect 22776 41370 22832 41372
rect 22856 41370 22912 41372
rect 22616 41318 22662 41370
rect 22662 41318 22672 41370
rect 22696 41318 22726 41370
rect 22726 41318 22738 41370
rect 22738 41318 22752 41370
rect 22776 41318 22790 41370
rect 22790 41318 22802 41370
rect 22802 41318 22832 41370
rect 22856 41318 22866 41370
rect 22866 41318 22912 41370
rect 22616 41316 22672 41318
rect 22696 41316 22752 41318
rect 22776 41316 22832 41318
rect 22856 41316 22912 41318
rect 27616 41370 27672 41372
rect 27696 41370 27752 41372
rect 27776 41370 27832 41372
rect 27856 41370 27912 41372
rect 27616 41318 27662 41370
rect 27662 41318 27672 41370
rect 27696 41318 27726 41370
rect 27726 41318 27738 41370
rect 27738 41318 27752 41370
rect 27776 41318 27790 41370
rect 27790 41318 27802 41370
rect 27802 41318 27832 41370
rect 27856 41318 27866 41370
rect 27866 41318 27912 41370
rect 27616 41316 27672 41318
rect 27696 41316 27752 41318
rect 27776 41316 27832 41318
rect 27856 41316 27912 41318
rect 32616 41370 32672 41372
rect 32696 41370 32752 41372
rect 32776 41370 32832 41372
rect 32856 41370 32912 41372
rect 32616 41318 32662 41370
rect 32662 41318 32672 41370
rect 32696 41318 32726 41370
rect 32726 41318 32738 41370
rect 32738 41318 32752 41370
rect 32776 41318 32790 41370
rect 32790 41318 32802 41370
rect 32802 41318 32832 41370
rect 32856 41318 32866 41370
rect 32866 41318 32912 41370
rect 32616 41316 32672 41318
rect 32696 41316 32752 41318
rect 32776 41316 32832 41318
rect 32856 41316 32912 41318
rect 37616 41370 37672 41372
rect 37696 41370 37752 41372
rect 37776 41370 37832 41372
rect 37856 41370 37912 41372
rect 37616 41318 37662 41370
rect 37662 41318 37672 41370
rect 37696 41318 37726 41370
rect 37726 41318 37738 41370
rect 37738 41318 37752 41370
rect 37776 41318 37790 41370
rect 37790 41318 37802 41370
rect 37802 41318 37832 41370
rect 37856 41318 37866 41370
rect 37866 41318 37912 41370
rect 37616 41316 37672 41318
rect 37696 41316 37752 41318
rect 37776 41316 37832 41318
rect 37856 41316 37912 41318
rect 42616 41370 42672 41372
rect 42696 41370 42752 41372
rect 42776 41370 42832 41372
rect 42856 41370 42912 41372
rect 42616 41318 42662 41370
rect 42662 41318 42672 41370
rect 42696 41318 42726 41370
rect 42726 41318 42738 41370
rect 42738 41318 42752 41370
rect 42776 41318 42790 41370
rect 42790 41318 42802 41370
rect 42802 41318 42832 41370
rect 42856 41318 42866 41370
rect 42866 41318 42912 41370
rect 42616 41316 42672 41318
rect 42696 41316 42752 41318
rect 42776 41316 42832 41318
rect 42856 41316 42912 41318
rect 47616 41370 47672 41372
rect 47696 41370 47752 41372
rect 47776 41370 47832 41372
rect 47856 41370 47912 41372
rect 47616 41318 47662 41370
rect 47662 41318 47672 41370
rect 47696 41318 47726 41370
rect 47726 41318 47738 41370
rect 47738 41318 47752 41370
rect 47776 41318 47790 41370
rect 47790 41318 47802 41370
rect 47802 41318 47832 41370
rect 47856 41318 47866 41370
rect 47866 41318 47912 41370
rect 47616 41316 47672 41318
rect 47696 41316 47752 41318
rect 47776 41316 47832 41318
rect 47856 41316 47912 41318
rect 52616 41370 52672 41372
rect 52696 41370 52752 41372
rect 52776 41370 52832 41372
rect 52856 41370 52912 41372
rect 52616 41318 52662 41370
rect 52662 41318 52672 41370
rect 52696 41318 52726 41370
rect 52726 41318 52738 41370
rect 52738 41318 52752 41370
rect 52776 41318 52790 41370
rect 52790 41318 52802 41370
rect 52802 41318 52832 41370
rect 52856 41318 52866 41370
rect 52866 41318 52912 41370
rect 52616 41316 52672 41318
rect 52696 41316 52752 41318
rect 52776 41316 52832 41318
rect 52856 41316 52912 41318
rect 57616 41370 57672 41372
rect 57696 41370 57752 41372
rect 57776 41370 57832 41372
rect 57856 41370 57912 41372
rect 57616 41318 57662 41370
rect 57662 41318 57672 41370
rect 57696 41318 57726 41370
rect 57726 41318 57738 41370
rect 57738 41318 57752 41370
rect 57776 41318 57790 41370
rect 57790 41318 57802 41370
rect 57802 41318 57832 41370
rect 57856 41318 57866 41370
rect 57866 41318 57912 41370
rect 57616 41316 57672 41318
rect 57696 41316 57752 41318
rect 57776 41316 57832 41318
rect 57856 41316 57912 41318
rect 58530 40876 58532 40896
rect 58532 40876 58584 40896
rect 58584 40876 58586 40896
rect 58530 40840 58586 40876
rect 1956 40826 2012 40828
rect 2036 40826 2092 40828
rect 2116 40826 2172 40828
rect 2196 40826 2252 40828
rect 1956 40774 2002 40826
rect 2002 40774 2012 40826
rect 2036 40774 2066 40826
rect 2066 40774 2078 40826
rect 2078 40774 2092 40826
rect 2116 40774 2130 40826
rect 2130 40774 2142 40826
rect 2142 40774 2172 40826
rect 2196 40774 2206 40826
rect 2206 40774 2252 40826
rect 1956 40772 2012 40774
rect 2036 40772 2092 40774
rect 2116 40772 2172 40774
rect 2196 40772 2252 40774
rect 6956 40826 7012 40828
rect 7036 40826 7092 40828
rect 7116 40826 7172 40828
rect 7196 40826 7252 40828
rect 6956 40774 7002 40826
rect 7002 40774 7012 40826
rect 7036 40774 7066 40826
rect 7066 40774 7078 40826
rect 7078 40774 7092 40826
rect 7116 40774 7130 40826
rect 7130 40774 7142 40826
rect 7142 40774 7172 40826
rect 7196 40774 7206 40826
rect 7206 40774 7252 40826
rect 6956 40772 7012 40774
rect 7036 40772 7092 40774
rect 7116 40772 7172 40774
rect 7196 40772 7252 40774
rect 11956 40826 12012 40828
rect 12036 40826 12092 40828
rect 12116 40826 12172 40828
rect 12196 40826 12252 40828
rect 11956 40774 12002 40826
rect 12002 40774 12012 40826
rect 12036 40774 12066 40826
rect 12066 40774 12078 40826
rect 12078 40774 12092 40826
rect 12116 40774 12130 40826
rect 12130 40774 12142 40826
rect 12142 40774 12172 40826
rect 12196 40774 12206 40826
rect 12206 40774 12252 40826
rect 11956 40772 12012 40774
rect 12036 40772 12092 40774
rect 12116 40772 12172 40774
rect 12196 40772 12252 40774
rect 16956 40826 17012 40828
rect 17036 40826 17092 40828
rect 17116 40826 17172 40828
rect 17196 40826 17252 40828
rect 16956 40774 17002 40826
rect 17002 40774 17012 40826
rect 17036 40774 17066 40826
rect 17066 40774 17078 40826
rect 17078 40774 17092 40826
rect 17116 40774 17130 40826
rect 17130 40774 17142 40826
rect 17142 40774 17172 40826
rect 17196 40774 17206 40826
rect 17206 40774 17252 40826
rect 16956 40772 17012 40774
rect 17036 40772 17092 40774
rect 17116 40772 17172 40774
rect 17196 40772 17252 40774
rect 21956 40826 22012 40828
rect 22036 40826 22092 40828
rect 22116 40826 22172 40828
rect 22196 40826 22252 40828
rect 21956 40774 22002 40826
rect 22002 40774 22012 40826
rect 22036 40774 22066 40826
rect 22066 40774 22078 40826
rect 22078 40774 22092 40826
rect 22116 40774 22130 40826
rect 22130 40774 22142 40826
rect 22142 40774 22172 40826
rect 22196 40774 22206 40826
rect 22206 40774 22252 40826
rect 21956 40772 22012 40774
rect 22036 40772 22092 40774
rect 22116 40772 22172 40774
rect 22196 40772 22252 40774
rect 26956 40826 27012 40828
rect 27036 40826 27092 40828
rect 27116 40826 27172 40828
rect 27196 40826 27252 40828
rect 26956 40774 27002 40826
rect 27002 40774 27012 40826
rect 27036 40774 27066 40826
rect 27066 40774 27078 40826
rect 27078 40774 27092 40826
rect 27116 40774 27130 40826
rect 27130 40774 27142 40826
rect 27142 40774 27172 40826
rect 27196 40774 27206 40826
rect 27206 40774 27252 40826
rect 26956 40772 27012 40774
rect 27036 40772 27092 40774
rect 27116 40772 27172 40774
rect 27196 40772 27252 40774
rect 31956 40826 32012 40828
rect 32036 40826 32092 40828
rect 32116 40826 32172 40828
rect 32196 40826 32252 40828
rect 31956 40774 32002 40826
rect 32002 40774 32012 40826
rect 32036 40774 32066 40826
rect 32066 40774 32078 40826
rect 32078 40774 32092 40826
rect 32116 40774 32130 40826
rect 32130 40774 32142 40826
rect 32142 40774 32172 40826
rect 32196 40774 32206 40826
rect 32206 40774 32252 40826
rect 31956 40772 32012 40774
rect 32036 40772 32092 40774
rect 32116 40772 32172 40774
rect 32196 40772 32252 40774
rect 36956 40826 37012 40828
rect 37036 40826 37092 40828
rect 37116 40826 37172 40828
rect 37196 40826 37252 40828
rect 36956 40774 37002 40826
rect 37002 40774 37012 40826
rect 37036 40774 37066 40826
rect 37066 40774 37078 40826
rect 37078 40774 37092 40826
rect 37116 40774 37130 40826
rect 37130 40774 37142 40826
rect 37142 40774 37172 40826
rect 37196 40774 37206 40826
rect 37206 40774 37252 40826
rect 36956 40772 37012 40774
rect 37036 40772 37092 40774
rect 37116 40772 37172 40774
rect 37196 40772 37252 40774
rect 41956 40826 42012 40828
rect 42036 40826 42092 40828
rect 42116 40826 42172 40828
rect 42196 40826 42252 40828
rect 41956 40774 42002 40826
rect 42002 40774 42012 40826
rect 42036 40774 42066 40826
rect 42066 40774 42078 40826
rect 42078 40774 42092 40826
rect 42116 40774 42130 40826
rect 42130 40774 42142 40826
rect 42142 40774 42172 40826
rect 42196 40774 42206 40826
rect 42206 40774 42252 40826
rect 41956 40772 42012 40774
rect 42036 40772 42092 40774
rect 42116 40772 42172 40774
rect 42196 40772 42252 40774
rect 46956 40826 47012 40828
rect 47036 40826 47092 40828
rect 47116 40826 47172 40828
rect 47196 40826 47252 40828
rect 46956 40774 47002 40826
rect 47002 40774 47012 40826
rect 47036 40774 47066 40826
rect 47066 40774 47078 40826
rect 47078 40774 47092 40826
rect 47116 40774 47130 40826
rect 47130 40774 47142 40826
rect 47142 40774 47172 40826
rect 47196 40774 47206 40826
rect 47206 40774 47252 40826
rect 46956 40772 47012 40774
rect 47036 40772 47092 40774
rect 47116 40772 47172 40774
rect 47196 40772 47252 40774
rect 51956 40826 52012 40828
rect 52036 40826 52092 40828
rect 52116 40826 52172 40828
rect 52196 40826 52252 40828
rect 51956 40774 52002 40826
rect 52002 40774 52012 40826
rect 52036 40774 52066 40826
rect 52066 40774 52078 40826
rect 52078 40774 52092 40826
rect 52116 40774 52130 40826
rect 52130 40774 52142 40826
rect 52142 40774 52172 40826
rect 52196 40774 52206 40826
rect 52206 40774 52252 40826
rect 51956 40772 52012 40774
rect 52036 40772 52092 40774
rect 52116 40772 52172 40774
rect 52196 40772 52252 40774
rect 56956 40826 57012 40828
rect 57036 40826 57092 40828
rect 57116 40826 57172 40828
rect 57196 40826 57252 40828
rect 56956 40774 57002 40826
rect 57002 40774 57012 40826
rect 57036 40774 57066 40826
rect 57066 40774 57078 40826
rect 57078 40774 57092 40826
rect 57116 40774 57130 40826
rect 57130 40774 57142 40826
rect 57142 40774 57172 40826
rect 57196 40774 57206 40826
rect 57206 40774 57252 40826
rect 56956 40772 57012 40774
rect 57036 40772 57092 40774
rect 57116 40772 57172 40774
rect 57196 40772 57252 40774
rect 2616 40282 2672 40284
rect 2696 40282 2752 40284
rect 2776 40282 2832 40284
rect 2856 40282 2912 40284
rect 2616 40230 2662 40282
rect 2662 40230 2672 40282
rect 2696 40230 2726 40282
rect 2726 40230 2738 40282
rect 2738 40230 2752 40282
rect 2776 40230 2790 40282
rect 2790 40230 2802 40282
rect 2802 40230 2832 40282
rect 2856 40230 2866 40282
rect 2866 40230 2912 40282
rect 2616 40228 2672 40230
rect 2696 40228 2752 40230
rect 2776 40228 2832 40230
rect 2856 40228 2912 40230
rect 7616 40282 7672 40284
rect 7696 40282 7752 40284
rect 7776 40282 7832 40284
rect 7856 40282 7912 40284
rect 7616 40230 7662 40282
rect 7662 40230 7672 40282
rect 7696 40230 7726 40282
rect 7726 40230 7738 40282
rect 7738 40230 7752 40282
rect 7776 40230 7790 40282
rect 7790 40230 7802 40282
rect 7802 40230 7832 40282
rect 7856 40230 7866 40282
rect 7866 40230 7912 40282
rect 7616 40228 7672 40230
rect 7696 40228 7752 40230
rect 7776 40228 7832 40230
rect 7856 40228 7912 40230
rect 12616 40282 12672 40284
rect 12696 40282 12752 40284
rect 12776 40282 12832 40284
rect 12856 40282 12912 40284
rect 12616 40230 12662 40282
rect 12662 40230 12672 40282
rect 12696 40230 12726 40282
rect 12726 40230 12738 40282
rect 12738 40230 12752 40282
rect 12776 40230 12790 40282
rect 12790 40230 12802 40282
rect 12802 40230 12832 40282
rect 12856 40230 12866 40282
rect 12866 40230 12912 40282
rect 12616 40228 12672 40230
rect 12696 40228 12752 40230
rect 12776 40228 12832 40230
rect 12856 40228 12912 40230
rect 17616 40282 17672 40284
rect 17696 40282 17752 40284
rect 17776 40282 17832 40284
rect 17856 40282 17912 40284
rect 17616 40230 17662 40282
rect 17662 40230 17672 40282
rect 17696 40230 17726 40282
rect 17726 40230 17738 40282
rect 17738 40230 17752 40282
rect 17776 40230 17790 40282
rect 17790 40230 17802 40282
rect 17802 40230 17832 40282
rect 17856 40230 17866 40282
rect 17866 40230 17912 40282
rect 17616 40228 17672 40230
rect 17696 40228 17752 40230
rect 17776 40228 17832 40230
rect 17856 40228 17912 40230
rect 22616 40282 22672 40284
rect 22696 40282 22752 40284
rect 22776 40282 22832 40284
rect 22856 40282 22912 40284
rect 22616 40230 22662 40282
rect 22662 40230 22672 40282
rect 22696 40230 22726 40282
rect 22726 40230 22738 40282
rect 22738 40230 22752 40282
rect 22776 40230 22790 40282
rect 22790 40230 22802 40282
rect 22802 40230 22832 40282
rect 22856 40230 22866 40282
rect 22866 40230 22912 40282
rect 22616 40228 22672 40230
rect 22696 40228 22752 40230
rect 22776 40228 22832 40230
rect 22856 40228 22912 40230
rect 27616 40282 27672 40284
rect 27696 40282 27752 40284
rect 27776 40282 27832 40284
rect 27856 40282 27912 40284
rect 27616 40230 27662 40282
rect 27662 40230 27672 40282
rect 27696 40230 27726 40282
rect 27726 40230 27738 40282
rect 27738 40230 27752 40282
rect 27776 40230 27790 40282
rect 27790 40230 27802 40282
rect 27802 40230 27832 40282
rect 27856 40230 27866 40282
rect 27866 40230 27912 40282
rect 27616 40228 27672 40230
rect 27696 40228 27752 40230
rect 27776 40228 27832 40230
rect 27856 40228 27912 40230
rect 32616 40282 32672 40284
rect 32696 40282 32752 40284
rect 32776 40282 32832 40284
rect 32856 40282 32912 40284
rect 32616 40230 32662 40282
rect 32662 40230 32672 40282
rect 32696 40230 32726 40282
rect 32726 40230 32738 40282
rect 32738 40230 32752 40282
rect 32776 40230 32790 40282
rect 32790 40230 32802 40282
rect 32802 40230 32832 40282
rect 32856 40230 32866 40282
rect 32866 40230 32912 40282
rect 32616 40228 32672 40230
rect 32696 40228 32752 40230
rect 32776 40228 32832 40230
rect 32856 40228 32912 40230
rect 37616 40282 37672 40284
rect 37696 40282 37752 40284
rect 37776 40282 37832 40284
rect 37856 40282 37912 40284
rect 37616 40230 37662 40282
rect 37662 40230 37672 40282
rect 37696 40230 37726 40282
rect 37726 40230 37738 40282
rect 37738 40230 37752 40282
rect 37776 40230 37790 40282
rect 37790 40230 37802 40282
rect 37802 40230 37832 40282
rect 37856 40230 37866 40282
rect 37866 40230 37912 40282
rect 37616 40228 37672 40230
rect 37696 40228 37752 40230
rect 37776 40228 37832 40230
rect 37856 40228 37912 40230
rect 42616 40282 42672 40284
rect 42696 40282 42752 40284
rect 42776 40282 42832 40284
rect 42856 40282 42912 40284
rect 42616 40230 42662 40282
rect 42662 40230 42672 40282
rect 42696 40230 42726 40282
rect 42726 40230 42738 40282
rect 42738 40230 42752 40282
rect 42776 40230 42790 40282
rect 42790 40230 42802 40282
rect 42802 40230 42832 40282
rect 42856 40230 42866 40282
rect 42866 40230 42912 40282
rect 42616 40228 42672 40230
rect 42696 40228 42752 40230
rect 42776 40228 42832 40230
rect 42856 40228 42912 40230
rect 47616 40282 47672 40284
rect 47696 40282 47752 40284
rect 47776 40282 47832 40284
rect 47856 40282 47912 40284
rect 47616 40230 47662 40282
rect 47662 40230 47672 40282
rect 47696 40230 47726 40282
rect 47726 40230 47738 40282
rect 47738 40230 47752 40282
rect 47776 40230 47790 40282
rect 47790 40230 47802 40282
rect 47802 40230 47832 40282
rect 47856 40230 47866 40282
rect 47866 40230 47912 40282
rect 47616 40228 47672 40230
rect 47696 40228 47752 40230
rect 47776 40228 47832 40230
rect 47856 40228 47912 40230
rect 52616 40282 52672 40284
rect 52696 40282 52752 40284
rect 52776 40282 52832 40284
rect 52856 40282 52912 40284
rect 52616 40230 52662 40282
rect 52662 40230 52672 40282
rect 52696 40230 52726 40282
rect 52726 40230 52738 40282
rect 52738 40230 52752 40282
rect 52776 40230 52790 40282
rect 52790 40230 52802 40282
rect 52802 40230 52832 40282
rect 52856 40230 52866 40282
rect 52866 40230 52912 40282
rect 52616 40228 52672 40230
rect 52696 40228 52752 40230
rect 52776 40228 52832 40230
rect 52856 40228 52912 40230
rect 57616 40282 57672 40284
rect 57696 40282 57752 40284
rect 57776 40282 57832 40284
rect 57856 40282 57912 40284
rect 57616 40230 57662 40282
rect 57662 40230 57672 40282
rect 57696 40230 57726 40282
rect 57726 40230 57738 40282
rect 57738 40230 57752 40282
rect 57776 40230 57790 40282
rect 57790 40230 57802 40282
rect 57802 40230 57832 40282
rect 57856 40230 57866 40282
rect 57866 40230 57912 40282
rect 57616 40228 57672 40230
rect 57696 40228 57752 40230
rect 57776 40228 57832 40230
rect 57856 40228 57912 40230
rect 58530 40024 58586 40080
rect 1956 39738 2012 39740
rect 2036 39738 2092 39740
rect 2116 39738 2172 39740
rect 2196 39738 2252 39740
rect 1956 39686 2002 39738
rect 2002 39686 2012 39738
rect 2036 39686 2066 39738
rect 2066 39686 2078 39738
rect 2078 39686 2092 39738
rect 2116 39686 2130 39738
rect 2130 39686 2142 39738
rect 2142 39686 2172 39738
rect 2196 39686 2206 39738
rect 2206 39686 2252 39738
rect 1956 39684 2012 39686
rect 2036 39684 2092 39686
rect 2116 39684 2172 39686
rect 2196 39684 2252 39686
rect 6956 39738 7012 39740
rect 7036 39738 7092 39740
rect 7116 39738 7172 39740
rect 7196 39738 7252 39740
rect 6956 39686 7002 39738
rect 7002 39686 7012 39738
rect 7036 39686 7066 39738
rect 7066 39686 7078 39738
rect 7078 39686 7092 39738
rect 7116 39686 7130 39738
rect 7130 39686 7142 39738
rect 7142 39686 7172 39738
rect 7196 39686 7206 39738
rect 7206 39686 7252 39738
rect 6956 39684 7012 39686
rect 7036 39684 7092 39686
rect 7116 39684 7172 39686
rect 7196 39684 7252 39686
rect 11956 39738 12012 39740
rect 12036 39738 12092 39740
rect 12116 39738 12172 39740
rect 12196 39738 12252 39740
rect 11956 39686 12002 39738
rect 12002 39686 12012 39738
rect 12036 39686 12066 39738
rect 12066 39686 12078 39738
rect 12078 39686 12092 39738
rect 12116 39686 12130 39738
rect 12130 39686 12142 39738
rect 12142 39686 12172 39738
rect 12196 39686 12206 39738
rect 12206 39686 12252 39738
rect 11956 39684 12012 39686
rect 12036 39684 12092 39686
rect 12116 39684 12172 39686
rect 12196 39684 12252 39686
rect 16956 39738 17012 39740
rect 17036 39738 17092 39740
rect 17116 39738 17172 39740
rect 17196 39738 17252 39740
rect 16956 39686 17002 39738
rect 17002 39686 17012 39738
rect 17036 39686 17066 39738
rect 17066 39686 17078 39738
rect 17078 39686 17092 39738
rect 17116 39686 17130 39738
rect 17130 39686 17142 39738
rect 17142 39686 17172 39738
rect 17196 39686 17206 39738
rect 17206 39686 17252 39738
rect 16956 39684 17012 39686
rect 17036 39684 17092 39686
rect 17116 39684 17172 39686
rect 17196 39684 17252 39686
rect 21956 39738 22012 39740
rect 22036 39738 22092 39740
rect 22116 39738 22172 39740
rect 22196 39738 22252 39740
rect 21956 39686 22002 39738
rect 22002 39686 22012 39738
rect 22036 39686 22066 39738
rect 22066 39686 22078 39738
rect 22078 39686 22092 39738
rect 22116 39686 22130 39738
rect 22130 39686 22142 39738
rect 22142 39686 22172 39738
rect 22196 39686 22206 39738
rect 22206 39686 22252 39738
rect 21956 39684 22012 39686
rect 22036 39684 22092 39686
rect 22116 39684 22172 39686
rect 22196 39684 22252 39686
rect 26956 39738 27012 39740
rect 27036 39738 27092 39740
rect 27116 39738 27172 39740
rect 27196 39738 27252 39740
rect 26956 39686 27002 39738
rect 27002 39686 27012 39738
rect 27036 39686 27066 39738
rect 27066 39686 27078 39738
rect 27078 39686 27092 39738
rect 27116 39686 27130 39738
rect 27130 39686 27142 39738
rect 27142 39686 27172 39738
rect 27196 39686 27206 39738
rect 27206 39686 27252 39738
rect 26956 39684 27012 39686
rect 27036 39684 27092 39686
rect 27116 39684 27172 39686
rect 27196 39684 27252 39686
rect 31956 39738 32012 39740
rect 32036 39738 32092 39740
rect 32116 39738 32172 39740
rect 32196 39738 32252 39740
rect 31956 39686 32002 39738
rect 32002 39686 32012 39738
rect 32036 39686 32066 39738
rect 32066 39686 32078 39738
rect 32078 39686 32092 39738
rect 32116 39686 32130 39738
rect 32130 39686 32142 39738
rect 32142 39686 32172 39738
rect 32196 39686 32206 39738
rect 32206 39686 32252 39738
rect 31956 39684 32012 39686
rect 32036 39684 32092 39686
rect 32116 39684 32172 39686
rect 32196 39684 32252 39686
rect 36956 39738 37012 39740
rect 37036 39738 37092 39740
rect 37116 39738 37172 39740
rect 37196 39738 37252 39740
rect 36956 39686 37002 39738
rect 37002 39686 37012 39738
rect 37036 39686 37066 39738
rect 37066 39686 37078 39738
rect 37078 39686 37092 39738
rect 37116 39686 37130 39738
rect 37130 39686 37142 39738
rect 37142 39686 37172 39738
rect 37196 39686 37206 39738
rect 37206 39686 37252 39738
rect 36956 39684 37012 39686
rect 37036 39684 37092 39686
rect 37116 39684 37172 39686
rect 37196 39684 37252 39686
rect 41956 39738 42012 39740
rect 42036 39738 42092 39740
rect 42116 39738 42172 39740
rect 42196 39738 42252 39740
rect 41956 39686 42002 39738
rect 42002 39686 42012 39738
rect 42036 39686 42066 39738
rect 42066 39686 42078 39738
rect 42078 39686 42092 39738
rect 42116 39686 42130 39738
rect 42130 39686 42142 39738
rect 42142 39686 42172 39738
rect 42196 39686 42206 39738
rect 42206 39686 42252 39738
rect 41956 39684 42012 39686
rect 42036 39684 42092 39686
rect 42116 39684 42172 39686
rect 42196 39684 42252 39686
rect 46956 39738 47012 39740
rect 47036 39738 47092 39740
rect 47116 39738 47172 39740
rect 47196 39738 47252 39740
rect 46956 39686 47002 39738
rect 47002 39686 47012 39738
rect 47036 39686 47066 39738
rect 47066 39686 47078 39738
rect 47078 39686 47092 39738
rect 47116 39686 47130 39738
rect 47130 39686 47142 39738
rect 47142 39686 47172 39738
rect 47196 39686 47206 39738
rect 47206 39686 47252 39738
rect 46956 39684 47012 39686
rect 47036 39684 47092 39686
rect 47116 39684 47172 39686
rect 47196 39684 47252 39686
rect 51956 39738 52012 39740
rect 52036 39738 52092 39740
rect 52116 39738 52172 39740
rect 52196 39738 52252 39740
rect 51956 39686 52002 39738
rect 52002 39686 52012 39738
rect 52036 39686 52066 39738
rect 52066 39686 52078 39738
rect 52078 39686 52092 39738
rect 52116 39686 52130 39738
rect 52130 39686 52142 39738
rect 52142 39686 52172 39738
rect 52196 39686 52206 39738
rect 52206 39686 52252 39738
rect 51956 39684 52012 39686
rect 52036 39684 52092 39686
rect 52116 39684 52172 39686
rect 52196 39684 52252 39686
rect 56956 39738 57012 39740
rect 57036 39738 57092 39740
rect 57116 39738 57172 39740
rect 57196 39738 57252 39740
rect 56956 39686 57002 39738
rect 57002 39686 57012 39738
rect 57036 39686 57066 39738
rect 57066 39686 57078 39738
rect 57078 39686 57092 39738
rect 57116 39686 57130 39738
rect 57130 39686 57142 39738
rect 57142 39686 57172 39738
rect 57196 39686 57206 39738
rect 57206 39686 57252 39738
rect 56956 39684 57012 39686
rect 57036 39684 57092 39686
rect 57116 39684 57172 39686
rect 57196 39684 57252 39686
rect 58530 39208 58586 39264
rect 2616 39194 2672 39196
rect 2696 39194 2752 39196
rect 2776 39194 2832 39196
rect 2856 39194 2912 39196
rect 2616 39142 2662 39194
rect 2662 39142 2672 39194
rect 2696 39142 2726 39194
rect 2726 39142 2738 39194
rect 2738 39142 2752 39194
rect 2776 39142 2790 39194
rect 2790 39142 2802 39194
rect 2802 39142 2832 39194
rect 2856 39142 2866 39194
rect 2866 39142 2912 39194
rect 2616 39140 2672 39142
rect 2696 39140 2752 39142
rect 2776 39140 2832 39142
rect 2856 39140 2912 39142
rect 7616 39194 7672 39196
rect 7696 39194 7752 39196
rect 7776 39194 7832 39196
rect 7856 39194 7912 39196
rect 7616 39142 7662 39194
rect 7662 39142 7672 39194
rect 7696 39142 7726 39194
rect 7726 39142 7738 39194
rect 7738 39142 7752 39194
rect 7776 39142 7790 39194
rect 7790 39142 7802 39194
rect 7802 39142 7832 39194
rect 7856 39142 7866 39194
rect 7866 39142 7912 39194
rect 7616 39140 7672 39142
rect 7696 39140 7752 39142
rect 7776 39140 7832 39142
rect 7856 39140 7912 39142
rect 12616 39194 12672 39196
rect 12696 39194 12752 39196
rect 12776 39194 12832 39196
rect 12856 39194 12912 39196
rect 12616 39142 12662 39194
rect 12662 39142 12672 39194
rect 12696 39142 12726 39194
rect 12726 39142 12738 39194
rect 12738 39142 12752 39194
rect 12776 39142 12790 39194
rect 12790 39142 12802 39194
rect 12802 39142 12832 39194
rect 12856 39142 12866 39194
rect 12866 39142 12912 39194
rect 12616 39140 12672 39142
rect 12696 39140 12752 39142
rect 12776 39140 12832 39142
rect 12856 39140 12912 39142
rect 17616 39194 17672 39196
rect 17696 39194 17752 39196
rect 17776 39194 17832 39196
rect 17856 39194 17912 39196
rect 17616 39142 17662 39194
rect 17662 39142 17672 39194
rect 17696 39142 17726 39194
rect 17726 39142 17738 39194
rect 17738 39142 17752 39194
rect 17776 39142 17790 39194
rect 17790 39142 17802 39194
rect 17802 39142 17832 39194
rect 17856 39142 17866 39194
rect 17866 39142 17912 39194
rect 17616 39140 17672 39142
rect 17696 39140 17752 39142
rect 17776 39140 17832 39142
rect 17856 39140 17912 39142
rect 22616 39194 22672 39196
rect 22696 39194 22752 39196
rect 22776 39194 22832 39196
rect 22856 39194 22912 39196
rect 22616 39142 22662 39194
rect 22662 39142 22672 39194
rect 22696 39142 22726 39194
rect 22726 39142 22738 39194
rect 22738 39142 22752 39194
rect 22776 39142 22790 39194
rect 22790 39142 22802 39194
rect 22802 39142 22832 39194
rect 22856 39142 22866 39194
rect 22866 39142 22912 39194
rect 22616 39140 22672 39142
rect 22696 39140 22752 39142
rect 22776 39140 22832 39142
rect 22856 39140 22912 39142
rect 27616 39194 27672 39196
rect 27696 39194 27752 39196
rect 27776 39194 27832 39196
rect 27856 39194 27912 39196
rect 27616 39142 27662 39194
rect 27662 39142 27672 39194
rect 27696 39142 27726 39194
rect 27726 39142 27738 39194
rect 27738 39142 27752 39194
rect 27776 39142 27790 39194
rect 27790 39142 27802 39194
rect 27802 39142 27832 39194
rect 27856 39142 27866 39194
rect 27866 39142 27912 39194
rect 27616 39140 27672 39142
rect 27696 39140 27752 39142
rect 27776 39140 27832 39142
rect 27856 39140 27912 39142
rect 32616 39194 32672 39196
rect 32696 39194 32752 39196
rect 32776 39194 32832 39196
rect 32856 39194 32912 39196
rect 32616 39142 32662 39194
rect 32662 39142 32672 39194
rect 32696 39142 32726 39194
rect 32726 39142 32738 39194
rect 32738 39142 32752 39194
rect 32776 39142 32790 39194
rect 32790 39142 32802 39194
rect 32802 39142 32832 39194
rect 32856 39142 32866 39194
rect 32866 39142 32912 39194
rect 32616 39140 32672 39142
rect 32696 39140 32752 39142
rect 32776 39140 32832 39142
rect 32856 39140 32912 39142
rect 37616 39194 37672 39196
rect 37696 39194 37752 39196
rect 37776 39194 37832 39196
rect 37856 39194 37912 39196
rect 37616 39142 37662 39194
rect 37662 39142 37672 39194
rect 37696 39142 37726 39194
rect 37726 39142 37738 39194
rect 37738 39142 37752 39194
rect 37776 39142 37790 39194
rect 37790 39142 37802 39194
rect 37802 39142 37832 39194
rect 37856 39142 37866 39194
rect 37866 39142 37912 39194
rect 37616 39140 37672 39142
rect 37696 39140 37752 39142
rect 37776 39140 37832 39142
rect 37856 39140 37912 39142
rect 42616 39194 42672 39196
rect 42696 39194 42752 39196
rect 42776 39194 42832 39196
rect 42856 39194 42912 39196
rect 42616 39142 42662 39194
rect 42662 39142 42672 39194
rect 42696 39142 42726 39194
rect 42726 39142 42738 39194
rect 42738 39142 42752 39194
rect 42776 39142 42790 39194
rect 42790 39142 42802 39194
rect 42802 39142 42832 39194
rect 42856 39142 42866 39194
rect 42866 39142 42912 39194
rect 42616 39140 42672 39142
rect 42696 39140 42752 39142
rect 42776 39140 42832 39142
rect 42856 39140 42912 39142
rect 47616 39194 47672 39196
rect 47696 39194 47752 39196
rect 47776 39194 47832 39196
rect 47856 39194 47912 39196
rect 47616 39142 47662 39194
rect 47662 39142 47672 39194
rect 47696 39142 47726 39194
rect 47726 39142 47738 39194
rect 47738 39142 47752 39194
rect 47776 39142 47790 39194
rect 47790 39142 47802 39194
rect 47802 39142 47832 39194
rect 47856 39142 47866 39194
rect 47866 39142 47912 39194
rect 47616 39140 47672 39142
rect 47696 39140 47752 39142
rect 47776 39140 47832 39142
rect 47856 39140 47912 39142
rect 52616 39194 52672 39196
rect 52696 39194 52752 39196
rect 52776 39194 52832 39196
rect 52856 39194 52912 39196
rect 52616 39142 52662 39194
rect 52662 39142 52672 39194
rect 52696 39142 52726 39194
rect 52726 39142 52738 39194
rect 52738 39142 52752 39194
rect 52776 39142 52790 39194
rect 52790 39142 52802 39194
rect 52802 39142 52832 39194
rect 52856 39142 52866 39194
rect 52866 39142 52912 39194
rect 52616 39140 52672 39142
rect 52696 39140 52752 39142
rect 52776 39140 52832 39142
rect 52856 39140 52912 39142
rect 57616 39194 57672 39196
rect 57696 39194 57752 39196
rect 57776 39194 57832 39196
rect 57856 39194 57912 39196
rect 57616 39142 57662 39194
rect 57662 39142 57672 39194
rect 57696 39142 57726 39194
rect 57726 39142 57738 39194
rect 57738 39142 57752 39194
rect 57776 39142 57790 39194
rect 57790 39142 57802 39194
rect 57802 39142 57832 39194
rect 57856 39142 57866 39194
rect 57866 39142 57912 39194
rect 57616 39140 57672 39142
rect 57696 39140 57752 39142
rect 57776 39140 57832 39142
rect 57856 39140 57912 39142
rect 1956 38650 2012 38652
rect 2036 38650 2092 38652
rect 2116 38650 2172 38652
rect 2196 38650 2252 38652
rect 1956 38598 2002 38650
rect 2002 38598 2012 38650
rect 2036 38598 2066 38650
rect 2066 38598 2078 38650
rect 2078 38598 2092 38650
rect 2116 38598 2130 38650
rect 2130 38598 2142 38650
rect 2142 38598 2172 38650
rect 2196 38598 2206 38650
rect 2206 38598 2252 38650
rect 1956 38596 2012 38598
rect 2036 38596 2092 38598
rect 2116 38596 2172 38598
rect 2196 38596 2252 38598
rect 6956 38650 7012 38652
rect 7036 38650 7092 38652
rect 7116 38650 7172 38652
rect 7196 38650 7252 38652
rect 6956 38598 7002 38650
rect 7002 38598 7012 38650
rect 7036 38598 7066 38650
rect 7066 38598 7078 38650
rect 7078 38598 7092 38650
rect 7116 38598 7130 38650
rect 7130 38598 7142 38650
rect 7142 38598 7172 38650
rect 7196 38598 7206 38650
rect 7206 38598 7252 38650
rect 6956 38596 7012 38598
rect 7036 38596 7092 38598
rect 7116 38596 7172 38598
rect 7196 38596 7252 38598
rect 11956 38650 12012 38652
rect 12036 38650 12092 38652
rect 12116 38650 12172 38652
rect 12196 38650 12252 38652
rect 11956 38598 12002 38650
rect 12002 38598 12012 38650
rect 12036 38598 12066 38650
rect 12066 38598 12078 38650
rect 12078 38598 12092 38650
rect 12116 38598 12130 38650
rect 12130 38598 12142 38650
rect 12142 38598 12172 38650
rect 12196 38598 12206 38650
rect 12206 38598 12252 38650
rect 11956 38596 12012 38598
rect 12036 38596 12092 38598
rect 12116 38596 12172 38598
rect 12196 38596 12252 38598
rect 16956 38650 17012 38652
rect 17036 38650 17092 38652
rect 17116 38650 17172 38652
rect 17196 38650 17252 38652
rect 16956 38598 17002 38650
rect 17002 38598 17012 38650
rect 17036 38598 17066 38650
rect 17066 38598 17078 38650
rect 17078 38598 17092 38650
rect 17116 38598 17130 38650
rect 17130 38598 17142 38650
rect 17142 38598 17172 38650
rect 17196 38598 17206 38650
rect 17206 38598 17252 38650
rect 16956 38596 17012 38598
rect 17036 38596 17092 38598
rect 17116 38596 17172 38598
rect 17196 38596 17252 38598
rect 21956 38650 22012 38652
rect 22036 38650 22092 38652
rect 22116 38650 22172 38652
rect 22196 38650 22252 38652
rect 21956 38598 22002 38650
rect 22002 38598 22012 38650
rect 22036 38598 22066 38650
rect 22066 38598 22078 38650
rect 22078 38598 22092 38650
rect 22116 38598 22130 38650
rect 22130 38598 22142 38650
rect 22142 38598 22172 38650
rect 22196 38598 22206 38650
rect 22206 38598 22252 38650
rect 21956 38596 22012 38598
rect 22036 38596 22092 38598
rect 22116 38596 22172 38598
rect 22196 38596 22252 38598
rect 26956 38650 27012 38652
rect 27036 38650 27092 38652
rect 27116 38650 27172 38652
rect 27196 38650 27252 38652
rect 26956 38598 27002 38650
rect 27002 38598 27012 38650
rect 27036 38598 27066 38650
rect 27066 38598 27078 38650
rect 27078 38598 27092 38650
rect 27116 38598 27130 38650
rect 27130 38598 27142 38650
rect 27142 38598 27172 38650
rect 27196 38598 27206 38650
rect 27206 38598 27252 38650
rect 26956 38596 27012 38598
rect 27036 38596 27092 38598
rect 27116 38596 27172 38598
rect 27196 38596 27252 38598
rect 31956 38650 32012 38652
rect 32036 38650 32092 38652
rect 32116 38650 32172 38652
rect 32196 38650 32252 38652
rect 31956 38598 32002 38650
rect 32002 38598 32012 38650
rect 32036 38598 32066 38650
rect 32066 38598 32078 38650
rect 32078 38598 32092 38650
rect 32116 38598 32130 38650
rect 32130 38598 32142 38650
rect 32142 38598 32172 38650
rect 32196 38598 32206 38650
rect 32206 38598 32252 38650
rect 31956 38596 32012 38598
rect 32036 38596 32092 38598
rect 32116 38596 32172 38598
rect 32196 38596 32252 38598
rect 36956 38650 37012 38652
rect 37036 38650 37092 38652
rect 37116 38650 37172 38652
rect 37196 38650 37252 38652
rect 36956 38598 37002 38650
rect 37002 38598 37012 38650
rect 37036 38598 37066 38650
rect 37066 38598 37078 38650
rect 37078 38598 37092 38650
rect 37116 38598 37130 38650
rect 37130 38598 37142 38650
rect 37142 38598 37172 38650
rect 37196 38598 37206 38650
rect 37206 38598 37252 38650
rect 36956 38596 37012 38598
rect 37036 38596 37092 38598
rect 37116 38596 37172 38598
rect 37196 38596 37252 38598
rect 41956 38650 42012 38652
rect 42036 38650 42092 38652
rect 42116 38650 42172 38652
rect 42196 38650 42252 38652
rect 41956 38598 42002 38650
rect 42002 38598 42012 38650
rect 42036 38598 42066 38650
rect 42066 38598 42078 38650
rect 42078 38598 42092 38650
rect 42116 38598 42130 38650
rect 42130 38598 42142 38650
rect 42142 38598 42172 38650
rect 42196 38598 42206 38650
rect 42206 38598 42252 38650
rect 41956 38596 42012 38598
rect 42036 38596 42092 38598
rect 42116 38596 42172 38598
rect 42196 38596 42252 38598
rect 46956 38650 47012 38652
rect 47036 38650 47092 38652
rect 47116 38650 47172 38652
rect 47196 38650 47252 38652
rect 46956 38598 47002 38650
rect 47002 38598 47012 38650
rect 47036 38598 47066 38650
rect 47066 38598 47078 38650
rect 47078 38598 47092 38650
rect 47116 38598 47130 38650
rect 47130 38598 47142 38650
rect 47142 38598 47172 38650
rect 47196 38598 47206 38650
rect 47206 38598 47252 38650
rect 46956 38596 47012 38598
rect 47036 38596 47092 38598
rect 47116 38596 47172 38598
rect 47196 38596 47252 38598
rect 51956 38650 52012 38652
rect 52036 38650 52092 38652
rect 52116 38650 52172 38652
rect 52196 38650 52252 38652
rect 51956 38598 52002 38650
rect 52002 38598 52012 38650
rect 52036 38598 52066 38650
rect 52066 38598 52078 38650
rect 52078 38598 52092 38650
rect 52116 38598 52130 38650
rect 52130 38598 52142 38650
rect 52142 38598 52172 38650
rect 52196 38598 52206 38650
rect 52206 38598 52252 38650
rect 51956 38596 52012 38598
rect 52036 38596 52092 38598
rect 52116 38596 52172 38598
rect 52196 38596 52252 38598
rect 56956 38650 57012 38652
rect 57036 38650 57092 38652
rect 57116 38650 57172 38652
rect 57196 38650 57252 38652
rect 56956 38598 57002 38650
rect 57002 38598 57012 38650
rect 57036 38598 57066 38650
rect 57066 38598 57078 38650
rect 57078 38598 57092 38650
rect 57116 38598 57130 38650
rect 57130 38598 57142 38650
rect 57142 38598 57172 38650
rect 57196 38598 57206 38650
rect 57206 38598 57252 38650
rect 56956 38596 57012 38598
rect 57036 38596 57092 38598
rect 57116 38596 57172 38598
rect 57196 38596 57252 38598
rect 58530 38392 58586 38448
rect 2616 38106 2672 38108
rect 2696 38106 2752 38108
rect 2776 38106 2832 38108
rect 2856 38106 2912 38108
rect 2616 38054 2662 38106
rect 2662 38054 2672 38106
rect 2696 38054 2726 38106
rect 2726 38054 2738 38106
rect 2738 38054 2752 38106
rect 2776 38054 2790 38106
rect 2790 38054 2802 38106
rect 2802 38054 2832 38106
rect 2856 38054 2866 38106
rect 2866 38054 2912 38106
rect 2616 38052 2672 38054
rect 2696 38052 2752 38054
rect 2776 38052 2832 38054
rect 2856 38052 2912 38054
rect 7616 38106 7672 38108
rect 7696 38106 7752 38108
rect 7776 38106 7832 38108
rect 7856 38106 7912 38108
rect 7616 38054 7662 38106
rect 7662 38054 7672 38106
rect 7696 38054 7726 38106
rect 7726 38054 7738 38106
rect 7738 38054 7752 38106
rect 7776 38054 7790 38106
rect 7790 38054 7802 38106
rect 7802 38054 7832 38106
rect 7856 38054 7866 38106
rect 7866 38054 7912 38106
rect 7616 38052 7672 38054
rect 7696 38052 7752 38054
rect 7776 38052 7832 38054
rect 7856 38052 7912 38054
rect 12616 38106 12672 38108
rect 12696 38106 12752 38108
rect 12776 38106 12832 38108
rect 12856 38106 12912 38108
rect 12616 38054 12662 38106
rect 12662 38054 12672 38106
rect 12696 38054 12726 38106
rect 12726 38054 12738 38106
rect 12738 38054 12752 38106
rect 12776 38054 12790 38106
rect 12790 38054 12802 38106
rect 12802 38054 12832 38106
rect 12856 38054 12866 38106
rect 12866 38054 12912 38106
rect 12616 38052 12672 38054
rect 12696 38052 12752 38054
rect 12776 38052 12832 38054
rect 12856 38052 12912 38054
rect 17616 38106 17672 38108
rect 17696 38106 17752 38108
rect 17776 38106 17832 38108
rect 17856 38106 17912 38108
rect 17616 38054 17662 38106
rect 17662 38054 17672 38106
rect 17696 38054 17726 38106
rect 17726 38054 17738 38106
rect 17738 38054 17752 38106
rect 17776 38054 17790 38106
rect 17790 38054 17802 38106
rect 17802 38054 17832 38106
rect 17856 38054 17866 38106
rect 17866 38054 17912 38106
rect 17616 38052 17672 38054
rect 17696 38052 17752 38054
rect 17776 38052 17832 38054
rect 17856 38052 17912 38054
rect 22616 38106 22672 38108
rect 22696 38106 22752 38108
rect 22776 38106 22832 38108
rect 22856 38106 22912 38108
rect 22616 38054 22662 38106
rect 22662 38054 22672 38106
rect 22696 38054 22726 38106
rect 22726 38054 22738 38106
rect 22738 38054 22752 38106
rect 22776 38054 22790 38106
rect 22790 38054 22802 38106
rect 22802 38054 22832 38106
rect 22856 38054 22866 38106
rect 22866 38054 22912 38106
rect 22616 38052 22672 38054
rect 22696 38052 22752 38054
rect 22776 38052 22832 38054
rect 22856 38052 22912 38054
rect 27616 38106 27672 38108
rect 27696 38106 27752 38108
rect 27776 38106 27832 38108
rect 27856 38106 27912 38108
rect 27616 38054 27662 38106
rect 27662 38054 27672 38106
rect 27696 38054 27726 38106
rect 27726 38054 27738 38106
rect 27738 38054 27752 38106
rect 27776 38054 27790 38106
rect 27790 38054 27802 38106
rect 27802 38054 27832 38106
rect 27856 38054 27866 38106
rect 27866 38054 27912 38106
rect 27616 38052 27672 38054
rect 27696 38052 27752 38054
rect 27776 38052 27832 38054
rect 27856 38052 27912 38054
rect 32616 38106 32672 38108
rect 32696 38106 32752 38108
rect 32776 38106 32832 38108
rect 32856 38106 32912 38108
rect 32616 38054 32662 38106
rect 32662 38054 32672 38106
rect 32696 38054 32726 38106
rect 32726 38054 32738 38106
rect 32738 38054 32752 38106
rect 32776 38054 32790 38106
rect 32790 38054 32802 38106
rect 32802 38054 32832 38106
rect 32856 38054 32866 38106
rect 32866 38054 32912 38106
rect 32616 38052 32672 38054
rect 32696 38052 32752 38054
rect 32776 38052 32832 38054
rect 32856 38052 32912 38054
rect 37616 38106 37672 38108
rect 37696 38106 37752 38108
rect 37776 38106 37832 38108
rect 37856 38106 37912 38108
rect 37616 38054 37662 38106
rect 37662 38054 37672 38106
rect 37696 38054 37726 38106
rect 37726 38054 37738 38106
rect 37738 38054 37752 38106
rect 37776 38054 37790 38106
rect 37790 38054 37802 38106
rect 37802 38054 37832 38106
rect 37856 38054 37866 38106
rect 37866 38054 37912 38106
rect 37616 38052 37672 38054
rect 37696 38052 37752 38054
rect 37776 38052 37832 38054
rect 37856 38052 37912 38054
rect 42616 38106 42672 38108
rect 42696 38106 42752 38108
rect 42776 38106 42832 38108
rect 42856 38106 42912 38108
rect 42616 38054 42662 38106
rect 42662 38054 42672 38106
rect 42696 38054 42726 38106
rect 42726 38054 42738 38106
rect 42738 38054 42752 38106
rect 42776 38054 42790 38106
rect 42790 38054 42802 38106
rect 42802 38054 42832 38106
rect 42856 38054 42866 38106
rect 42866 38054 42912 38106
rect 42616 38052 42672 38054
rect 42696 38052 42752 38054
rect 42776 38052 42832 38054
rect 42856 38052 42912 38054
rect 47616 38106 47672 38108
rect 47696 38106 47752 38108
rect 47776 38106 47832 38108
rect 47856 38106 47912 38108
rect 47616 38054 47662 38106
rect 47662 38054 47672 38106
rect 47696 38054 47726 38106
rect 47726 38054 47738 38106
rect 47738 38054 47752 38106
rect 47776 38054 47790 38106
rect 47790 38054 47802 38106
rect 47802 38054 47832 38106
rect 47856 38054 47866 38106
rect 47866 38054 47912 38106
rect 47616 38052 47672 38054
rect 47696 38052 47752 38054
rect 47776 38052 47832 38054
rect 47856 38052 47912 38054
rect 52616 38106 52672 38108
rect 52696 38106 52752 38108
rect 52776 38106 52832 38108
rect 52856 38106 52912 38108
rect 52616 38054 52662 38106
rect 52662 38054 52672 38106
rect 52696 38054 52726 38106
rect 52726 38054 52738 38106
rect 52738 38054 52752 38106
rect 52776 38054 52790 38106
rect 52790 38054 52802 38106
rect 52802 38054 52832 38106
rect 52856 38054 52866 38106
rect 52866 38054 52912 38106
rect 52616 38052 52672 38054
rect 52696 38052 52752 38054
rect 52776 38052 52832 38054
rect 52856 38052 52912 38054
rect 57616 38106 57672 38108
rect 57696 38106 57752 38108
rect 57776 38106 57832 38108
rect 57856 38106 57912 38108
rect 57616 38054 57662 38106
rect 57662 38054 57672 38106
rect 57696 38054 57726 38106
rect 57726 38054 57738 38106
rect 57738 38054 57752 38106
rect 57776 38054 57790 38106
rect 57790 38054 57802 38106
rect 57802 38054 57832 38106
rect 57856 38054 57866 38106
rect 57866 38054 57912 38106
rect 57616 38052 57672 38054
rect 57696 38052 57752 38054
rect 57776 38052 57832 38054
rect 57856 38052 57912 38054
rect 58530 37612 58532 37632
rect 58532 37612 58584 37632
rect 58584 37612 58586 37632
rect 58530 37576 58586 37612
rect 1956 37562 2012 37564
rect 2036 37562 2092 37564
rect 2116 37562 2172 37564
rect 2196 37562 2252 37564
rect 1956 37510 2002 37562
rect 2002 37510 2012 37562
rect 2036 37510 2066 37562
rect 2066 37510 2078 37562
rect 2078 37510 2092 37562
rect 2116 37510 2130 37562
rect 2130 37510 2142 37562
rect 2142 37510 2172 37562
rect 2196 37510 2206 37562
rect 2206 37510 2252 37562
rect 1956 37508 2012 37510
rect 2036 37508 2092 37510
rect 2116 37508 2172 37510
rect 2196 37508 2252 37510
rect 6956 37562 7012 37564
rect 7036 37562 7092 37564
rect 7116 37562 7172 37564
rect 7196 37562 7252 37564
rect 6956 37510 7002 37562
rect 7002 37510 7012 37562
rect 7036 37510 7066 37562
rect 7066 37510 7078 37562
rect 7078 37510 7092 37562
rect 7116 37510 7130 37562
rect 7130 37510 7142 37562
rect 7142 37510 7172 37562
rect 7196 37510 7206 37562
rect 7206 37510 7252 37562
rect 6956 37508 7012 37510
rect 7036 37508 7092 37510
rect 7116 37508 7172 37510
rect 7196 37508 7252 37510
rect 11956 37562 12012 37564
rect 12036 37562 12092 37564
rect 12116 37562 12172 37564
rect 12196 37562 12252 37564
rect 11956 37510 12002 37562
rect 12002 37510 12012 37562
rect 12036 37510 12066 37562
rect 12066 37510 12078 37562
rect 12078 37510 12092 37562
rect 12116 37510 12130 37562
rect 12130 37510 12142 37562
rect 12142 37510 12172 37562
rect 12196 37510 12206 37562
rect 12206 37510 12252 37562
rect 11956 37508 12012 37510
rect 12036 37508 12092 37510
rect 12116 37508 12172 37510
rect 12196 37508 12252 37510
rect 16956 37562 17012 37564
rect 17036 37562 17092 37564
rect 17116 37562 17172 37564
rect 17196 37562 17252 37564
rect 16956 37510 17002 37562
rect 17002 37510 17012 37562
rect 17036 37510 17066 37562
rect 17066 37510 17078 37562
rect 17078 37510 17092 37562
rect 17116 37510 17130 37562
rect 17130 37510 17142 37562
rect 17142 37510 17172 37562
rect 17196 37510 17206 37562
rect 17206 37510 17252 37562
rect 16956 37508 17012 37510
rect 17036 37508 17092 37510
rect 17116 37508 17172 37510
rect 17196 37508 17252 37510
rect 21956 37562 22012 37564
rect 22036 37562 22092 37564
rect 22116 37562 22172 37564
rect 22196 37562 22252 37564
rect 21956 37510 22002 37562
rect 22002 37510 22012 37562
rect 22036 37510 22066 37562
rect 22066 37510 22078 37562
rect 22078 37510 22092 37562
rect 22116 37510 22130 37562
rect 22130 37510 22142 37562
rect 22142 37510 22172 37562
rect 22196 37510 22206 37562
rect 22206 37510 22252 37562
rect 21956 37508 22012 37510
rect 22036 37508 22092 37510
rect 22116 37508 22172 37510
rect 22196 37508 22252 37510
rect 26956 37562 27012 37564
rect 27036 37562 27092 37564
rect 27116 37562 27172 37564
rect 27196 37562 27252 37564
rect 26956 37510 27002 37562
rect 27002 37510 27012 37562
rect 27036 37510 27066 37562
rect 27066 37510 27078 37562
rect 27078 37510 27092 37562
rect 27116 37510 27130 37562
rect 27130 37510 27142 37562
rect 27142 37510 27172 37562
rect 27196 37510 27206 37562
rect 27206 37510 27252 37562
rect 26956 37508 27012 37510
rect 27036 37508 27092 37510
rect 27116 37508 27172 37510
rect 27196 37508 27252 37510
rect 31956 37562 32012 37564
rect 32036 37562 32092 37564
rect 32116 37562 32172 37564
rect 32196 37562 32252 37564
rect 31956 37510 32002 37562
rect 32002 37510 32012 37562
rect 32036 37510 32066 37562
rect 32066 37510 32078 37562
rect 32078 37510 32092 37562
rect 32116 37510 32130 37562
rect 32130 37510 32142 37562
rect 32142 37510 32172 37562
rect 32196 37510 32206 37562
rect 32206 37510 32252 37562
rect 31956 37508 32012 37510
rect 32036 37508 32092 37510
rect 32116 37508 32172 37510
rect 32196 37508 32252 37510
rect 36956 37562 37012 37564
rect 37036 37562 37092 37564
rect 37116 37562 37172 37564
rect 37196 37562 37252 37564
rect 36956 37510 37002 37562
rect 37002 37510 37012 37562
rect 37036 37510 37066 37562
rect 37066 37510 37078 37562
rect 37078 37510 37092 37562
rect 37116 37510 37130 37562
rect 37130 37510 37142 37562
rect 37142 37510 37172 37562
rect 37196 37510 37206 37562
rect 37206 37510 37252 37562
rect 36956 37508 37012 37510
rect 37036 37508 37092 37510
rect 37116 37508 37172 37510
rect 37196 37508 37252 37510
rect 41956 37562 42012 37564
rect 42036 37562 42092 37564
rect 42116 37562 42172 37564
rect 42196 37562 42252 37564
rect 41956 37510 42002 37562
rect 42002 37510 42012 37562
rect 42036 37510 42066 37562
rect 42066 37510 42078 37562
rect 42078 37510 42092 37562
rect 42116 37510 42130 37562
rect 42130 37510 42142 37562
rect 42142 37510 42172 37562
rect 42196 37510 42206 37562
rect 42206 37510 42252 37562
rect 41956 37508 42012 37510
rect 42036 37508 42092 37510
rect 42116 37508 42172 37510
rect 42196 37508 42252 37510
rect 46956 37562 47012 37564
rect 47036 37562 47092 37564
rect 47116 37562 47172 37564
rect 47196 37562 47252 37564
rect 46956 37510 47002 37562
rect 47002 37510 47012 37562
rect 47036 37510 47066 37562
rect 47066 37510 47078 37562
rect 47078 37510 47092 37562
rect 47116 37510 47130 37562
rect 47130 37510 47142 37562
rect 47142 37510 47172 37562
rect 47196 37510 47206 37562
rect 47206 37510 47252 37562
rect 46956 37508 47012 37510
rect 47036 37508 47092 37510
rect 47116 37508 47172 37510
rect 47196 37508 47252 37510
rect 51956 37562 52012 37564
rect 52036 37562 52092 37564
rect 52116 37562 52172 37564
rect 52196 37562 52252 37564
rect 51956 37510 52002 37562
rect 52002 37510 52012 37562
rect 52036 37510 52066 37562
rect 52066 37510 52078 37562
rect 52078 37510 52092 37562
rect 52116 37510 52130 37562
rect 52130 37510 52142 37562
rect 52142 37510 52172 37562
rect 52196 37510 52206 37562
rect 52206 37510 52252 37562
rect 51956 37508 52012 37510
rect 52036 37508 52092 37510
rect 52116 37508 52172 37510
rect 52196 37508 52252 37510
rect 56956 37562 57012 37564
rect 57036 37562 57092 37564
rect 57116 37562 57172 37564
rect 57196 37562 57252 37564
rect 56956 37510 57002 37562
rect 57002 37510 57012 37562
rect 57036 37510 57066 37562
rect 57066 37510 57078 37562
rect 57078 37510 57092 37562
rect 57116 37510 57130 37562
rect 57130 37510 57142 37562
rect 57142 37510 57172 37562
rect 57196 37510 57206 37562
rect 57206 37510 57252 37562
rect 56956 37508 57012 37510
rect 57036 37508 57092 37510
rect 57116 37508 57172 37510
rect 57196 37508 57252 37510
rect 2616 37018 2672 37020
rect 2696 37018 2752 37020
rect 2776 37018 2832 37020
rect 2856 37018 2912 37020
rect 2616 36966 2662 37018
rect 2662 36966 2672 37018
rect 2696 36966 2726 37018
rect 2726 36966 2738 37018
rect 2738 36966 2752 37018
rect 2776 36966 2790 37018
rect 2790 36966 2802 37018
rect 2802 36966 2832 37018
rect 2856 36966 2866 37018
rect 2866 36966 2912 37018
rect 2616 36964 2672 36966
rect 2696 36964 2752 36966
rect 2776 36964 2832 36966
rect 2856 36964 2912 36966
rect 7616 37018 7672 37020
rect 7696 37018 7752 37020
rect 7776 37018 7832 37020
rect 7856 37018 7912 37020
rect 7616 36966 7662 37018
rect 7662 36966 7672 37018
rect 7696 36966 7726 37018
rect 7726 36966 7738 37018
rect 7738 36966 7752 37018
rect 7776 36966 7790 37018
rect 7790 36966 7802 37018
rect 7802 36966 7832 37018
rect 7856 36966 7866 37018
rect 7866 36966 7912 37018
rect 7616 36964 7672 36966
rect 7696 36964 7752 36966
rect 7776 36964 7832 36966
rect 7856 36964 7912 36966
rect 12616 37018 12672 37020
rect 12696 37018 12752 37020
rect 12776 37018 12832 37020
rect 12856 37018 12912 37020
rect 12616 36966 12662 37018
rect 12662 36966 12672 37018
rect 12696 36966 12726 37018
rect 12726 36966 12738 37018
rect 12738 36966 12752 37018
rect 12776 36966 12790 37018
rect 12790 36966 12802 37018
rect 12802 36966 12832 37018
rect 12856 36966 12866 37018
rect 12866 36966 12912 37018
rect 12616 36964 12672 36966
rect 12696 36964 12752 36966
rect 12776 36964 12832 36966
rect 12856 36964 12912 36966
rect 17616 37018 17672 37020
rect 17696 37018 17752 37020
rect 17776 37018 17832 37020
rect 17856 37018 17912 37020
rect 17616 36966 17662 37018
rect 17662 36966 17672 37018
rect 17696 36966 17726 37018
rect 17726 36966 17738 37018
rect 17738 36966 17752 37018
rect 17776 36966 17790 37018
rect 17790 36966 17802 37018
rect 17802 36966 17832 37018
rect 17856 36966 17866 37018
rect 17866 36966 17912 37018
rect 17616 36964 17672 36966
rect 17696 36964 17752 36966
rect 17776 36964 17832 36966
rect 17856 36964 17912 36966
rect 22616 37018 22672 37020
rect 22696 37018 22752 37020
rect 22776 37018 22832 37020
rect 22856 37018 22912 37020
rect 22616 36966 22662 37018
rect 22662 36966 22672 37018
rect 22696 36966 22726 37018
rect 22726 36966 22738 37018
rect 22738 36966 22752 37018
rect 22776 36966 22790 37018
rect 22790 36966 22802 37018
rect 22802 36966 22832 37018
rect 22856 36966 22866 37018
rect 22866 36966 22912 37018
rect 22616 36964 22672 36966
rect 22696 36964 22752 36966
rect 22776 36964 22832 36966
rect 22856 36964 22912 36966
rect 27616 37018 27672 37020
rect 27696 37018 27752 37020
rect 27776 37018 27832 37020
rect 27856 37018 27912 37020
rect 27616 36966 27662 37018
rect 27662 36966 27672 37018
rect 27696 36966 27726 37018
rect 27726 36966 27738 37018
rect 27738 36966 27752 37018
rect 27776 36966 27790 37018
rect 27790 36966 27802 37018
rect 27802 36966 27832 37018
rect 27856 36966 27866 37018
rect 27866 36966 27912 37018
rect 27616 36964 27672 36966
rect 27696 36964 27752 36966
rect 27776 36964 27832 36966
rect 27856 36964 27912 36966
rect 32616 37018 32672 37020
rect 32696 37018 32752 37020
rect 32776 37018 32832 37020
rect 32856 37018 32912 37020
rect 32616 36966 32662 37018
rect 32662 36966 32672 37018
rect 32696 36966 32726 37018
rect 32726 36966 32738 37018
rect 32738 36966 32752 37018
rect 32776 36966 32790 37018
rect 32790 36966 32802 37018
rect 32802 36966 32832 37018
rect 32856 36966 32866 37018
rect 32866 36966 32912 37018
rect 32616 36964 32672 36966
rect 32696 36964 32752 36966
rect 32776 36964 32832 36966
rect 32856 36964 32912 36966
rect 37616 37018 37672 37020
rect 37696 37018 37752 37020
rect 37776 37018 37832 37020
rect 37856 37018 37912 37020
rect 37616 36966 37662 37018
rect 37662 36966 37672 37018
rect 37696 36966 37726 37018
rect 37726 36966 37738 37018
rect 37738 36966 37752 37018
rect 37776 36966 37790 37018
rect 37790 36966 37802 37018
rect 37802 36966 37832 37018
rect 37856 36966 37866 37018
rect 37866 36966 37912 37018
rect 37616 36964 37672 36966
rect 37696 36964 37752 36966
rect 37776 36964 37832 36966
rect 37856 36964 37912 36966
rect 42616 37018 42672 37020
rect 42696 37018 42752 37020
rect 42776 37018 42832 37020
rect 42856 37018 42912 37020
rect 42616 36966 42662 37018
rect 42662 36966 42672 37018
rect 42696 36966 42726 37018
rect 42726 36966 42738 37018
rect 42738 36966 42752 37018
rect 42776 36966 42790 37018
rect 42790 36966 42802 37018
rect 42802 36966 42832 37018
rect 42856 36966 42866 37018
rect 42866 36966 42912 37018
rect 42616 36964 42672 36966
rect 42696 36964 42752 36966
rect 42776 36964 42832 36966
rect 42856 36964 42912 36966
rect 47616 37018 47672 37020
rect 47696 37018 47752 37020
rect 47776 37018 47832 37020
rect 47856 37018 47912 37020
rect 47616 36966 47662 37018
rect 47662 36966 47672 37018
rect 47696 36966 47726 37018
rect 47726 36966 47738 37018
rect 47738 36966 47752 37018
rect 47776 36966 47790 37018
rect 47790 36966 47802 37018
rect 47802 36966 47832 37018
rect 47856 36966 47866 37018
rect 47866 36966 47912 37018
rect 47616 36964 47672 36966
rect 47696 36964 47752 36966
rect 47776 36964 47832 36966
rect 47856 36964 47912 36966
rect 52616 37018 52672 37020
rect 52696 37018 52752 37020
rect 52776 37018 52832 37020
rect 52856 37018 52912 37020
rect 52616 36966 52662 37018
rect 52662 36966 52672 37018
rect 52696 36966 52726 37018
rect 52726 36966 52738 37018
rect 52738 36966 52752 37018
rect 52776 36966 52790 37018
rect 52790 36966 52802 37018
rect 52802 36966 52832 37018
rect 52856 36966 52866 37018
rect 52866 36966 52912 37018
rect 52616 36964 52672 36966
rect 52696 36964 52752 36966
rect 52776 36964 52832 36966
rect 52856 36964 52912 36966
rect 57616 37018 57672 37020
rect 57696 37018 57752 37020
rect 57776 37018 57832 37020
rect 57856 37018 57912 37020
rect 57616 36966 57662 37018
rect 57662 36966 57672 37018
rect 57696 36966 57726 37018
rect 57726 36966 57738 37018
rect 57738 36966 57752 37018
rect 57776 36966 57790 37018
rect 57790 36966 57802 37018
rect 57802 36966 57832 37018
rect 57856 36966 57866 37018
rect 57866 36966 57912 37018
rect 57616 36964 57672 36966
rect 57696 36964 57752 36966
rect 57776 36964 57832 36966
rect 57856 36964 57912 36966
rect 58530 36760 58586 36816
rect 1956 36474 2012 36476
rect 2036 36474 2092 36476
rect 2116 36474 2172 36476
rect 2196 36474 2252 36476
rect 1956 36422 2002 36474
rect 2002 36422 2012 36474
rect 2036 36422 2066 36474
rect 2066 36422 2078 36474
rect 2078 36422 2092 36474
rect 2116 36422 2130 36474
rect 2130 36422 2142 36474
rect 2142 36422 2172 36474
rect 2196 36422 2206 36474
rect 2206 36422 2252 36474
rect 1956 36420 2012 36422
rect 2036 36420 2092 36422
rect 2116 36420 2172 36422
rect 2196 36420 2252 36422
rect 6956 36474 7012 36476
rect 7036 36474 7092 36476
rect 7116 36474 7172 36476
rect 7196 36474 7252 36476
rect 6956 36422 7002 36474
rect 7002 36422 7012 36474
rect 7036 36422 7066 36474
rect 7066 36422 7078 36474
rect 7078 36422 7092 36474
rect 7116 36422 7130 36474
rect 7130 36422 7142 36474
rect 7142 36422 7172 36474
rect 7196 36422 7206 36474
rect 7206 36422 7252 36474
rect 6956 36420 7012 36422
rect 7036 36420 7092 36422
rect 7116 36420 7172 36422
rect 7196 36420 7252 36422
rect 11956 36474 12012 36476
rect 12036 36474 12092 36476
rect 12116 36474 12172 36476
rect 12196 36474 12252 36476
rect 11956 36422 12002 36474
rect 12002 36422 12012 36474
rect 12036 36422 12066 36474
rect 12066 36422 12078 36474
rect 12078 36422 12092 36474
rect 12116 36422 12130 36474
rect 12130 36422 12142 36474
rect 12142 36422 12172 36474
rect 12196 36422 12206 36474
rect 12206 36422 12252 36474
rect 11956 36420 12012 36422
rect 12036 36420 12092 36422
rect 12116 36420 12172 36422
rect 12196 36420 12252 36422
rect 16956 36474 17012 36476
rect 17036 36474 17092 36476
rect 17116 36474 17172 36476
rect 17196 36474 17252 36476
rect 16956 36422 17002 36474
rect 17002 36422 17012 36474
rect 17036 36422 17066 36474
rect 17066 36422 17078 36474
rect 17078 36422 17092 36474
rect 17116 36422 17130 36474
rect 17130 36422 17142 36474
rect 17142 36422 17172 36474
rect 17196 36422 17206 36474
rect 17206 36422 17252 36474
rect 16956 36420 17012 36422
rect 17036 36420 17092 36422
rect 17116 36420 17172 36422
rect 17196 36420 17252 36422
rect 21956 36474 22012 36476
rect 22036 36474 22092 36476
rect 22116 36474 22172 36476
rect 22196 36474 22252 36476
rect 21956 36422 22002 36474
rect 22002 36422 22012 36474
rect 22036 36422 22066 36474
rect 22066 36422 22078 36474
rect 22078 36422 22092 36474
rect 22116 36422 22130 36474
rect 22130 36422 22142 36474
rect 22142 36422 22172 36474
rect 22196 36422 22206 36474
rect 22206 36422 22252 36474
rect 21956 36420 22012 36422
rect 22036 36420 22092 36422
rect 22116 36420 22172 36422
rect 22196 36420 22252 36422
rect 26956 36474 27012 36476
rect 27036 36474 27092 36476
rect 27116 36474 27172 36476
rect 27196 36474 27252 36476
rect 26956 36422 27002 36474
rect 27002 36422 27012 36474
rect 27036 36422 27066 36474
rect 27066 36422 27078 36474
rect 27078 36422 27092 36474
rect 27116 36422 27130 36474
rect 27130 36422 27142 36474
rect 27142 36422 27172 36474
rect 27196 36422 27206 36474
rect 27206 36422 27252 36474
rect 26956 36420 27012 36422
rect 27036 36420 27092 36422
rect 27116 36420 27172 36422
rect 27196 36420 27252 36422
rect 31956 36474 32012 36476
rect 32036 36474 32092 36476
rect 32116 36474 32172 36476
rect 32196 36474 32252 36476
rect 31956 36422 32002 36474
rect 32002 36422 32012 36474
rect 32036 36422 32066 36474
rect 32066 36422 32078 36474
rect 32078 36422 32092 36474
rect 32116 36422 32130 36474
rect 32130 36422 32142 36474
rect 32142 36422 32172 36474
rect 32196 36422 32206 36474
rect 32206 36422 32252 36474
rect 31956 36420 32012 36422
rect 32036 36420 32092 36422
rect 32116 36420 32172 36422
rect 32196 36420 32252 36422
rect 36956 36474 37012 36476
rect 37036 36474 37092 36476
rect 37116 36474 37172 36476
rect 37196 36474 37252 36476
rect 36956 36422 37002 36474
rect 37002 36422 37012 36474
rect 37036 36422 37066 36474
rect 37066 36422 37078 36474
rect 37078 36422 37092 36474
rect 37116 36422 37130 36474
rect 37130 36422 37142 36474
rect 37142 36422 37172 36474
rect 37196 36422 37206 36474
rect 37206 36422 37252 36474
rect 36956 36420 37012 36422
rect 37036 36420 37092 36422
rect 37116 36420 37172 36422
rect 37196 36420 37252 36422
rect 41956 36474 42012 36476
rect 42036 36474 42092 36476
rect 42116 36474 42172 36476
rect 42196 36474 42252 36476
rect 41956 36422 42002 36474
rect 42002 36422 42012 36474
rect 42036 36422 42066 36474
rect 42066 36422 42078 36474
rect 42078 36422 42092 36474
rect 42116 36422 42130 36474
rect 42130 36422 42142 36474
rect 42142 36422 42172 36474
rect 42196 36422 42206 36474
rect 42206 36422 42252 36474
rect 41956 36420 42012 36422
rect 42036 36420 42092 36422
rect 42116 36420 42172 36422
rect 42196 36420 42252 36422
rect 46956 36474 47012 36476
rect 47036 36474 47092 36476
rect 47116 36474 47172 36476
rect 47196 36474 47252 36476
rect 46956 36422 47002 36474
rect 47002 36422 47012 36474
rect 47036 36422 47066 36474
rect 47066 36422 47078 36474
rect 47078 36422 47092 36474
rect 47116 36422 47130 36474
rect 47130 36422 47142 36474
rect 47142 36422 47172 36474
rect 47196 36422 47206 36474
rect 47206 36422 47252 36474
rect 46956 36420 47012 36422
rect 47036 36420 47092 36422
rect 47116 36420 47172 36422
rect 47196 36420 47252 36422
rect 51956 36474 52012 36476
rect 52036 36474 52092 36476
rect 52116 36474 52172 36476
rect 52196 36474 52252 36476
rect 51956 36422 52002 36474
rect 52002 36422 52012 36474
rect 52036 36422 52066 36474
rect 52066 36422 52078 36474
rect 52078 36422 52092 36474
rect 52116 36422 52130 36474
rect 52130 36422 52142 36474
rect 52142 36422 52172 36474
rect 52196 36422 52206 36474
rect 52206 36422 52252 36474
rect 51956 36420 52012 36422
rect 52036 36420 52092 36422
rect 52116 36420 52172 36422
rect 52196 36420 52252 36422
rect 56956 36474 57012 36476
rect 57036 36474 57092 36476
rect 57116 36474 57172 36476
rect 57196 36474 57252 36476
rect 56956 36422 57002 36474
rect 57002 36422 57012 36474
rect 57036 36422 57066 36474
rect 57066 36422 57078 36474
rect 57078 36422 57092 36474
rect 57116 36422 57130 36474
rect 57130 36422 57142 36474
rect 57142 36422 57172 36474
rect 57196 36422 57206 36474
rect 57206 36422 57252 36474
rect 56956 36420 57012 36422
rect 57036 36420 57092 36422
rect 57116 36420 57172 36422
rect 57196 36420 57252 36422
rect 58530 35944 58586 36000
rect 2616 35930 2672 35932
rect 2696 35930 2752 35932
rect 2776 35930 2832 35932
rect 2856 35930 2912 35932
rect 2616 35878 2662 35930
rect 2662 35878 2672 35930
rect 2696 35878 2726 35930
rect 2726 35878 2738 35930
rect 2738 35878 2752 35930
rect 2776 35878 2790 35930
rect 2790 35878 2802 35930
rect 2802 35878 2832 35930
rect 2856 35878 2866 35930
rect 2866 35878 2912 35930
rect 2616 35876 2672 35878
rect 2696 35876 2752 35878
rect 2776 35876 2832 35878
rect 2856 35876 2912 35878
rect 7616 35930 7672 35932
rect 7696 35930 7752 35932
rect 7776 35930 7832 35932
rect 7856 35930 7912 35932
rect 7616 35878 7662 35930
rect 7662 35878 7672 35930
rect 7696 35878 7726 35930
rect 7726 35878 7738 35930
rect 7738 35878 7752 35930
rect 7776 35878 7790 35930
rect 7790 35878 7802 35930
rect 7802 35878 7832 35930
rect 7856 35878 7866 35930
rect 7866 35878 7912 35930
rect 7616 35876 7672 35878
rect 7696 35876 7752 35878
rect 7776 35876 7832 35878
rect 7856 35876 7912 35878
rect 12616 35930 12672 35932
rect 12696 35930 12752 35932
rect 12776 35930 12832 35932
rect 12856 35930 12912 35932
rect 12616 35878 12662 35930
rect 12662 35878 12672 35930
rect 12696 35878 12726 35930
rect 12726 35878 12738 35930
rect 12738 35878 12752 35930
rect 12776 35878 12790 35930
rect 12790 35878 12802 35930
rect 12802 35878 12832 35930
rect 12856 35878 12866 35930
rect 12866 35878 12912 35930
rect 12616 35876 12672 35878
rect 12696 35876 12752 35878
rect 12776 35876 12832 35878
rect 12856 35876 12912 35878
rect 17616 35930 17672 35932
rect 17696 35930 17752 35932
rect 17776 35930 17832 35932
rect 17856 35930 17912 35932
rect 17616 35878 17662 35930
rect 17662 35878 17672 35930
rect 17696 35878 17726 35930
rect 17726 35878 17738 35930
rect 17738 35878 17752 35930
rect 17776 35878 17790 35930
rect 17790 35878 17802 35930
rect 17802 35878 17832 35930
rect 17856 35878 17866 35930
rect 17866 35878 17912 35930
rect 17616 35876 17672 35878
rect 17696 35876 17752 35878
rect 17776 35876 17832 35878
rect 17856 35876 17912 35878
rect 22616 35930 22672 35932
rect 22696 35930 22752 35932
rect 22776 35930 22832 35932
rect 22856 35930 22912 35932
rect 22616 35878 22662 35930
rect 22662 35878 22672 35930
rect 22696 35878 22726 35930
rect 22726 35878 22738 35930
rect 22738 35878 22752 35930
rect 22776 35878 22790 35930
rect 22790 35878 22802 35930
rect 22802 35878 22832 35930
rect 22856 35878 22866 35930
rect 22866 35878 22912 35930
rect 22616 35876 22672 35878
rect 22696 35876 22752 35878
rect 22776 35876 22832 35878
rect 22856 35876 22912 35878
rect 27616 35930 27672 35932
rect 27696 35930 27752 35932
rect 27776 35930 27832 35932
rect 27856 35930 27912 35932
rect 27616 35878 27662 35930
rect 27662 35878 27672 35930
rect 27696 35878 27726 35930
rect 27726 35878 27738 35930
rect 27738 35878 27752 35930
rect 27776 35878 27790 35930
rect 27790 35878 27802 35930
rect 27802 35878 27832 35930
rect 27856 35878 27866 35930
rect 27866 35878 27912 35930
rect 27616 35876 27672 35878
rect 27696 35876 27752 35878
rect 27776 35876 27832 35878
rect 27856 35876 27912 35878
rect 32616 35930 32672 35932
rect 32696 35930 32752 35932
rect 32776 35930 32832 35932
rect 32856 35930 32912 35932
rect 32616 35878 32662 35930
rect 32662 35878 32672 35930
rect 32696 35878 32726 35930
rect 32726 35878 32738 35930
rect 32738 35878 32752 35930
rect 32776 35878 32790 35930
rect 32790 35878 32802 35930
rect 32802 35878 32832 35930
rect 32856 35878 32866 35930
rect 32866 35878 32912 35930
rect 32616 35876 32672 35878
rect 32696 35876 32752 35878
rect 32776 35876 32832 35878
rect 32856 35876 32912 35878
rect 37616 35930 37672 35932
rect 37696 35930 37752 35932
rect 37776 35930 37832 35932
rect 37856 35930 37912 35932
rect 37616 35878 37662 35930
rect 37662 35878 37672 35930
rect 37696 35878 37726 35930
rect 37726 35878 37738 35930
rect 37738 35878 37752 35930
rect 37776 35878 37790 35930
rect 37790 35878 37802 35930
rect 37802 35878 37832 35930
rect 37856 35878 37866 35930
rect 37866 35878 37912 35930
rect 37616 35876 37672 35878
rect 37696 35876 37752 35878
rect 37776 35876 37832 35878
rect 37856 35876 37912 35878
rect 42616 35930 42672 35932
rect 42696 35930 42752 35932
rect 42776 35930 42832 35932
rect 42856 35930 42912 35932
rect 42616 35878 42662 35930
rect 42662 35878 42672 35930
rect 42696 35878 42726 35930
rect 42726 35878 42738 35930
rect 42738 35878 42752 35930
rect 42776 35878 42790 35930
rect 42790 35878 42802 35930
rect 42802 35878 42832 35930
rect 42856 35878 42866 35930
rect 42866 35878 42912 35930
rect 42616 35876 42672 35878
rect 42696 35876 42752 35878
rect 42776 35876 42832 35878
rect 42856 35876 42912 35878
rect 47616 35930 47672 35932
rect 47696 35930 47752 35932
rect 47776 35930 47832 35932
rect 47856 35930 47912 35932
rect 47616 35878 47662 35930
rect 47662 35878 47672 35930
rect 47696 35878 47726 35930
rect 47726 35878 47738 35930
rect 47738 35878 47752 35930
rect 47776 35878 47790 35930
rect 47790 35878 47802 35930
rect 47802 35878 47832 35930
rect 47856 35878 47866 35930
rect 47866 35878 47912 35930
rect 47616 35876 47672 35878
rect 47696 35876 47752 35878
rect 47776 35876 47832 35878
rect 47856 35876 47912 35878
rect 52616 35930 52672 35932
rect 52696 35930 52752 35932
rect 52776 35930 52832 35932
rect 52856 35930 52912 35932
rect 52616 35878 52662 35930
rect 52662 35878 52672 35930
rect 52696 35878 52726 35930
rect 52726 35878 52738 35930
rect 52738 35878 52752 35930
rect 52776 35878 52790 35930
rect 52790 35878 52802 35930
rect 52802 35878 52832 35930
rect 52856 35878 52866 35930
rect 52866 35878 52912 35930
rect 52616 35876 52672 35878
rect 52696 35876 52752 35878
rect 52776 35876 52832 35878
rect 52856 35876 52912 35878
rect 57616 35930 57672 35932
rect 57696 35930 57752 35932
rect 57776 35930 57832 35932
rect 57856 35930 57912 35932
rect 57616 35878 57662 35930
rect 57662 35878 57672 35930
rect 57696 35878 57726 35930
rect 57726 35878 57738 35930
rect 57738 35878 57752 35930
rect 57776 35878 57790 35930
rect 57790 35878 57802 35930
rect 57802 35878 57832 35930
rect 57856 35878 57866 35930
rect 57866 35878 57912 35930
rect 57616 35876 57672 35878
rect 57696 35876 57752 35878
rect 57776 35876 57832 35878
rect 57856 35876 57912 35878
rect 1956 35386 2012 35388
rect 2036 35386 2092 35388
rect 2116 35386 2172 35388
rect 2196 35386 2252 35388
rect 1956 35334 2002 35386
rect 2002 35334 2012 35386
rect 2036 35334 2066 35386
rect 2066 35334 2078 35386
rect 2078 35334 2092 35386
rect 2116 35334 2130 35386
rect 2130 35334 2142 35386
rect 2142 35334 2172 35386
rect 2196 35334 2206 35386
rect 2206 35334 2252 35386
rect 1956 35332 2012 35334
rect 2036 35332 2092 35334
rect 2116 35332 2172 35334
rect 2196 35332 2252 35334
rect 6956 35386 7012 35388
rect 7036 35386 7092 35388
rect 7116 35386 7172 35388
rect 7196 35386 7252 35388
rect 6956 35334 7002 35386
rect 7002 35334 7012 35386
rect 7036 35334 7066 35386
rect 7066 35334 7078 35386
rect 7078 35334 7092 35386
rect 7116 35334 7130 35386
rect 7130 35334 7142 35386
rect 7142 35334 7172 35386
rect 7196 35334 7206 35386
rect 7206 35334 7252 35386
rect 6956 35332 7012 35334
rect 7036 35332 7092 35334
rect 7116 35332 7172 35334
rect 7196 35332 7252 35334
rect 11956 35386 12012 35388
rect 12036 35386 12092 35388
rect 12116 35386 12172 35388
rect 12196 35386 12252 35388
rect 11956 35334 12002 35386
rect 12002 35334 12012 35386
rect 12036 35334 12066 35386
rect 12066 35334 12078 35386
rect 12078 35334 12092 35386
rect 12116 35334 12130 35386
rect 12130 35334 12142 35386
rect 12142 35334 12172 35386
rect 12196 35334 12206 35386
rect 12206 35334 12252 35386
rect 11956 35332 12012 35334
rect 12036 35332 12092 35334
rect 12116 35332 12172 35334
rect 12196 35332 12252 35334
rect 16956 35386 17012 35388
rect 17036 35386 17092 35388
rect 17116 35386 17172 35388
rect 17196 35386 17252 35388
rect 16956 35334 17002 35386
rect 17002 35334 17012 35386
rect 17036 35334 17066 35386
rect 17066 35334 17078 35386
rect 17078 35334 17092 35386
rect 17116 35334 17130 35386
rect 17130 35334 17142 35386
rect 17142 35334 17172 35386
rect 17196 35334 17206 35386
rect 17206 35334 17252 35386
rect 16956 35332 17012 35334
rect 17036 35332 17092 35334
rect 17116 35332 17172 35334
rect 17196 35332 17252 35334
rect 21956 35386 22012 35388
rect 22036 35386 22092 35388
rect 22116 35386 22172 35388
rect 22196 35386 22252 35388
rect 21956 35334 22002 35386
rect 22002 35334 22012 35386
rect 22036 35334 22066 35386
rect 22066 35334 22078 35386
rect 22078 35334 22092 35386
rect 22116 35334 22130 35386
rect 22130 35334 22142 35386
rect 22142 35334 22172 35386
rect 22196 35334 22206 35386
rect 22206 35334 22252 35386
rect 21956 35332 22012 35334
rect 22036 35332 22092 35334
rect 22116 35332 22172 35334
rect 22196 35332 22252 35334
rect 26956 35386 27012 35388
rect 27036 35386 27092 35388
rect 27116 35386 27172 35388
rect 27196 35386 27252 35388
rect 26956 35334 27002 35386
rect 27002 35334 27012 35386
rect 27036 35334 27066 35386
rect 27066 35334 27078 35386
rect 27078 35334 27092 35386
rect 27116 35334 27130 35386
rect 27130 35334 27142 35386
rect 27142 35334 27172 35386
rect 27196 35334 27206 35386
rect 27206 35334 27252 35386
rect 26956 35332 27012 35334
rect 27036 35332 27092 35334
rect 27116 35332 27172 35334
rect 27196 35332 27252 35334
rect 31956 35386 32012 35388
rect 32036 35386 32092 35388
rect 32116 35386 32172 35388
rect 32196 35386 32252 35388
rect 31956 35334 32002 35386
rect 32002 35334 32012 35386
rect 32036 35334 32066 35386
rect 32066 35334 32078 35386
rect 32078 35334 32092 35386
rect 32116 35334 32130 35386
rect 32130 35334 32142 35386
rect 32142 35334 32172 35386
rect 32196 35334 32206 35386
rect 32206 35334 32252 35386
rect 31956 35332 32012 35334
rect 32036 35332 32092 35334
rect 32116 35332 32172 35334
rect 32196 35332 32252 35334
rect 36956 35386 37012 35388
rect 37036 35386 37092 35388
rect 37116 35386 37172 35388
rect 37196 35386 37252 35388
rect 36956 35334 37002 35386
rect 37002 35334 37012 35386
rect 37036 35334 37066 35386
rect 37066 35334 37078 35386
rect 37078 35334 37092 35386
rect 37116 35334 37130 35386
rect 37130 35334 37142 35386
rect 37142 35334 37172 35386
rect 37196 35334 37206 35386
rect 37206 35334 37252 35386
rect 36956 35332 37012 35334
rect 37036 35332 37092 35334
rect 37116 35332 37172 35334
rect 37196 35332 37252 35334
rect 41956 35386 42012 35388
rect 42036 35386 42092 35388
rect 42116 35386 42172 35388
rect 42196 35386 42252 35388
rect 41956 35334 42002 35386
rect 42002 35334 42012 35386
rect 42036 35334 42066 35386
rect 42066 35334 42078 35386
rect 42078 35334 42092 35386
rect 42116 35334 42130 35386
rect 42130 35334 42142 35386
rect 42142 35334 42172 35386
rect 42196 35334 42206 35386
rect 42206 35334 42252 35386
rect 41956 35332 42012 35334
rect 42036 35332 42092 35334
rect 42116 35332 42172 35334
rect 42196 35332 42252 35334
rect 46956 35386 47012 35388
rect 47036 35386 47092 35388
rect 47116 35386 47172 35388
rect 47196 35386 47252 35388
rect 46956 35334 47002 35386
rect 47002 35334 47012 35386
rect 47036 35334 47066 35386
rect 47066 35334 47078 35386
rect 47078 35334 47092 35386
rect 47116 35334 47130 35386
rect 47130 35334 47142 35386
rect 47142 35334 47172 35386
rect 47196 35334 47206 35386
rect 47206 35334 47252 35386
rect 46956 35332 47012 35334
rect 47036 35332 47092 35334
rect 47116 35332 47172 35334
rect 47196 35332 47252 35334
rect 51956 35386 52012 35388
rect 52036 35386 52092 35388
rect 52116 35386 52172 35388
rect 52196 35386 52252 35388
rect 51956 35334 52002 35386
rect 52002 35334 52012 35386
rect 52036 35334 52066 35386
rect 52066 35334 52078 35386
rect 52078 35334 52092 35386
rect 52116 35334 52130 35386
rect 52130 35334 52142 35386
rect 52142 35334 52172 35386
rect 52196 35334 52206 35386
rect 52206 35334 52252 35386
rect 51956 35332 52012 35334
rect 52036 35332 52092 35334
rect 52116 35332 52172 35334
rect 52196 35332 52252 35334
rect 56956 35386 57012 35388
rect 57036 35386 57092 35388
rect 57116 35386 57172 35388
rect 57196 35386 57252 35388
rect 56956 35334 57002 35386
rect 57002 35334 57012 35386
rect 57036 35334 57066 35386
rect 57066 35334 57078 35386
rect 57078 35334 57092 35386
rect 57116 35334 57130 35386
rect 57130 35334 57142 35386
rect 57142 35334 57172 35386
rect 57196 35334 57206 35386
rect 57206 35334 57252 35386
rect 56956 35332 57012 35334
rect 57036 35332 57092 35334
rect 57116 35332 57172 35334
rect 57196 35332 57252 35334
rect 58530 35128 58586 35184
rect 2616 34842 2672 34844
rect 2696 34842 2752 34844
rect 2776 34842 2832 34844
rect 2856 34842 2912 34844
rect 2616 34790 2662 34842
rect 2662 34790 2672 34842
rect 2696 34790 2726 34842
rect 2726 34790 2738 34842
rect 2738 34790 2752 34842
rect 2776 34790 2790 34842
rect 2790 34790 2802 34842
rect 2802 34790 2832 34842
rect 2856 34790 2866 34842
rect 2866 34790 2912 34842
rect 2616 34788 2672 34790
rect 2696 34788 2752 34790
rect 2776 34788 2832 34790
rect 2856 34788 2912 34790
rect 7616 34842 7672 34844
rect 7696 34842 7752 34844
rect 7776 34842 7832 34844
rect 7856 34842 7912 34844
rect 7616 34790 7662 34842
rect 7662 34790 7672 34842
rect 7696 34790 7726 34842
rect 7726 34790 7738 34842
rect 7738 34790 7752 34842
rect 7776 34790 7790 34842
rect 7790 34790 7802 34842
rect 7802 34790 7832 34842
rect 7856 34790 7866 34842
rect 7866 34790 7912 34842
rect 7616 34788 7672 34790
rect 7696 34788 7752 34790
rect 7776 34788 7832 34790
rect 7856 34788 7912 34790
rect 12616 34842 12672 34844
rect 12696 34842 12752 34844
rect 12776 34842 12832 34844
rect 12856 34842 12912 34844
rect 12616 34790 12662 34842
rect 12662 34790 12672 34842
rect 12696 34790 12726 34842
rect 12726 34790 12738 34842
rect 12738 34790 12752 34842
rect 12776 34790 12790 34842
rect 12790 34790 12802 34842
rect 12802 34790 12832 34842
rect 12856 34790 12866 34842
rect 12866 34790 12912 34842
rect 12616 34788 12672 34790
rect 12696 34788 12752 34790
rect 12776 34788 12832 34790
rect 12856 34788 12912 34790
rect 17616 34842 17672 34844
rect 17696 34842 17752 34844
rect 17776 34842 17832 34844
rect 17856 34842 17912 34844
rect 17616 34790 17662 34842
rect 17662 34790 17672 34842
rect 17696 34790 17726 34842
rect 17726 34790 17738 34842
rect 17738 34790 17752 34842
rect 17776 34790 17790 34842
rect 17790 34790 17802 34842
rect 17802 34790 17832 34842
rect 17856 34790 17866 34842
rect 17866 34790 17912 34842
rect 17616 34788 17672 34790
rect 17696 34788 17752 34790
rect 17776 34788 17832 34790
rect 17856 34788 17912 34790
rect 22616 34842 22672 34844
rect 22696 34842 22752 34844
rect 22776 34842 22832 34844
rect 22856 34842 22912 34844
rect 22616 34790 22662 34842
rect 22662 34790 22672 34842
rect 22696 34790 22726 34842
rect 22726 34790 22738 34842
rect 22738 34790 22752 34842
rect 22776 34790 22790 34842
rect 22790 34790 22802 34842
rect 22802 34790 22832 34842
rect 22856 34790 22866 34842
rect 22866 34790 22912 34842
rect 22616 34788 22672 34790
rect 22696 34788 22752 34790
rect 22776 34788 22832 34790
rect 22856 34788 22912 34790
rect 27616 34842 27672 34844
rect 27696 34842 27752 34844
rect 27776 34842 27832 34844
rect 27856 34842 27912 34844
rect 27616 34790 27662 34842
rect 27662 34790 27672 34842
rect 27696 34790 27726 34842
rect 27726 34790 27738 34842
rect 27738 34790 27752 34842
rect 27776 34790 27790 34842
rect 27790 34790 27802 34842
rect 27802 34790 27832 34842
rect 27856 34790 27866 34842
rect 27866 34790 27912 34842
rect 27616 34788 27672 34790
rect 27696 34788 27752 34790
rect 27776 34788 27832 34790
rect 27856 34788 27912 34790
rect 32616 34842 32672 34844
rect 32696 34842 32752 34844
rect 32776 34842 32832 34844
rect 32856 34842 32912 34844
rect 32616 34790 32662 34842
rect 32662 34790 32672 34842
rect 32696 34790 32726 34842
rect 32726 34790 32738 34842
rect 32738 34790 32752 34842
rect 32776 34790 32790 34842
rect 32790 34790 32802 34842
rect 32802 34790 32832 34842
rect 32856 34790 32866 34842
rect 32866 34790 32912 34842
rect 32616 34788 32672 34790
rect 32696 34788 32752 34790
rect 32776 34788 32832 34790
rect 32856 34788 32912 34790
rect 37616 34842 37672 34844
rect 37696 34842 37752 34844
rect 37776 34842 37832 34844
rect 37856 34842 37912 34844
rect 37616 34790 37662 34842
rect 37662 34790 37672 34842
rect 37696 34790 37726 34842
rect 37726 34790 37738 34842
rect 37738 34790 37752 34842
rect 37776 34790 37790 34842
rect 37790 34790 37802 34842
rect 37802 34790 37832 34842
rect 37856 34790 37866 34842
rect 37866 34790 37912 34842
rect 37616 34788 37672 34790
rect 37696 34788 37752 34790
rect 37776 34788 37832 34790
rect 37856 34788 37912 34790
rect 42616 34842 42672 34844
rect 42696 34842 42752 34844
rect 42776 34842 42832 34844
rect 42856 34842 42912 34844
rect 42616 34790 42662 34842
rect 42662 34790 42672 34842
rect 42696 34790 42726 34842
rect 42726 34790 42738 34842
rect 42738 34790 42752 34842
rect 42776 34790 42790 34842
rect 42790 34790 42802 34842
rect 42802 34790 42832 34842
rect 42856 34790 42866 34842
rect 42866 34790 42912 34842
rect 42616 34788 42672 34790
rect 42696 34788 42752 34790
rect 42776 34788 42832 34790
rect 42856 34788 42912 34790
rect 47616 34842 47672 34844
rect 47696 34842 47752 34844
rect 47776 34842 47832 34844
rect 47856 34842 47912 34844
rect 47616 34790 47662 34842
rect 47662 34790 47672 34842
rect 47696 34790 47726 34842
rect 47726 34790 47738 34842
rect 47738 34790 47752 34842
rect 47776 34790 47790 34842
rect 47790 34790 47802 34842
rect 47802 34790 47832 34842
rect 47856 34790 47866 34842
rect 47866 34790 47912 34842
rect 47616 34788 47672 34790
rect 47696 34788 47752 34790
rect 47776 34788 47832 34790
rect 47856 34788 47912 34790
rect 52616 34842 52672 34844
rect 52696 34842 52752 34844
rect 52776 34842 52832 34844
rect 52856 34842 52912 34844
rect 52616 34790 52662 34842
rect 52662 34790 52672 34842
rect 52696 34790 52726 34842
rect 52726 34790 52738 34842
rect 52738 34790 52752 34842
rect 52776 34790 52790 34842
rect 52790 34790 52802 34842
rect 52802 34790 52832 34842
rect 52856 34790 52866 34842
rect 52866 34790 52912 34842
rect 52616 34788 52672 34790
rect 52696 34788 52752 34790
rect 52776 34788 52832 34790
rect 52856 34788 52912 34790
rect 57616 34842 57672 34844
rect 57696 34842 57752 34844
rect 57776 34842 57832 34844
rect 57856 34842 57912 34844
rect 57616 34790 57662 34842
rect 57662 34790 57672 34842
rect 57696 34790 57726 34842
rect 57726 34790 57738 34842
rect 57738 34790 57752 34842
rect 57776 34790 57790 34842
rect 57790 34790 57802 34842
rect 57802 34790 57832 34842
rect 57856 34790 57866 34842
rect 57866 34790 57912 34842
rect 57616 34788 57672 34790
rect 57696 34788 57752 34790
rect 57776 34788 57832 34790
rect 57856 34788 57912 34790
rect 58530 34348 58532 34368
rect 58532 34348 58584 34368
rect 58584 34348 58586 34368
rect 58530 34312 58586 34348
rect 1956 34298 2012 34300
rect 2036 34298 2092 34300
rect 2116 34298 2172 34300
rect 2196 34298 2252 34300
rect 1956 34246 2002 34298
rect 2002 34246 2012 34298
rect 2036 34246 2066 34298
rect 2066 34246 2078 34298
rect 2078 34246 2092 34298
rect 2116 34246 2130 34298
rect 2130 34246 2142 34298
rect 2142 34246 2172 34298
rect 2196 34246 2206 34298
rect 2206 34246 2252 34298
rect 1956 34244 2012 34246
rect 2036 34244 2092 34246
rect 2116 34244 2172 34246
rect 2196 34244 2252 34246
rect 6956 34298 7012 34300
rect 7036 34298 7092 34300
rect 7116 34298 7172 34300
rect 7196 34298 7252 34300
rect 6956 34246 7002 34298
rect 7002 34246 7012 34298
rect 7036 34246 7066 34298
rect 7066 34246 7078 34298
rect 7078 34246 7092 34298
rect 7116 34246 7130 34298
rect 7130 34246 7142 34298
rect 7142 34246 7172 34298
rect 7196 34246 7206 34298
rect 7206 34246 7252 34298
rect 6956 34244 7012 34246
rect 7036 34244 7092 34246
rect 7116 34244 7172 34246
rect 7196 34244 7252 34246
rect 11956 34298 12012 34300
rect 12036 34298 12092 34300
rect 12116 34298 12172 34300
rect 12196 34298 12252 34300
rect 11956 34246 12002 34298
rect 12002 34246 12012 34298
rect 12036 34246 12066 34298
rect 12066 34246 12078 34298
rect 12078 34246 12092 34298
rect 12116 34246 12130 34298
rect 12130 34246 12142 34298
rect 12142 34246 12172 34298
rect 12196 34246 12206 34298
rect 12206 34246 12252 34298
rect 11956 34244 12012 34246
rect 12036 34244 12092 34246
rect 12116 34244 12172 34246
rect 12196 34244 12252 34246
rect 16956 34298 17012 34300
rect 17036 34298 17092 34300
rect 17116 34298 17172 34300
rect 17196 34298 17252 34300
rect 16956 34246 17002 34298
rect 17002 34246 17012 34298
rect 17036 34246 17066 34298
rect 17066 34246 17078 34298
rect 17078 34246 17092 34298
rect 17116 34246 17130 34298
rect 17130 34246 17142 34298
rect 17142 34246 17172 34298
rect 17196 34246 17206 34298
rect 17206 34246 17252 34298
rect 16956 34244 17012 34246
rect 17036 34244 17092 34246
rect 17116 34244 17172 34246
rect 17196 34244 17252 34246
rect 21956 34298 22012 34300
rect 22036 34298 22092 34300
rect 22116 34298 22172 34300
rect 22196 34298 22252 34300
rect 21956 34246 22002 34298
rect 22002 34246 22012 34298
rect 22036 34246 22066 34298
rect 22066 34246 22078 34298
rect 22078 34246 22092 34298
rect 22116 34246 22130 34298
rect 22130 34246 22142 34298
rect 22142 34246 22172 34298
rect 22196 34246 22206 34298
rect 22206 34246 22252 34298
rect 21956 34244 22012 34246
rect 22036 34244 22092 34246
rect 22116 34244 22172 34246
rect 22196 34244 22252 34246
rect 26956 34298 27012 34300
rect 27036 34298 27092 34300
rect 27116 34298 27172 34300
rect 27196 34298 27252 34300
rect 26956 34246 27002 34298
rect 27002 34246 27012 34298
rect 27036 34246 27066 34298
rect 27066 34246 27078 34298
rect 27078 34246 27092 34298
rect 27116 34246 27130 34298
rect 27130 34246 27142 34298
rect 27142 34246 27172 34298
rect 27196 34246 27206 34298
rect 27206 34246 27252 34298
rect 26956 34244 27012 34246
rect 27036 34244 27092 34246
rect 27116 34244 27172 34246
rect 27196 34244 27252 34246
rect 31956 34298 32012 34300
rect 32036 34298 32092 34300
rect 32116 34298 32172 34300
rect 32196 34298 32252 34300
rect 31956 34246 32002 34298
rect 32002 34246 32012 34298
rect 32036 34246 32066 34298
rect 32066 34246 32078 34298
rect 32078 34246 32092 34298
rect 32116 34246 32130 34298
rect 32130 34246 32142 34298
rect 32142 34246 32172 34298
rect 32196 34246 32206 34298
rect 32206 34246 32252 34298
rect 31956 34244 32012 34246
rect 32036 34244 32092 34246
rect 32116 34244 32172 34246
rect 32196 34244 32252 34246
rect 36956 34298 37012 34300
rect 37036 34298 37092 34300
rect 37116 34298 37172 34300
rect 37196 34298 37252 34300
rect 36956 34246 37002 34298
rect 37002 34246 37012 34298
rect 37036 34246 37066 34298
rect 37066 34246 37078 34298
rect 37078 34246 37092 34298
rect 37116 34246 37130 34298
rect 37130 34246 37142 34298
rect 37142 34246 37172 34298
rect 37196 34246 37206 34298
rect 37206 34246 37252 34298
rect 36956 34244 37012 34246
rect 37036 34244 37092 34246
rect 37116 34244 37172 34246
rect 37196 34244 37252 34246
rect 41956 34298 42012 34300
rect 42036 34298 42092 34300
rect 42116 34298 42172 34300
rect 42196 34298 42252 34300
rect 41956 34246 42002 34298
rect 42002 34246 42012 34298
rect 42036 34246 42066 34298
rect 42066 34246 42078 34298
rect 42078 34246 42092 34298
rect 42116 34246 42130 34298
rect 42130 34246 42142 34298
rect 42142 34246 42172 34298
rect 42196 34246 42206 34298
rect 42206 34246 42252 34298
rect 41956 34244 42012 34246
rect 42036 34244 42092 34246
rect 42116 34244 42172 34246
rect 42196 34244 42252 34246
rect 46956 34298 47012 34300
rect 47036 34298 47092 34300
rect 47116 34298 47172 34300
rect 47196 34298 47252 34300
rect 46956 34246 47002 34298
rect 47002 34246 47012 34298
rect 47036 34246 47066 34298
rect 47066 34246 47078 34298
rect 47078 34246 47092 34298
rect 47116 34246 47130 34298
rect 47130 34246 47142 34298
rect 47142 34246 47172 34298
rect 47196 34246 47206 34298
rect 47206 34246 47252 34298
rect 46956 34244 47012 34246
rect 47036 34244 47092 34246
rect 47116 34244 47172 34246
rect 47196 34244 47252 34246
rect 51956 34298 52012 34300
rect 52036 34298 52092 34300
rect 52116 34298 52172 34300
rect 52196 34298 52252 34300
rect 51956 34246 52002 34298
rect 52002 34246 52012 34298
rect 52036 34246 52066 34298
rect 52066 34246 52078 34298
rect 52078 34246 52092 34298
rect 52116 34246 52130 34298
rect 52130 34246 52142 34298
rect 52142 34246 52172 34298
rect 52196 34246 52206 34298
rect 52206 34246 52252 34298
rect 51956 34244 52012 34246
rect 52036 34244 52092 34246
rect 52116 34244 52172 34246
rect 52196 34244 52252 34246
rect 56956 34298 57012 34300
rect 57036 34298 57092 34300
rect 57116 34298 57172 34300
rect 57196 34298 57252 34300
rect 56956 34246 57002 34298
rect 57002 34246 57012 34298
rect 57036 34246 57066 34298
rect 57066 34246 57078 34298
rect 57078 34246 57092 34298
rect 57116 34246 57130 34298
rect 57130 34246 57142 34298
rect 57142 34246 57172 34298
rect 57196 34246 57206 34298
rect 57206 34246 57252 34298
rect 56956 34244 57012 34246
rect 57036 34244 57092 34246
rect 57116 34244 57172 34246
rect 57196 34244 57252 34246
rect 2616 33754 2672 33756
rect 2696 33754 2752 33756
rect 2776 33754 2832 33756
rect 2856 33754 2912 33756
rect 2616 33702 2662 33754
rect 2662 33702 2672 33754
rect 2696 33702 2726 33754
rect 2726 33702 2738 33754
rect 2738 33702 2752 33754
rect 2776 33702 2790 33754
rect 2790 33702 2802 33754
rect 2802 33702 2832 33754
rect 2856 33702 2866 33754
rect 2866 33702 2912 33754
rect 2616 33700 2672 33702
rect 2696 33700 2752 33702
rect 2776 33700 2832 33702
rect 2856 33700 2912 33702
rect 7616 33754 7672 33756
rect 7696 33754 7752 33756
rect 7776 33754 7832 33756
rect 7856 33754 7912 33756
rect 7616 33702 7662 33754
rect 7662 33702 7672 33754
rect 7696 33702 7726 33754
rect 7726 33702 7738 33754
rect 7738 33702 7752 33754
rect 7776 33702 7790 33754
rect 7790 33702 7802 33754
rect 7802 33702 7832 33754
rect 7856 33702 7866 33754
rect 7866 33702 7912 33754
rect 7616 33700 7672 33702
rect 7696 33700 7752 33702
rect 7776 33700 7832 33702
rect 7856 33700 7912 33702
rect 12616 33754 12672 33756
rect 12696 33754 12752 33756
rect 12776 33754 12832 33756
rect 12856 33754 12912 33756
rect 12616 33702 12662 33754
rect 12662 33702 12672 33754
rect 12696 33702 12726 33754
rect 12726 33702 12738 33754
rect 12738 33702 12752 33754
rect 12776 33702 12790 33754
rect 12790 33702 12802 33754
rect 12802 33702 12832 33754
rect 12856 33702 12866 33754
rect 12866 33702 12912 33754
rect 12616 33700 12672 33702
rect 12696 33700 12752 33702
rect 12776 33700 12832 33702
rect 12856 33700 12912 33702
rect 17616 33754 17672 33756
rect 17696 33754 17752 33756
rect 17776 33754 17832 33756
rect 17856 33754 17912 33756
rect 17616 33702 17662 33754
rect 17662 33702 17672 33754
rect 17696 33702 17726 33754
rect 17726 33702 17738 33754
rect 17738 33702 17752 33754
rect 17776 33702 17790 33754
rect 17790 33702 17802 33754
rect 17802 33702 17832 33754
rect 17856 33702 17866 33754
rect 17866 33702 17912 33754
rect 17616 33700 17672 33702
rect 17696 33700 17752 33702
rect 17776 33700 17832 33702
rect 17856 33700 17912 33702
rect 22616 33754 22672 33756
rect 22696 33754 22752 33756
rect 22776 33754 22832 33756
rect 22856 33754 22912 33756
rect 22616 33702 22662 33754
rect 22662 33702 22672 33754
rect 22696 33702 22726 33754
rect 22726 33702 22738 33754
rect 22738 33702 22752 33754
rect 22776 33702 22790 33754
rect 22790 33702 22802 33754
rect 22802 33702 22832 33754
rect 22856 33702 22866 33754
rect 22866 33702 22912 33754
rect 22616 33700 22672 33702
rect 22696 33700 22752 33702
rect 22776 33700 22832 33702
rect 22856 33700 22912 33702
rect 27616 33754 27672 33756
rect 27696 33754 27752 33756
rect 27776 33754 27832 33756
rect 27856 33754 27912 33756
rect 27616 33702 27662 33754
rect 27662 33702 27672 33754
rect 27696 33702 27726 33754
rect 27726 33702 27738 33754
rect 27738 33702 27752 33754
rect 27776 33702 27790 33754
rect 27790 33702 27802 33754
rect 27802 33702 27832 33754
rect 27856 33702 27866 33754
rect 27866 33702 27912 33754
rect 27616 33700 27672 33702
rect 27696 33700 27752 33702
rect 27776 33700 27832 33702
rect 27856 33700 27912 33702
rect 32616 33754 32672 33756
rect 32696 33754 32752 33756
rect 32776 33754 32832 33756
rect 32856 33754 32912 33756
rect 32616 33702 32662 33754
rect 32662 33702 32672 33754
rect 32696 33702 32726 33754
rect 32726 33702 32738 33754
rect 32738 33702 32752 33754
rect 32776 33702 32790 33754
rect 32790 33702 32802 33754
rect 32802 33702 32832 33754
rect 32856 33702 32866 33754
rect 32866 33702 32912 33754
rect 32616 33700 32672 33702
rect 32696 33700 32752 33702
rect 32776 33700 32832 33702
rect 32856 33700 32912 33702
rect 37616 33754 37672 33756
rect 37696 33754 37752 33756
rect 37776 33754 37832 33756
rect 37856 33754 37912 33756
rect 37616 33702 37662 33754
rect 37662 33702 37672 33754
rect 37696 33702 37726 33754
rect 37726 33702 37738 33754
rect 37738 33702 37752 33754
rect 37776 33702 37790 33754
rect 37790 33702 37802 33754
rect 37802 33702 37832 33754
rect 37856 33702 37866 33754
rect 37866 33702 37912 33754
rect 37616 33700 37672 33702
rect 37696 33700 37752 33702
rect 37776 33700 37832 33702
rect 37856 33700 37912 33702
rect 42616 33754 42672 33756
rect 42696 33754 42752 33756
rect 42776 33754 42832 33756
rect 42856 33754 42912 33756
rect 42616 33702 42662 33754
rect 42662 33702 42672 33754
rect 42696 33702 42726 33754
rect 42726 33702 42738 33754
rect 42738 33702 42752 33754
rect 42776 33702 42790 33754
rect 42790 33702 42802 33754
rect 42802 33702 42832 33754
rect 42856 33702 42866 33754
rect 42866 33702 42912 33754
rect 42616 33700 42672 33702
rect 42696 33700 42752 33702
rect 42776 33700 42832 33702
rect 42856 33700 42912 33702
rect 47616 33754 47672 33756
rect 47696 33754 47752 33756
rect 47776 33754 47832 33756
rect 47856 33754 47912 33756
rect 47616 33702 47662 33754
rect 47662 33702 47672 33754
rect 47696 33702 47726 33754
rect 47726 33702 47738 33754
rect 47738 33702 47752 33754
rect 47776 33702 47790 33754
rect 47790 33702 47802 33754
rect 47802 33702 47832 33754
rect 47856 33702 47866 33754
rect 47866 33702 47912 33754
rect 47616 33700 47672 33702
rect 47696 33700 47752 33702
rect 47776 33700 47832 33702
rect 47856 33700 47912 33702
rect 52616 33754 52672 33756
rect 52696 33754 52752 33756
rect 52776 33754 52832 33756
rect 52856 33754 52912 33756
rect 52616 33702 52662 33754
rect 52662 33702 52672 33754
rect 52696 33702 52726 33754
rect 52726 33702 52738 33754
rect 52738 33702 52752 33754
rect 52776 33702 52790 33754
rect 52790 33702 52802 33754
rect 52802 33702 52832 33754
rect 52856 33702 52866 33754
rect 52866 33702 52912 33754
rect 52616 33700 52672 33702
rect 52696 33700 52752 33702
rect 52776 33700 52832 33702
rect 52856 33700 52912 33702
rect 57616 33754 57672 33756
rect 57696 33754 57752 33756
rect 57776 33754 57832 33756
rect 57856 33754 57912 33756
rect 57616 33702 57662 33754
rect 57662 33702 57672 33754
rect 57696 33702 57726 33754
rect 57726 33702 57738 33754
rect 57738 33702 57752 33754
rect 57776 33702 57790 33754
rect 57790 33702 57802 33754
rect 57802 33702 57832 33754
rect 57856 33702 57866 33754
rect 57866 33702 57912 33754
rect 57616 33700 57672 33702
rect 57696 33700 57752 33702
rect 57776 33700 57832 33702
rect 57856 33700 57912 33702
rect 58530 33496 58586 33552
rect 1956 33210 2012 33212
rect 2036 33210 2092 33212
rect 2116 33210 2172 33212
rect 2196 33210 2252 33212
rect 1956 33158 2002 33210
rect 2002 33158 2012 33210
rect 2036 33158 2066 33210
rect 2066 33158 2078 33210
rect 2078 33158 2092 33210
rect 2116 33158 2130 33210
rect 2130 33158 2142 33210
rect 2142 33158 2172 33210
rect 2196 33158 2206 33210
rect 2206 33158 2252 33210
rect 1956 33156 2012 33158
rect 2036 33156 2092 33158
rect 2116 33156 2172 33158
rect 2196 33156 2252 33158
rect 6956 33210 7012 33212
rect 7036 33210 7092 33212
rect 7116 33210 7172 33212
rect 7196 33210 7252 33212
rect 6956 33158 7002 33210
rect 7002 33158 7012 33210
rect 7036 33158 7066 33210
rect 7066 33158 7078 33210
rect 7078 33158 7092 33210
rect 7116 33158 7130 33210
rect 7130 33158 7142 33210
rect 7142 33158 7172 33210
rect 7196 33158 7206 33210
rect 7206 33158 7252 33210
rect 6956 33156 7012 33158
rect 7036 33156 7092 33158
rect 7116 33156 7172 33158
rect 7196 33156 7252 33158
rect 11956 33210 12012 33212
rect 12036 33210 12092 33212
rect 12116 33210 12172 33212
rect 12196 33210 12252 33212
rect 11956 33158 12002 33210
rect 12002 33158 12012 33210
rect 12036 33158 12066 33210
rect 12066 33158 12078 33210
rect 12078 33158 12092 33210
rect 12116 33158 12130 33210
rect 12130 33158 12142 33210
rect 12142 33158 12172 33210
rect 12196 33158 12206 33210
rect 12206 33158 12252 33210
rect 11956 33156 12012 33158
rect 12036 33156 12092 33158
rect 12116 33156 12172 33158
rect 12196 33156 12252 33158
rect 16956 33210 17012 33212
rect 17036 33210 17092 33212
rect 17116 33210 17172 33212
rect 17196 33210 17252 33212
rect 16956 33158 17002 33210
rect 17002 33158 17012 33210
rect 17036 33158 17066 33210
rect 17066 33158 17078 33210
rect 17078 33158 17092 33210
rect 17116 33158 17130 33210
rect 17130 33158 17142 33210
rect 17142 33158 17172 33210
rect 17196 33158 17206 33210
rect 17206 33158 17252 33210
rect 16956 33156 17012 33158
rect 17036 33156 17092 33158
rect 17116 33156 17172 33158
rect 17196 33156 17252 33158
rect 21956 33210 22012 33212
rect 22036 33210 22092 33212
rect 22116 33210 22172 33212
rect 22196 33210 22252 33212
rect 21956 33158 22002 33210
rect 22002 33158 22012 33210
rect 22036 33158 22066 33210
rect 22066 33158 22078 33210
rect 22078 33158 22092 33210
rect 22116 33158 22130 33210
rect 22130 33158 22142 33210
rect 22142 33158 22172 33210
rect 22196 33158 22206 33210
rect 22206 33158 22252 33210
rect 21956 33156 22012 33158
rect 22036 33156 22092 33158
rect 22116 33156 22172 33158
rect 22196 33156 22252 33158
rect 26956 33210 27012 33212
rect 27036 33210 27092 33212
rect 27116 33210 27172 33212
rect 27196 33210 27252 33212
rect 26956 33158 27002 33210
rect 27002 33158 27012 33210
rect 27036 33158 27066 33210
rect 27066 33158 27078 33210
rect 27078 33158 27092 33210
rect 27116 33158 27130 33210
rect 27130 33158 27142 33210
rect 27142 33158 27172 33210
rect 27196 33158 27206 33210
rect 27206 33158 27252 33210
rect 26956 33156 27012 33158
rect 27036 33156 27092 33158
rect 27116 33156 27172 33158
rect 27196 33156 27252 33158
rect 31956 33210 32012 33212
rect 32036 33210 32092 33212
rect 32116 33210 32172 33212
rect 32196 33210 32252 33212
rect 31956 33158 32002 33210
rect 32002 33158 32012 33210
rect 32036 33158 32066 33210
rect 32066 33158 32078 33210
rect 32078 33158 32092 33210
rect 32116 33158 32130 33210
rect 32130 33158 32142 33210
rect 32142 33158 32172 33210
rect 32196 33158 32206 33210
rect 32206 33158 32252 33210
rect 31956 33156 32012 33158
rect 32036 33156 32092 33158
rect 32116 33156 32172 33158
rect 32196 33156 32252 33158
rect 36956 33210 37012 33212
rect 37036 33210 37092 33212
rect 37116 33210 37172 33212
rect 37196 33210 37252 33212
rect 36956 33158 37002 33210
rect 37002 33158 37012 33210
rect 37036 33158 37066 33210
rect 37066 33158 37078 33210
rect 37078 33158 37092 33210
rect 37116 33158 37130 33210
rect 37130 33158 37142 33210
rect 37142 33158 37172 33210
rect 37196 33158 37206 33210
rect 37206 33158 37252 33210
rect 36956 33156 37012 33158
rect 37036 33156 37092 33158
rect 37116 33156 37172 33158
rect 37196 33156 37252 33158
rect 41956 33210 42012 33212
rect 42036 33210 42092 33212
rect 42116 33210 42172 33212
rect 42196 33210 42252 33212
rect 41956 33158 42002 33210
rect 42002 33158 42012 33210
rect 42036 33158 42066 33210
rect 42066 33158 42078 33210
rect 42078 33158 42092 33210
rect 42116 33158 42130 33210
rect 42130 33158 42142 33210
rect 42142 33158 42172 33210
rect 42196 33158 42206 33210
rect 42206 33158 42252 33210
rect 41956 33156 42012 33158
rect 42036 33156 42092 33158
rect 42116 33156 42172 33158
rect 42196 33156 42252 33158
rect 46956 33210 47012 33212
rect 47036 33210 47092 33212
rect 47116 33210 47172 33212
rect 47196 33210 47252 33212
rect 46956 33158 47002 33210
rect 47002 33158 47012 33210
rect 47036 33158 47066 33210
rect 47066 33158 47078 33210
rect 47078 33158 47092 33210
rect 47116 33158 47130 33210
rect 47130 33158 47142 33210
rect 47142 33158 47172 33210
rect 47196 33158 47206 33210
rect 47206 33158 47252 33210
rect 46956 33156 47012 33158
rect 47036 33156 47092 33158
rect 47116 33156 47172 33158
rect 47196 33156 47252 33158
rect 51956 33210 52012 33212
rect 52036 33210 52092 33212
rect 52116 33210 52172 33212
rect 52196 33210 52252 33212
rect 51956 33158 52002 33210
rect 52002 33158 52012 33210
rect 52036 33158 52066 33210
rect 52066 33158 52078 33210
rect 52078 33158 52092 33210
rect 52116 33158 52130 33210
rect 52130 33158 52142 33210
rect 52142 33158 52172 33210
rect 52196 33158 52206 33210
rect 52206 33158 52252 33210
rect 51956 33156 52012 33158
rect 52036 33156 52092 33158
rect 52116 33156 52172 33158
rect 52196 33156 52252 33158
rect 56956 33210 57012 33212
rect 57036 33210 57092 33212
rect 57116 33210 57172 33212
rect 57196 33210 57252 33212
rect 56956 33158 57002 33210
rect 57002 33158 57012 33210
rect 57036 33158 57066 33210
rect 57066 33158 57078 33210
rect 57078 33158 57092 33210
rect 57116 33158 57130 33210
rect 57130 33158 57142 33210
rect 57142 33158 57172 33210
rect 57196 33158 57206 33210
rect 57206 33158 57252 33210
rect 56956 33156 57012 33158
rect 57036 33156 57092 33158
rect 57116 33156 57172 33158
rect 57196 33156 57252 33158
rect 58530 32680 58586 32736
rect 2616 32666 2672 32668
rect 2696 32666 2752 32668
rect 2776 32666 2832 32668
rect 2856 32666 2912 32668
rect 2616 32614 2662 32666
rect 2662 32614 2672 32666
rect 2696 32614 2726 32666
rect 2726 32614 2738 32666
rect 2738 32614 2752 32666
rect 2776 32614 2790 32666
rect 2790 32614 2802 32666
rect 2802 32614 2832 32666
rect 2856 32614 2866 32666
rect 2866 32614 2912 32666
rect 2616 32612 2672 32614
rect 2696 32612 2752 32614
rect 2776 32612 2832 32614
rect 2856 32612 2912 32614
rect 7616 32666 7672 32668
rect 7696 32666 7752 32668
rect 7776 32666 7832 32668
rect 7856 32666 7912 32668
rect 7616 32614 7662 32666
rect 7662 32614 7672 32666
rect 7696 32614 7726 32666
rect 7726 32614 7738 32666
rect 7738 32614 7752 32666
rect 7776 32614 7790 32666
rect 7790 32614 7802 32666
rect 7802 32614 7832 32666
rect 7856 32614 7866 32666
rect 7866 32614 7912 32666
rect 7616 32612 7672 32614
rect 7696 32612 7752 32614
rect 7776 32612 7832 32614
rect 7856 32612 7912 32614
rect 12616 32666 12672 32668
rect 12696 32666 12752 32668
rect 12776 32666 12832 32668
rect 12856 32666 12912 32668
rect 12616 32614 12662 32666
rect 12662 32614 12672 32666
rect 12696 32614 12726 32666
rect 12726 32614 12738 32666
rect 12738 32614 12752 32666
rect 12776 32614 12790 32666
rect 12790 32614 12802 32666
rect 12802 32614 12832 32666
rect 12856 32614 12866 32666
rect 12866 32614 12912 32666
rect 12616 32612 12672 32614
rect 12696 32612 12752 32614
rect 12776 32612 12832 32614
rect 12856 32612 12912 32614
rect 17616 32666 17672 32668
rect 17696 32666 17752 32668
rect 17776 32666 17832 32668
rect 17856 32666 17912 32668
rect 17616 32614 17662 32666
rect 17662 32614 17672 32666
rect 17696 32614 17726 32666
rect 17726 32614 17738 32666
rect 17738 32614 17752 32666
rect 17776 32614 17790 32666
rect 17790 32614 17802 32666
rect 17802 32614 17832 32666
rect 17856 32614 17866 32666
rect 17866 32614 17912 32666
rect 17616 32612 17672 32614
rect 17696 32612 17752 32614
rect 17776 32612 17832 32614
rect 17856 32612 17912 32614
rect 22616 32666 22672 32668
rect 22696 32666 22752 32668
rect 22776 32666 22832 32668
rect 22856 32666 22912 32668
rect 22616 32614 22662 32666
rect 22662 32614 22672 32666
rect 22696 32614 22726 32666
rect 22726 32614 22738 32666
rect 22738 32614 22752 32666
rect 22776 32614 22790 32666
rect 22790 32614 22802 32666
rect 22802 32614 22832 32666
rect 22856 32614 22866 32666
rect 22866 32614 22912 32666
rect 22616 32612 22672 32614
rect 22696 32612 22752 32614
rect 22776 32612 22832 32614
rect 22856 32612 22912 32614
rect 27616 32666 27672 32668
rect 27696 32666 27752 32668
rect 27776 32666 27832 32668
rect 27856 32666 27912 32668
rect 27616 32614 27662 32666
rect 27662 32614 27672 32666
rect 27696 32614 27726 32666
rect 27726 32614 27738 32666
rect 27738 32614 27752 32666
rect 27776 32614 27790 32666
rect 27790 32614 27802 32666
rect 27802 32614 27832 32666
rect 27856 32614 27866 32666
rect 27866 32614 27912 32666
rect 27616 32612 27672 32614
rect 27696 32612 27752 32614
rect 27776 32612 27832 32614
rect 27856 32612 27912 32614
rect 32616 32666 32672 32668
rect 32696 32666 32752 32668
rect 32776 32666 32832 32668
rect 32856 32666 32912 32668
rect 32616 32614 32662 32666
rect 32662 32614 32672 32666
rect 32696 32614 32726 32666
rect 32726 32614 32738 32666
rect 32738 32614 32752 32666
rect 32776 32614 32790 32666
rect 32790 32614 32802 32666
rect 32802 32614 32832 32666
rect 32856 32614 32866 32666
rect 32866 32614 32912 32666
rect 32616 32612 32672 32614
rect 32696 32612 32752 32614
rect 32776 32612 32832 32614
rect 32856 32612 32912 32614
rect 37616 32666 37672 32668
rect 37696 32666 37752 32668
rect 37776 32666 37832 32668
rect 37856 32666 37912 32668
rect 37616 32614 37662 32666
rect 37662 32614 37672 32666
rect 37696 32614 37726 32666
rect 37726 32614 37738 32666
rect 37738 32614 37752 32666
rect 37776 32614 37790 32666
rect 37790 32614 37802 32666
rect 37802 32614 37832 32666
rect 37856 32614 37866 32666
rect 37866 32614 37912 32666
rect 37616 32612 37672 32614
rect 37696 32612 37752 32614
rect 37776 32612 37832 32614
rect 37856 32612 37912 32614
rect 42616 32666 42672 32668
rect 42696 32666 42752 32668
rect 42776 32666 42832 32668
rect 42856 32666 42912 32668
rect 42616 32614 42662 32666
rect 42662 32614 42672 32666
rect 42696 32614 42726 32666
rect 42726 32614 42738 32666
rect 42738 32614 42752 32666
rect 42776 32614 42790 32666
rect 42790 32614 42802 32666
rect 42802 32614 42832 32666
rect 42856 32614 42866 32666
rect 42866 32614 42912 32666
rect 42616 32612 42672 32614
rect 42696 32612 42752 32614
rect 42776 32612 42832 32614
rect 42856 32612 42912 32614
rect 47616 32666 47672 32668
rect 47696 32666 47752 32668
rect 47776 32666 47832 32668
rect 47856 32666 47912 32668
rect 47616 32614 47662 32666
rect 47662 32614 47672 32666
rect 47696 32614 47726 32666
rect 47726 32614 47738 32666
rect 47738 32614 47752 32666
rect 47776 32614 47790 32666
rect 47790 32614 47802 32666
rect 47802 32614 47832 32666
rect 47856 32614 47866 32666
rect 47866 32614 47912 32666
rect 47616 32612 47672 32614
rect 47696 32612 47752 32614
rect 47776 32612 47832 32614
rect 47856 32612 47912 32614
rect 52616 32666 52672 32668
rect 52696 32666 52752 32668
rect 52776 32666 52832 32668
rect 52856 32666 52912 32668
rect 52616 32614 52662 32666
rect 52662 32614 52672 32666
rect 52696 32614 52726 32666
rect 52726 32614 52738 32666
rect 52738 32614 52752 32666
rect 52776 32614 52790 32666
rect 52790 32614 52802 32666
rect 52802 32614 52832 32666
rect 52856 32614 52866 32666
rect 52866 32614 52912 32666
rect 52616 32612 52672 32614
rect 52696 32612 52752 32614
rect 52776 32612 52832 32614
rect 52856 32612 52912 32614
rect 57616 32666 57672 32668
rect 57696 32666 57752 32668
rect 57776 32666 57832 32668
rect 57856 32666 57912 32668
rect 57616 32614 57662 32666
rect 57662 32614 57672 32666
rect 57696 32614 57726 32666
rect 57726 32614 57738 32666
rect 57738 32614 57752 32666
rect 57776 32614 57790 32666
rect 57790 32614 57802 32666
rect 57802 32614 57832 32666
rect 57856 32614 57866 32666
rect 57866 32614 57912 32666
rect 57616 32612 57672 32614
rect 57696 32612 57752 32614
rect 57776 32612 57832 32614
rect 57856 32612 57912 32614
rect 1956 32122 2012 32124
rect 2036 32122 2092 32124
rect 2116 32122 2172 32124
rect 2196 32122 2252 32124
rect 1956 32070 2002 32122
rect 2002 32070 2012 32122
rect 2036 32070 2066 32122
rect 2066 32070 2078 32122
rect 2078 32070 2092 32122
rect 2116 32070 2130 32122
rect 2130 32070 2142 32122
rect 2142 32070 2172 32122
rect 2196 32070 2206 32122
rect 2206 32070 2252 32122
rect 1956 32068 2012 32070
rect 2036 32068 2092 32070
rect 2116 32068 2172 32070
rect 2196 32068 2252 32070
rect 6956 32122 7012 32124
rect 7036 32122 7092 32124
rect 7116 32122 7172 32124
rect 7196 32122 7252 32124
rect 6956 32070 7002 32122
rect 7002 32070 7012 32122
rect 7036 32070 7066 32122
rect 7066 32070 7078 32122
rect 7078 32070 7092 32122
rect 7116 32070 7130 32122
rect 7130 32070 7142 32122
rect 7142 32070 7172 32122
rect 7196 32070 7206 32122
rect 7206 32070 7252 32122
rect 6956 32068 7012 32070
rect 7036 32068 7092 32070
rect 7116 32068 7172 32070
rect 7196 32068 7252 32070
rect 11956 32122 12012 32124
rect 12036 32122 12092 32124
rect 12116 32122 12172 32124
rect 12196 32122 12252 32124
rect 11956 32070 12002 32122
rect 12002 32070 12012 32122
rect 12036 32070 12066 32122
rect 12066 32070 12078 32122
rect 12078 32070 12092 32122
rect 12116 32070 12130 32122
rect 12130 32070 12142 32122
rect 12142 32070 12172 32122
rect 12196 32070 12206 32122
rect 12206 32070 12252 32122
rect 11956 32068 12012 32070
rect 12036 32068 12092 32070
rect 12116 32068 12172 32070
rect 12196 32068 12252 32070
rect 16956 32122 17012 32124
rect 17036 32122 17092 32124
rect 17116 32122 17172 32124
rect 17196 32122 17252 32124
rect 16956 32070 17002 32122
rect 17002 32070 17012 32122
rect 17036 32070 17066 32122
rect 17066 32070 17078 32122
rect 17078 32070 17092 32122
rect 17116 32070 17130 32122
rect 17130 32070 17142 32122
rect 17142 32070 17172 32122
rect 17196 32070 17206 32122
rect 17206 32070 17252 32122
rect 16956 32068 17012 32070
rect 17036 32068 17092 32070
rect 17116 32068 17172 32070
rect 17196 32068 17252 32070
rect 21956 32122 22012 32124
rect 22036 32122 22092 32124
rect 22116 32122 22172 32124
rect 22196 32122 22252 32124
rect 21956 32070 22002 32122
rect 22002 32070 22012 32122
rect 22036 32070 22066 32122
rect 22066 32070 22078 32122
rect 22078 32070 22092 32122
rect 22116 32070 22130 32122
rect 22130 32070 22142 32122
rect 22142 32070 22172 32122
rect 22196 32070 22206 32122
rect 22206 32070 22252 32122
rect 21956 32068 22012 32070
rect 22036 32068 22092 32070
rect 22116 32068 22172 32070
rect 22196 32068 22252 32070
rect 26956 32122 27012 32124
rect 27036 32122 27092 32124
rect 27116 32122 27172 32124
rect 27196 32122 27252 32124
rect 26956 32070 27002 32122
rect 27002 32070 27012 32122
rect 27036 32070 27066 32122
rect 27066 32070 27078 32122
rect 27078 32070 27092 32122
rect 27116 32070 27130 32122
rect 27130 32070 27142 32122
rect 27142 32070 27172 32122
rect 27196 32070 27206 32122
rect 27206 32070 27252 32122
rect 26956 32068 27012 32070
rect 27036 32068 27092 32070
rect 27116 32068 27172 32070
rect 27196 32068 27252 32070
rect 31956 32122 32012 32124
rect 32036 32122 32092 32124
rect 32116 32122 32172 32124
rect 32196 32122 32252 32124
rect 31956 32070 32002 32122
rect 32002 32070 32012 32122
rect 32036 32070 32066 32122
rect 32066 32070 32078 32122
rect 32078 32070 32092 32122
rect 32116 32070 32130 32122
rect 32130 32070 32142 32122
rect 32142 32070 32172 32122
rect 32196 32070 32206 32122
rect 32206 32070 32252 32122
rect 31956 32068 32012 32070
rect 32036 32068 32092 32070
rect 32116 32068 32172 32070
rect 32196 32068 32252 32070
rect 36956 32122 37012 32124
rect 37036 32122 37092 32124
rect 37116 32122 37172 32124
rect 37196 32122 37252 32124
rect 36956 32070 37002 32122
rect 37002 32070 37012 32122
rect 37036 32070 37066 32122
rect 37066 32070 37078 32122
rect 37078 32070 37092 32122
rect 37116 32070 37130 32122
rect 37130 32070 37142 32122
rect 37142 32070 37172 32122
rect 37196 32070 37206 32122
rect 37206 32070 37252 32122
rect 36956 32068 37012 32070
rect 37036 32068 37092 32070
rect 37116 32068 37172 32070
rect 37196 32068 37252 32070
rect 41956 32122 42012 32124
rect 42036 32122 42092 32124
rect 42116 32122 42172 32124
rect 42196 32122 42252 32124
rect 41956 32070 42002 32122
rect 42002 32070 42012 32122
rect 42036 32070 42066 32122
rect 42066 32070 42078 32122
rect 42078 32070 42092 32122
rect 42116 32070 42130 32122
rect 42130 32070 42142 32122
rect 42142 32070 42172 32122
rect 42196 32070 42206 32122
rect 42206 32070 42252 32122
rect 41956 32068 42012 32070
rect 42036 32068 42092 32070
rect 42116 32068 42172 32070
rect 42196 32068 42252 32070
rect 46956 32122 47012 32124
rect 47036 32122 47092 32124
rect 47116 32122 47172 32124
rect 47196 32122 47252 32124
rect 46956 32070 47002 32122
rect 47002 32070 47012 32122
rect 47036 32070 47066 32122
rect 47066 32070 47078 32122
rect 47078 32070 47092 32122
rect 47116 32070 47130 32122
rect 47130 32070 47142 32122
rect 47142 32070 47172 32122
rect 47196 32070 47206 32122
rect 47206 32070 47252 32122
rect 46956 32068 47012 32070
rect 47036 32068 47092 32070
rect 47116 32068 47172 32070
rect 47196 32068 47252 32070
rect 51956 32122 52012 32124
rect 52036 32122 52092 32124
rect 52116 32122 52172 32124
rect 52196 32122 52252 32124
rect 51956 32070 52002 32122
rect 52002 32070 52012 32122
rect 52036 32070 52066 32122
rect 52066 32070 52078 32122
rect 52078 32070 52092 32122
rect 52116 32070 52130 32122
rect 52130 32070 52142 32122
rect 52142 32070 52172 32122
rect 52196 32070 52206 32122
rect 52206 32070 52252 32122
rect 51956 32068 52012 32070
rect 52036 32068 52092 32070
rect 52116 32068 52172 32070
rect 52196 32068 52252 32070
rect 56956 32122 57012 32124
rect 57036 32122 57092 32124
rect 57116 32122 57172 32124
rect 57196 32122 57252 32124
rect 56956 32070 57002 32122
rect 57002 32070 57012 32122
rect 57036 32070 57066 32122
rect 57066 32070 57078 32122
rect 57078 32070 57092 32122
rect 57116 32070 57130 32122
rect 57130 32070 57142 32122
rect 57142 32070 57172 32122
rect 57196 32070 57206 32122
rect 57206 32070 57252 32122
rect 56956 32068 57012 32070
rect 57036 32068 57092 32070
rect 57116 32068 57172 32070
rect 57196 32068 57252 32070
rect 58530 31864 58586 31920
rect 2616 31578 2672 31580
rect 2696 31578 2752 31580
rect 2776 31578 2832 31580
rect 2856 31578 2912 31580
rect 2616 31526 2662 31578
rect 2662 31526 2672 31578
rect 2696 31526 2726 31578
rect 2726 31526 2738 31578
rect 2738 31526 2752 31578
rect 2776 31526 2790 31578
rect 2790 31526 2802 31578
rect 2802 31526 2832 31578
rect 2856 31526 2866 31578
rect 2866 31526 2912 31578
rect 2616 31524 2672 31526
rect 2696 31524 2752 31526
rect 2776 31524 2832 31526
rect 2856 31524 2912 31526
rect 7616 31578 7672 31580
rect 7696 31578 7752 31580
rect 7776 31578 7832 31580
rect 7856 31578 7912 31580
rect 7616 31526 7662 31578
rect 7662 31526 7672 31578
rect 7696 31526 7726 31578
rect 7726 31526 7738 31578
rect 7738 31526 7752 31578
rect 7776 31526 7790 31578
rect 7790 31526 7802 31578
rect 7802 31526 7832 31578
rect 7856 31526 7866 31578
rect 7866 31526 7912 31578
rect 7616 31524 7672 31526
rect 7696 31524 7752 31526
rect 7776 31524 7832 31526
rect 7856 31524 7912 31526
rect 12616 31578 12672 31580
rect 12696 31578 12752 31580
rect 12776 31578 12832 31580
rect 12856 31578 12912 31580
rect 12616 31526 12662 31578
rect 12662 31526 12672 31578
rect 12696 31526 12726 31578
rect 12726 31526 12738 31578
rect 12738 31526 12752 31578
rect 12776 31526 12790 31578
rect 12790 31526 12802 31578
rect 12802 31526 12832 31578
rect 12856 31526 12866 31578
rect 12866 31526 12912 31578
rect 12616 31524 12672 31526
rect 12696 31524 12752 31526
rect 12776 31524 12832 31526
rect 12856 31524 12912 31526
rect 17616 31578 17672 31580
rect 17696 31578 17752 31580
rect 17776 31578 17832 31580
rect 17856 31578 17912 31580
rect 17616 31526 17662 31578
rect 17662 31526 17672 31578
rect 17696 31526 17726 31578
rect 17726 31526 17738 31578
rect 17738 31526 17752 31578
rect 17776 31526 17790 31578
rect 17790 31526 17802 31578
rect 17802 31526 17832 31578
rect 17856 31526 17866 31578
rect 17866 31526 17912 31578
rect 17616 31524 17672 31526
rect 17696 31524 17752 31526
rect 17776 31524 17832 31526
rect 17856 31524 17912 31526
rect 22616 31578 22672 31580
rect 22696 31578 22752 31580
rect 22776 31578 22832 31580
rect 22856 31578 22912 31580
rect 22616 31526 22662 31578
rect 22662 31526 22672 31578
rect 22696 31526 22726 31578
rect 22726 31526 22738 31578
rect 22738 31526 22752 31578
rect 22776 31526 22790 31578
rect 22790 31526 22802 31578
rect 22802 31526 22832 31578
rect 22856 31526 22866 31578
rect 22866 31526 22912 31578
rect 22616 31524 22672 31526
rect 22696 31524 22752 31526
rect 22776 31524 22832 31526
rect 22856 31524 22912 31526
rect 27616 31578 27672 31580
rect 27696 31578 27752 31580
rect 27776 31578 27832 31580
rect 27856 31578 27912 31580
rect 27616 31526 27662 31578
rect 27662 31526 27672 31578
rect 27696 31526 27726 31578
rect 27726 31526 27738 31578
rect 27738 31526 27752 31578
rect 27776 31526 27790 31578
rect 27790 31526 27802 31578
rect 27802 31526 27832 31578
rect 27856 31526 27866 31578
rect 27866 31526 27912 31578
rect 27616 31524 27672 31526
rect 27696 31524 27752 31526
rect 27776 31524 27832 31526
rect 27856 31524 27912 31526
rect 32616 31578 32672 31580
rect 32696 31578 32752 31580
rect 32776 31578 32832 31580
rect 32856 31578 32912 31580
rect 32616 31526 32662 31578
rect 32662 31526 32672 31578
rect 32696 31526 32726 31578
rect 32726 31526 32738 31578
rect 32738 31526 32752 31578
rect 32776 31526 32790 31578
rect 32790 31526 32802 31578
rect 32802 31526 32832 31578
rect 32856 31526 32866 31578
rect 32866 31526 32912 31578
rect 32616 31524 32672 31526
rect 32696 31524 32752 31526
rect 32776 31524 32832 31526
rect 32856 31524 32912 31526
rect 37616 31578 37672 31580
rect 37696 31578 37752 31580
rect 37776 31578 37832 31580
rect 37856 31578 37912 31580
rect 37616 31526 37662 31578
rect 37662 31526 37672 31578
rect 37696 31526 37726 31578
rect 37726 31526 37738 31578
rect 37738 31526 37752 31578
rect 37776 31526 37790 31578
rect 37790 31526 37802 31578
rect 37802 31526 37832 31578
rect 37856 31526 37866 31578
rect 37866 31526 37912 31578
rect 37616 31524 37672 31526
rect 37696 31524 37752 31526
rect 37776 31524 37832 31526
rect 37856 31524 37912 31526
rect 42616 31578 42672 31580
rect 42696 31578 42752 31580
rect 42776 31578 42832 31580
rect 42856 31578 42912 31580
rect 42616 31526 42662 31578
rect 42662 31526 42672 31578
rect 42696 31526 42726 31578
rect 42726 31526 42738 31578
rect 42738 31526 42752 31578
rect 42776 31526 42790 31578
rect 42790 31526 42802 31578
rect 42802 31526 42832 31578
rect 42856 31526 42866 31578
rect 42866 31526 42912 31578
rect 42616 31524 42672 31526
rect 42696 31524 42752 31526
rect 42776 31524 42832 31526
rect 42856 31524 42912 31526
rect 47616 31578 47672 31580
rect 47696 31578 47752 31580
rect 47776 31578 47832 31580
rect 47856 31578 47912 31580
rect 47616 31526 47662 31578
rect 47662 31526 47672 31578
rect 47696 31526 47726 31578
rect 47726 31526 47738 31578
rect 47738 31526 47752 31578
rect 47776 31526 47790 31578
rect 47790 31526 47802 31578
rect 47802 31526 47832 31578
rect 47856 31526 47866 31578
rect 47866 31526 47912 31578
rect 47616 31524 47672 31526
rect 47696 31524 47752 31526
rect 47776 31524 47832 31526
rect 47856 31524 47912 31526
rect 52616 31578 52672 31580
rect 52696 31578 52752 31580
rect 52776 31578 52832 31580
rect 52856 31578 52912 31580
rect 52616 31526 52662 31578
rect 52662 31526 52672 31578
rect 52696 31526 52726 31578
rect 52726 31526 52738 31578
rect 52738 31526 52752 31578
rect 52776 31526 52790 31578
rect 52790 31526 52802 31578
rect 52802 31526 52832 31578
rect 52856 31526 52866 31578
rect 52866 31526 52912 31578
rect 52616 31524 52672 31526
rect 52696 31524 52752 31526
rect 52776 31524 52832 31526
rect 52856 31524 52912 31526
rect 57616 31578 57672 31580
rect 57696 31578 57752 31580
rect 57776 31578 57832 31580
rect 57856 31578 57912 31580
rect 57616 31526 57662 31578
rect 57662 31526 57672 31578
rect 57696 31526 57726 31578
rect 57726 31526 57738 31578
rect 57738 31526 57752 31578
rect 57776 31526 57790 31578
rect 57790 31526 57802 31578
rect 57802 31526 57832 31578
rect 57856 31526 57866 31578
rect 57866 31526 57912 31578
rect 57616 31524 57672 31526
rect 57696 31524 57752 31526
rect 57776 31524 57832 31526
rect 57856 31524 57912 31526
rect 58530 31084 58532 31104
rect 58532 31084 58584 31104
rect 58584 31084 58586 31104
rect 58530 31048 58586 31084
rect 1956 31034 2012 31036
rect 2036 31034 2092 31036
rect 2116 31034 2172 31036
rect 2196 31034 2252 31036
rect 1956 30982 2002 31034
rect 2002 30982 2012 31034
rect 2036 30982 2066 31034
rect 2066 30982 2078 31034
rect 2078 30982 2092 31034
rect 2116 30982 2130 31034
rect 2130 30982 2142 31034
rect 2142 30982 2172 31034
rect 2196 30982 2206 31034
rect 2206 30982 2252 31034
rect 1956 30980 2012 30982
rect 2036 30980 2092 30982
rect 2116 30980 2172 30982
rect 2196 30980 2252 30982
rect 6956 31034 7012 31036
rect 7036 31034 7092 31036
rect 7116 31034 7172 31036
rect 7196 31034 7252 31036
rect 6956 30982 7002 31034
rect 7002 30982 7012 31034
rect 7036 30982 7066 31034
rect 7066 30982 7078 31034
rect 7078 30982 7092 31034
rect 7116 30982 7130 31034
rect 7130 30982 7142 31034
rect 7142 30982 7172 31034
rect 7196 30982 7206 31034
rect 7206 30982 7252 31034
rect 6956 30980 7012 30982
rect 7036 30980 7092 30982
rect 7116 30980 7172 30982
rect 7196 30980 7252 30982
rect 11956 31034 12012 31036
rect 12036 31034 12092 31036
rect 12116 31034 12172 31036
rect 12196 31034 12252 31036
rect 11956 30982 12002 31034
rect 12002 30982 12012 31034
rect 12036 30982 12066 31034
rect 12066 30982 12078 31034
rect 12078 30982 12092 31034
rect 12116 30982 12130 31034
rect 12130 30982 12142 31034
rect 12142 30982 12172 31034
rect 12196 30982 12206 31034
rect 12206 30982 12252 31034
rect 11956 30980 12012 30982
rect 12036 30980 12092 30982
rect 12116 30980 12172 30982
rect 12196 30980 12252 30982
rect 16956 31034 17012 31036
rect 17036 31034 17092 31036
rect 17116 31034 17172 31036
rect 17196 31034 17252 31036
rect 16956 30982 17002 31034
rect 17002 30982 17012 31034
rect 17036 30982 17066 31034
rect 17066 30982 17078 31034
rect 17078 30982 17092 31034
rect 17116 30982 17130 31034
rect 17130 30982 17142 31034
rect 17142 30982 17172 31034
rect 17196 30982 17206 31034
rect 17206 30982 17252 31034
rect 16956 30980 17012 30982
rect 17036 30980 17092 30982
rect 17116 30980 17172 30982
rect 17196 30980 17252 30982
rect 21956 31034 22012 31036
rect 22036 31034 22092 31036
rect 22116 31034 22172 31036
rect 22196 31034 22252 31036
rect 21956 30982 22002 31034
rect 22002 30982 22012 31034
rect 22036 30982 22066 31034
rect 22066 30982 22078 31034
rect 22078 30982 22092 31034
rect 22116 30982 22130 31034
rect 22130 30982 22142 31034
rect 22142 30982 22172 31034
rect 22196 30982 22206 31034
rect 22206 30982 22252 31034
rect 21956 30980 22012 30982
rect 22036 30980 22092 30982
rect 22116 30980 22172 30982
rect 22196 30980 22252 30982
rect 26956 31034 27012 31036
rect 27036 31034 27092 31036
rect 27116 31034 27172 31036
rect 27196 31034 27252 31036
rect 26956 30982 27002 31034
rect 27002 30982 27012 31034
rect 27036 30982 27066 31034
rect 27066 30982 27078 31034
rect 27078 30982 27092 31034
rect 27116 30982 27130 31034
rect 27130 30982 27142 31034
rect 27142 30982 27172 31034
rect 27196 30982 27206 31034
rect 27206 30982 27252 31034
rect 26956 30980 27012 30982
rect 27036 30980 27092 30982
rect 27116 30980 27172 30982
rect 27196 30980 27252 30982
rect 31956 31034 32012 31036
rect 32036 31034 32092 31036
rect 32116 31034 32172 31036
rect 32196 31034 32252 31036
rect 31956 30982 32002 31034
rect 32002 30982 32012 31034
rect 32036 30982 32066 31034
rect 32066 30982 32078 31034
rect 32078 30982 32092 31034
rect 32116 30982 32130 31034
rect 32130 30982 32142 31034
rect 32142 30982 32172 31034
rect 32196 30982 32206 31034
rect 32206 30982 32252 31034
rect 31956 30980 32012 30982
rect 32036 30980 32092 30982
rect 32116 30980 32172 30982
rect 32196 30980 32252 30982
rect 36956 31034 37012 31036
rect 37036 31034 37092 31036
rect 37116 31034 37172 31036
rect 37196 31034 37252 31036
rect 36956 30982 37002 31034
rect 37002 30982 37012 31034
rect 37036 30982 37066 31034
rect 37066 30982 37078 31034
rect 37078 30982 37092 31034
rect 37116 30982 37130 31034
rect 37130 30982 37142 31034
rect 37142 30982 37172 31034
rect 37196 30982 37206 31034
rect 37206 30982 37252 31034
rect 36956 30980 37012 30982
rect 37036 30980 37092 30982
rect 37116 30980 37172 30982
rect 37196 30980 37252 30982
rect 41956 31034 42012 31036
rect 42036 31034 42092 31036
rect 42116 31034 42172 31036
rect 42196 31034 42252 31036
rect 41956 30982 42002 31034
rect 42002 30982 42012 31034
rect 42036 30982 42066 31034
rect 42066 30982 42078 31034
rect 42078 30982 42092 31034
rect 42116 30982 42130 31034
rect 42130 30982 42142 31034
rect 42142 30982 42172 31034
rect 42196 30982 42206 31034
rect 42206 30982 42252 31034
rect 41956 30980 42012 30982
rect 42036 30980 42092 30982
rect 42116 30980 42172 30982
rect 42196 30980 42252 30982
rect 46956 31034 47012 31036
rect 47036 31034 47092 31036
rect 47116 31034 47172 31036
rect 47196 31034 47252 31036
rect 46956 30982 47002 31034
rect 47002 30982 47012 31034
rect 47036 30982 47066 31034
rect 47066 30982 47078 31034
rect 47078 30982 47092 31034
rect 47116 30982 47130 31034
rect 47130 30982 47142 31034
rect 47142 30982 47172 31034
rect 47196 30982 47206 31034
rect 47206 30982 47252 31034
rect 46956 30980 47012 30982
rect 47036 30980 47092 30982
rect 47116 30980 47172 30982
rect 47196 30980 47252 30982
rect 51956 31034 52012 31036
rect 52036 31034 52092 31036
rect 52116 31034 52172 31036
rect 52196 31034 52252 31036
rect 51956 30982 52002 31034
rect 52002 30982 52012 31034
rect 52036 30982 52066 31034
rect 52066 30982 52078 31034
rect 52078 30982 52092 31034
rect 52116 30982 52130 31034
rect 52130 30982 52142 31034
rect 52142 30982 52172 31034
rect 52196 30982 52206 31034
rect 52206 30982 52252 31034
rect 51956 30980 52012 30982
rect 52036 30980 52092 30982
rect 52116 30980 52172 30982
rect 52196 30980 52252 30982
rect 56956 31034 57012 31036
rect 57036 31034 57092 31036
rect 57116 31034 57172 31036
rect 57196 31034 57252 31036
rect 56956 30982 57002 31034
rect 57002 30982 57012 31034
rect 57036 30982 57066 31034
rect 57066 30982 57078 31034
rect 57078 30982 57092 31034
rect 57116 30982 57130 31034
rect 57130 30982 57142 31034
rect 57142 30982 57172 31034
rect 57196 30982 57206 31034
rect 57206 30982 57252 31034
rect 56956 30980 57012 30982
rect 57036 30980 57092 30982
rect 57116 30980 57172 30982
rect 57196 30980 57252 30982
rect 2616 30490 2672 30492
rect 2696 30490 2752 30492
rect 2776 30490 2832 30492
rect 2856 30490 2912 30492
rect 2616 30438 2662 30490
rect 2662 30438 2672 30490
rect 2696 30438 2726 30490
rect 2726 30438 2738 30490
rect 2738 30438 2752 30490
rect 2776 30438 2790 30490
rect 2790 30438 2802 30490
rect 2802 30438 2832 30490
rect 2856 30438 2866 30490
rect 2866 30438 2912 30490
rect 2616 30436 2672 30438
rect 2696 30436 2752 30438
rect 2776 30436 2832 30438
rect 2856 30436 2912 30438
rect 7616 30490 7672 30492
rect 7696 30490 7752 30492
rect 7776 30490 7832 30492
rect 7856 30490 7912 30492
rect 7616 30438 7662 30490
rect 7662 30438 7672 30490
rect 7696 30438 7726 30490
rect 7726 30438 7738 30490
rect 7738 30438 7752 30490
rect 7776 30438 7790 30490
rect 7790 30438 7802 30490
rect 7802 30438 7832 30490
rect 7856 30438 7866 30490
rect 7866 30438 7912 30490
rect 7616 30436 7672 30438
rect 7696 30436 7752 30438
rect 7776 30436 7832 30438
rect 7856 30436 7912 30438
rect 12616 30490 12672 30492
rect 12696 30490 12752 30492
rect 12776 30490 12832 30492
rect 12856 30490 12912 30492
rect 12616 30438 12662 30490
rect 12662 30438 12672 30490
rect 12696 30438 12726 30490
rect 12726 30438 12738 30490
rect 12738 30438 12752 30490
rect 12776 30438 12790 30490
rect 12790 30438 12802 30490
rect 12802 30438 12832 30490
rect 12856 30438 12866 30490
rect 12866 30438 12912 30490
rect 12616 30436 12672 30438
rect 12696 30436 12752 30438
rect 12776 30436 12832 30438
rect 12856 30436 12912 30438
rect 17616 30490 17672 30492
rect 17696 30490 17752 30492
rect 17776 30490 17832 30492
rect 17856 30490 17912 30492
rect 17616 30438 17662 30490
rect 17662 30438 17672 30490
rect 17696 30438 17726 30490
rect 17726 30438 17738 30490
rect 17738 30438 17752 30490
rect 17776 30438 17790 30490
rect 17790 30438 17802 30490
rect 17802 30438 17832 30490
rect 17856 30438 17866 30490
rect 17866 30438 17912 30490
rect 17616 30436 17672 30438
rect 17696 30436 17752 30438
rect 17776 30436 17832 30438
rect 17856 30436 17912 30438
rect 22616 30490 22672 30492
rect 22696 30490 22752 30492
rect 22776 30490 22832 30492
rect 22856 30490 22912 30492
rect 22616 30438 22662 30490
rect 22662 30438 22672 30490
rect 22696 30438 22726 30490
rect 22726 30438 22738 30490
rect 22738 30438 22752 30490
rect 22776 30438 22790 30490
rect 22790 30438 22802 30490
rect 22802 30438 22832 30490
rect 22856 30438 22866 30490
rect 22866 30438 22912 30490
rect 22616 30436 22672 30438
rect 22696 30436 22752 30438
rect 22776 30436 22832 30438
rect 22856 30436 22912 30438
rect 27616 30490 27672 30492
rect 27696 30490 27752 30492
rect 27776 30490 27832 30492
rect 27856 30490 27912 30492
rect 27616 30438 27662 30490
rect 27662 30438 27672 30490
rect 27696 30438 27726 30490
rect 27726 30438 27738 30490
rect 27738 30438 27752 30490
rect 27776 30438 27790 30490
rect 27790 30438 27802 30490
rect 27802 30438 27832 30490
rect 27856 30438 27866 30490
rect 27866 30438 27912 30490
rect 27616 30436 27672 30438
rect 27696 30436 27752 30438
rect 27776 30436 27832 30438
rect 27856 30436 27912 30438
rect 32616 30490 32672 30492
rect 32696 30490 32752 30492
rect 32776 30490 32832 30492
rect 32856 30490 32912 30492
rect 32616 30438 32662 30490
rect 32662 30438 32672 30490
rect 32696 30438 32726 30490
rect 32726 30438 32738 30490
rect 32738 30438 32752 30490
rect 32776 30438 32790 30490
rect 32790 30438 32802 30490
rect 32802 30438 32832 30490
rect 32856 30438 32866 30490
rect 32866 30438 32912 30490
rect 32616 30436 32672 30438
rect 32696 30436 32752 30438
rect 32776 30436 32832 30438
rect 32856 30436 32912 30438
rect 37616 30490 37672 30492
rect 37696 30490 37752 30492
rect 37776 30490 37832 30492
rect 37856 30490 37912 30492
rect 37616 30438 37662 30490
rect 37662 30438 37672 30490
rect 37696 30438 37726 30490
rect 37726 30438 37738 30490
rect 37738 30438 37752 30490
rect 37776 30438 37790 30490
rect 37790 30438 37802 30490
rect 37802 30438 37832 30490
rect 37856 30438 37866 30490
rect 37866 30438 37912 30490
rect 37616 30436 37672 30438
rect 37696 30436 37752 30438
rect 37776 30436 37832 30438
rect 37856 30436 37912 30438
rect 42616 30490 42672 30492
rect 42696 30490 42752 30492
rect 42776 30490 42832 30492
rect 42856 30490 42912 30492
rect 42616 30438 42662 30490
rect 42662 30438 42672 30490
rect 42696 30438 42726 30490
rect 42726 30438 42738 30490
rect 42738 30438 42752 30490
rect 42776 30438 42790 30490
rect 42790 30438 42802 30490
rect 42802 30438 42832 30490
rect 42856 30438 42866 30490
rect 42866 30438 42912 30490
rect 42616 30436 42672 30438
rect 42696 30436 42752 30438
rect 42776 30436 42832 30438
rect 42856 30436 42912 30438
rect 47616 30490 47672 30492
rect 47696 30490 47752 30492
rect 47776 30490 47832 30492
rect 47856 30490 47912 30492
rect 47616 30438 47662 30490
rect 47662 30438 47672 30490
rect 47696 30438 47726 30490
rect 47726 30438 47738 30490
rect 47738 30438 47752 30490
rect 47776 30438 47790 30490
rect 47790 30438 47802 30490
rect 47802 30438 47832 30490
rect 47856 30438 47866 30490
rect 47866 30438 47912 30490
rect 47616 30436 47672 30438
rect 47696 30436 47752 30438
rect 47776 30436 47832 30438
rect 47856 30436 47912 30438
rect 52616 30490 52672 30492
rect 52696 30490 52752 30492
rect 52776 30490 52832 30492
rect 52856 30490 52912 30492
rect 52616 30438 52662 30490
rect 52662 30438 52672 30490
rect 52696 30438 52726 30490
rect 52726 30438 52738 30490
rect 52738 30438 52752 30490
rect 52776 30438 52790 30490
rect 52790 30438 52802 30490
rect 52802 30438 52832 30490
rect 52856 30438 52866 30490
rect 52866 30438 52912 30490
rect 52616 30436 52672 30438
rect 52696 30436 52752 30438
rect 52776 30436 52832 30438
rect 52856 30436 52912 30438
rect 57616 30490 57672 30492
rect 57696 30490 57752 30492
rect 57776 30490 57832 30492
rect 57856 30490 57912 30492
rect 57616 30438 57662 30490
rect 57662 30438 57672 30490
rect 57696 30438 57726 30490
rect 57726 30438 57738 30490
rect 57738 30438 57752 30490
rect 57776 30438 57790 30490
rect 57790 30438 57802 30490
rect 57802 30438 57832 30490
rect 57856 30438 57866 30490
rect 57866 30438 57912 30490
rect 57616 30436 57672 30438
rect 57696 30436 57752 30438
rect 57776 30436 57832 30438
rect 57856 30436 57912 30438
rect 58530 30232 58586 30288
rect 1956 29946 2012 29948
rect 2036 29946 2092 29948
rect 2116 29946 2172 29948
rect 2196 29946 2252 29948
rect 1956 29894 2002 29946
rect 2002 29894 2012 29946
rect 2036 29894 2066 29946
rect 2066 29894 2078 29946
rect 2078 29894 2092 29946
rect 2116 29894 2130 29946
rect 2130 29894 2142 29946
rect 2142 29894 2172 29946
rect 2196 29894 2206 29946
rect 2206 29894 2252 29946
rect 1956 29892 2012 29894
rect 2036 29892 2092 29894
rect 2116 29892 2172 29894
rect 2196 29892 2252 29894
rect 6956 29946 7012 29948
rect 7036 29946 7092 29948
rect 7116 29946 7172 29948
rect 7196 29946 7252 29948
rect 6956 29894 7002 29946
rect 7002 29894 7012 29946
rect 7036 29894 7066 29946
rect 7066 29894 7078 29946
rect 7078 29894 7092 29946
rect 7116 29894 7130 29946
rect 7130 29894 7142 29946
rect 7142 29894 7172 29946
rect 7196 29894 7206 29946
rect 7206 29894 7252 29946
rect 6956 29892 7012 29894
rect 7036 29892 7092 29894
rect 7116 29892 7172 29894
rect 7196 29892 7252 29894
rect 11956 29946 12012 29948
rect 12036 29946 12092 29948
rect 12116 29946 12172 29948
rect 12196 29946 12252 29948
rect 11956 29894 12002 29946
rect 12002 29894 12012 29946
rect 12036 29894 12066 29946
rect 12066 29894 12078 29946
rect 12078 29894 12092 29946
rect 12116 29894 12130 29946
rect 12130 29894 12142 29946
rect 12142 29894 12172 29946
rect 12196 29894 12206 29946
rect 12206 29894 12252 29946
rect 11956 29892 12012 29894
rect 12036 29892 12092 29894
rect 12116 29892 12172 29894
rect 12196 29892 12252 29894
rect 16956 29946 17012 29948
rect 17036 29946 17092 29948
rect 17116 29946 17172 29948
rect 17196 29946 17252 29948
rect 16956 29894 17002 29946
rect 17002 29894 17012 29946
rect 17036 29894 17066 29946
rect 17066 29894 17078 29946
rect 17078 29894 17092 29946
rect 17116 29894 17130 29946
rect 17130 29894 17142 29946
rect 17142 29894 17172 29946
rect 17196 29894 17206 29946
rect 17206 29894 17252 29946
rect 16956 29892 17012 29894
rect 17036 29892 17092 29894
rect 17116 29892 17172 29894
rect 17196 29892 17252 29894
rect 21956 29946 22012 29948
rect 22036 29946 22092 29948
rect 22116 29946 22172 29948
rect 22196 29946 22252 29948
rect 21956 29894 22002 29946
rect 22002 29894 22012 29946
rect 22036 29894 22066 29946
rect 22066 29894 22078 29946
rect 22078 29894 22092 29946
rect 22116 29894 22130 29946
rect 22130 29894 22142 29946
rect 22142 29894 22172 29946
rect 22196 29894 22206 29946
rect 22206 29894 22252 29946
rect 21956 29892 22012 29894
rect 22036 29892 22092 29894
rect 22116 29892 22172 29894
rect 22196 29892 22252 29894
rect 26956 29946 27012 29948
rect 27036 29946 27092 29948
rect 27116 29946 27172 29948
rect 27196 29946 27252 29948
rect 26956 29894 27002 29946
rect 27002 29894 27012 29946
rect 27036 29894 27066 29946
rect 27066 29894 27078 29946
rect 27078 29894 27092 29946
rect 27116 29894 27130 29946
rect 27130 29894 27142 29946
rect 27142 29894 27172 29946
rect 27196 29894 27206 29946
rect 27206 29894 27252 29946
rect 26956 29892 27012 29894
rect 27036 29892 27092 29894
rect 27116 29892 27172 29894
rect 27196 29892 27252 29894
rect 31956 29946 32012 29948
rect 32036 29946 32092 29948
rect 32116 29946 32172 29948
rect 32196 29946 32252 29948
rect 31956 29894 32002 29946
rect 32002 29894 32012 29946
rect 32036 29894 32066 29946
rect 32066 29894 32078 29946
rect 32078 29894 32092 29946
rect 32116 29894 32130 29946
rect 32130 29894 32142 29946
rect 32142 29894 32172 29946
rect 32196 29894 32206 29946
rect 32206 29894 32252 29946
rect 31956 29892 32012 29894
rect 32036 29892 32092 29894
rect 32116 29892 32172 29894
rect 32196 29892 32252 29894
rect 36956 29946 37012 29948
rect 37036 29946 37092 29948
rect 37116 29946 37172 29948
rect 37196 29946 37252 29948
rect 36956 29894 37002 29946
rect 37002 29894 37012 29946
rect 37036 29894 37066 29946
rect 37066 29894 37078 29946
rect 37078 29894 37092 29946
rect 37116 29894 37130 29946
rect 37130 29894 37142 29946
rect 37142 29894 37172 29946
rect 37196 29894 37206 29946
rect 37206 29894 37252 29946
rect 36956 29892 37012 29894
rect 37036 29892 37092 29894
rect 37116 29892 37172 29894
rect 37196 29892 37252 29894
rect 41956 29946 42012 29948
rect 42036 29946 42092 29948
rect 42116 29946 42172 29948
rect 42196 29946 42252 29948
rect 41956 29894 42002 29946
rect 42002 29894 42012 29946
rect 42036 29894 42066 29946
rect 42066 29894 42078 29946
rect 42078 29894 42092 29946
rect 42116 29894 42130 29946
rect 42130 29894 42142 29946
rect 42142 29894 42172 29946
rect 42196 29894 42206 29946
rect 42206 29894 42252 29946
rect 41956 29892 42012 29894
rect 42036 29892 42092 29894
rect 42116 29892 42172 29894
rect 42196 29892 42252 29894
rect 46956 29946 47012 29948
rect 47036 29946 47092 29948
rect 47116 29946 47172 29948
rect 47196 29946 47252 29948
rect 46956 29894 47002 29946
rect 47002 29894 47012 29946
rect 47036 29894 47066 29946
rect 47066 29894 47078 29946
rect 47078 29894 47092 29946
rect 47116 29894 47130 29946
rect 47130 29894 47142 29946
rect 47142 29894 47172 29946
rect 47196 29894 47206 29946
rect 47206 29894 47252 29946
rect 46956 29892 47012 29894
rect 47036 29892 47092 29894
rect 47116 29892 47172 29894
rect 47196 29892 47252 29894
rect 51956 29946 52012 29948
rect 52036 29946 52092 29948
rect 52116 29946 52172 29948
rect 52196 29946 52252 29948
rect 51956 29894 52002 29946
rect 52002 29894 52012 29946
rect 52036 29894 52066 29946
rect 52066 29894 52078 29946
rect 52078 29894 52092 29946
rect 52116 29894 52130 29946
rect 52130 29894 52142 29946
rect 52142 29894 52172 29946
rect 52196 29894 52206 29946
rect 52206 29894 52252 29946
rect 51956 29892 52012 29894
rect 52036 29892 52092 29894
rect 52116 29892 52172 29894
rect 52196 29892 52252 29894
rect 56956 29946 57012 29948
rect 57036 29946 57092 29948
rect 57116 29946 57172 29948
rect 57196 29946 57252 29948
rect 56956 29894 57002 29946
rect 57002 29894 57012 29946
rect 57036 29894 57066 29946
rect 57066 29894 57078 29946
rect 57078 29894 57092 29946
rect 57116 29894 57130 29946
rect 57130 29894 57142 29946
rect 57142 29894 57172 29946
rect 57196 29894 57206 29946
rect 57206 29894 57252 29946
rect 56956 29892 57012 29894
rect 57036 29892 57092 29894
rect 57116 29892 57172 29894
rect 57196 29892 57252 29894
rect 58530 29416 58586 29472
rect 2616 29402 2672 29404
rect 2696 29402 2752 29404
rect 2776 29402 2832 29404
rect 2856 29402 2912 29404
rect 2616 29350 2662 29402
rect 2662 29350 2672 29402
rect 2696 29350 2726 29402
rect 2726 29350 2738 29402
rect 2738 29350 2752 29402
rect 2776 29350 2790 29402
rect 2790 29350 2802 29402
rect 2802 29350 2832 29402
rect 2856 29350 2866 29402
rect 2866 29350 2912 29402
rect 2616 29348 2672 29350
rect 2696 29348 2752 29350
rect 2776 29348 2832 29350
rect 2856 29348 2912 29350
rect 7616 29402 7672 29404
rect 7696 29402 7752 29404
rect 7776 29402 7832 29404
rect 7856 29402 7912 29404
rect 7616 29350 7662 29402
rect 7662 29350 7672 29402
rect 7696 29350 7726 29402
rect 7726 29350 7738 29402
rect 7738 29350 7752 29402
rect 7776 29350 7790 29402
rect 7790 29350 7802 29402
rect 7802 29350 7832 29402
rect 7856 29350 7866 29402
rect 7866 29350 7912 29402
rect 7616 29348 7672 29350
rect 7696 29348 7752 29350
rect 7776 29348 7832 29350
rect 7856 29348 7912 29350
rect 12616 29402 12672 29404
rect 12696 29402 12752 29404
rect 12776 29402 12832 29404
rect 12856 29402 12912 29404
rect 12616 29350 12662 29402
rect 12662 29350 12672 29402
rect 12696 29350 12726 29402
rect 12726 29350 12738 29402
rect 12738 29350 12752 29402
rect 12776 29350 12790 29402
rect 12790 29350 12802 29402
rect 12802 29350 12832 29402
rect 12856 29350 12866 29402
rect 12866 29350 12912 29402
rect 12616 29348 12672 29350
rect 12696 29348 12752 29350
rect 12776 29348 12832 29350
rect 12856 29348 12912 29350
rect 17616 29402 17672 29404
rect 17696 29402 17752 29404
rect 17776 29402 17832 29404
rect 17856 29402 17912 29404
rect 17616 29350 17662 29402
rect 17662 29350 17672 29402
rect 17696 29350 17726 29402
rect 17726 29350 17738 29402
rect 17738 29350 17752 29402
rect 17776 29350 17790 29402
rect 17790 29350 17802 29402
rect 17802 29350 17832 29402
rect 17856 29350 17866 29402
rect 17866 29350 17912 29402
rect 17616 29348 17672 29350
rect 17696 29348 17752 29350
rect 17776 29348 17832 29350
rect 17856 29348 17912 29350
rect 22616 29402 22672 29404
rect 22696 29402 22752 29404
rect 22776 29402 22832 29404
rect 22856 29402 22912 29404
rect 22616 29350 22662 29402
rect 22662 29350 22672 29402
rect 22696 29350 22726 29402
rect 22726 29350 22738 29402
rect 22738 29350 22752 29402
rect 22776 29350 22790 29402
rect 22790 29350 22802 29402
rect 22802 29350 22832 29402
rect 22856 29350 22866 29402
rect 22866 29350 22912 29402
rect 22616 29348 22672 29350
rect 22696 29348 22752 29350
rect 22776 29348 22832 29350
rect 22856 29348 22912 29350
rect 27616 29402 27672 29404
rect 27696 29402 27752 29404
rect 27776 29402 27832 29404
rect 27856 29402 27912 29404
rect 27616 29350 27662 29402
rect 27662 29350 27672 29402
rect 27696 29350 27726 29402
rect 27726 29350 27738 29402
rect 27738 29350 27752 29402
rect 27776 29350 27790 29402
rect 27790 29350 27802 29402
rect 27802 29350 27832 29402
rect 27856 29350 27866 29402
rect 27866 29350 27912 29402
rect 27616 29348 27672 29350
rect 27696 29348 27752 29350
rect 27776 29348 27832 29350
rect 27856 29348 27912 29350
rect 32616 29402 32672 29404
rect 32696 29402 32752 29404
rect 32776 29402 32832 29404
rect 32856 29402 32912 29404
rect 32616 29350 32662 29402
rect 32662 29350 32672 29402
rect 32696 29350 32726 29402
rect 32726 29350 32738 29402
rect 32738 29350 32752 29402
rect 32776 29350 32790 29402
rect 32790 29350 32802 29402
rect 32802 29350 32832 29402
rect 32856 29350 32866 29402
rect 32866 29350 32912 29402
rect 32616 29348 32672 29350
rect 32696 29348 32752 29350
rect 32776 29348 32832 29350
rect 32856 29348 32912 29350
rect 37616 29402 37672 29404
rect 37696 29402 37752 29404
rect 37776 29402 37832 29404
rect 37856 29402 37912 29404
rect 37616 29350 37662 29402
rect 37662 29350 37672 29402
rect 37696 29350 37726 29402
rect 37726 29350 37738 29402
rect 37738 29350 37752 29402
rect 37776 29350 37790 29402
rect 37790 29350 37802 29402
rect 37802 29350 37832 29402
rect 37856 29350 37866 29402
rect 37866 29350 37912 29402
rect 37616 29348 37672 29350
rect 37696 29348 37752 29350
rect 37776 29348 37832 29350
rect 37856 29348 37912 29350
rect 42616 29402 42672 29404
rect 42696 29402 42752 29404
rect 42776 29402 42832 29404
rect 42856 29402 42912 29404
rect 42616 29350 42662 29402
rect 42662 29350 42672 29402
rect 42696 29350 42726 29402
rect 42726 29350 42738 29402
rect 42738 29350 42752 29402
rect 42776 29350 42790 29402
rect 42790 29350 42802 29402
rect 42802 29350 42832 29402
rect 42856 29350 42866 29402
rect 42866 29350 42912 29402
rect 42616 29348 42672 29350
rect 42696 29348 42752 29350
rect 42776 29348 42832 29350
rect 42856 29348 42912 29350
rect 47616 29402 47672 29404
rect 47696 29402 47752 29404
rect 47776 29402 47832 29404
rect 47856 29402 47912 29404
rect 47616 29350 47662 29402
rect 47662 29350 47672 29402
rect 47696 29350 47726 29402
rect 47726 29350 47738 29402
rect 47738 29350 47752 29402
rect 47776 29350 47790 29402
rect 47790 29350 47802 29402
rect 47802 29350 47832 29402
rect 47856 29350 47866 29402
rect 47866 29350 47912 29402
rect 47616 29348 47672 29350
rect 47696 29348 47752 29350
rect 47776 29348 47832 29350
rect 47856 29348 47912 29350
rect 52616 29402 52672 29404
rect 52696 29402 52752 29404
rect 52776 29402 52832 29404
rect 52856 29402 52912 29404
rect 52616 29350 52662 29402
rect 52662 29350 52672 29402
rect 52696 29350 52726 29402
rect 52726 29350 52738 29402
rect 52738 29350 52752 29402
rect 52776 29350 52790 29402
rect 52790 29350 52802 29402
rect 52802 29350 52832 29402
rect 52856 29350 52866 29402
rect 52866 29350 52912 29402
rect 52616 29348 52672 29350
rect 52696 29348 52752 29350
rect 52776 29348 52832 29350
rect 52856 29348 52912 29350
rect 57616 29402 57672 29404
rect 57696 29402 57752 29404
rect 57776 29402 57832 29404
rect 57856 29402 57912 29404
rect 57616 29350 57662 29402
rect 57662 29350 57672 29402
rect 57696 29350 57726 29402
rect 57726 29350 57738 29402
rect 57738 29350 57752 29402
rect 57776 29350 57790 29402
rect 57790 29350 57802 29402
rect 57802 29350 57832 29402
rect 57856 29350 57866 29402
rect 57866 29350 57912 29402
rect 57616 29348 57672 29350
rect 57696 29348 57752 29350
rect 57776 29348 57832 29350
rect 57856 29348 57912 29350
rect 1956 28858 2012 28860
rect 2036 28858 2092 28860
rect 2116 28858 2172 28860
rect 2196 28858 2252 28860
rect 1956 28806 2002 28858
rect 2002 28806 2012 28858
rect 2036 28806 2066 28858
rect 2066 28806 2078 28858
rect 2078 28806 2092 28858
rect 2116 28806 2130 28858
rect 2130 28806 2142 28858
rect 2142 28806 2172 28858
rect 2196 28806 2206 28858
rect 2206 28806 2252 28858
rect 1956 28804 2012 28806
rect 2036 28804 2092 28806
rect 2116 28804 2172 28806
rect 2196 28804 2252 28806
rect 6956 28858 7012 28860
rect 7036 28858 7092 28860
rect 7116 28858 7172 28860
rect 7196 28858 7252 28860
rect 6956 28806 7002 28858
rect 7002 28806 7012 28858
rect 7036 28806 7066 28858
rect 7066 28806 7078 28858
rect 7078 28806 7092 28858
rect 7116 28806 7130 28858
rect 7130 28806 7142 28858
rect 7142 28806 7172 28858
rect 7196 28806 7206 28858
rect 7206 28806 7252 28858
rect 6956 28804 7012 28806
rect 7036 28804 7092 28806
rect 7116 28804 7172 28806
rect 7196 28804 7252 28806
rect 11956 28858 12012 28860
rect 12036 28858 12092 28860
rect 12116 28858 12172 28860
rect 12196 28858 12252 28860
rect 11956 28806 12002 28858
rect 12002 28806 12012 28858
rect 12036 28806 12066 28858
rect 12066 28806 12078 28858
rect 12078 28806 12092 28858
rect 12116 28806 12130 28858
rect 12130 28806 12142 28858
rect 12142 28806 12172 28858
rect 12196 28806 12206 28858
rect 12206 28806 12252 28858
rect 11956 28804 12012 28806
rect 12036 28804 12092 28806
rect 12116 28804 12172 28806
rect 12196 28804 12252 28806
rect 16956 28858 17012 28860
rect 17036 28858 17092 28860
rect 17116 28858 17172 28860
rect 17196 28858 17252 28860
rect 16956 28806 17002 28858
rect 17002 28806 17012 28858
rect 17036 28806 17066 28858
rect 17066 28806 17078 28858
rect 17078 28806 17092 28858
rect 17116 28806 17130 28858
rect 17130 28806 17142 28858
rect 17142 28806 17172 28858
rect 17196 28806 17206 28858
rect 17206 28806 17252 28858
rect 16956 28804 17012 28806
rect 17036 28804 17092 28806
rect 17116 28804 17172 28806
rect 17196 28804 17252 28806
rect 21956 28858 22012 28860
rect 22036 28858 22092 28860
rect 22116 28858 22172 28860
rect 22196 28858 22252 28860
rect 21956 28806 22002 28858
rect 22002 28806 22012 28858
rect 22036 28806 22066 28858
rect 22066 28806 22078 28858
rect 22078 28806 22092 28858
rect 22116 28806 22130 28858
rect 22130 28806 22142 28858
rect 22142 28806 22172 28858
rect 22196 28806 22206 28858
rect 22206 28806 22252 28858
rect 21956 28804 22012 28806
rect 22036 28804 22092 28806
rect 22116 28804 22172 28806
rect 22196 28804 22252 28806
rect 26956 28858 27012 28860
rect 27036 28858 27092 28860
rect 27116 28858 27172 28860
rect 27196 28858 27252 28860
rect 26956 28806 27002 28858
rect 27002 28806 27012 28858
rect 27036 28806 27066 28858
rect 27066 28806 27078 28858
rect 27078 28806 27092 28858
rect 27116 28806 27130 28858
rect 27130 28806 27142 28858
rect 27142 28806 27172 28858
rect 27196 28806 27206 28858
rect 27206 28806 27252 28858
rect 26956 28804 27012 28806
rect 27036 28804 27092 28806
rect 27116 28804 27172 28806
rect 27196 28804 27252 28806
rect 31956 28858 32012 28860
rect 32036 28858 32092 28860
rect 32116 28858 32172 28860
rect 32196 28858 32252 28860
rect 31956 28806 32002 28858
rect 32002 28806 32012 28858
rect 32036 28806 32066 28858
rect 32066 28806 32078 28858
rect 32078 28806 32092 28858
rect 32116 28806 32130 28858
rect 32130 28806 32142 28858
rect 32142 28806 32172 28858
rect 32196 28806 32206 28858
rect 32206 28806 32252 28858
rect 31956 28804 32012 28806
rect 32036 28804 32092 28806
rect 32116 28804 32172 28806
rect 32196 28804 32252 28806
rect 36956 28858 37012 28860
rect 37036 28858 37092 28860
rect 37116 28858 37172 28860
rect 37196 28858 37252 28860
rect 36956 28806 37002 28858
rect 37002 28806 37012 28858
rect 37036 28806 37066 28858
rect 37066 28806 37078 28858
rect 37078 28806 37092 28858
rect 37116 28806 37130 28858
rect 37130 28806 37142 28858
rect 37142 28806 37172 28858
rect 37196 28806 37206 28858
rect 37206 28806 37252 28858
rect 36956 28804 37012 28806
rect 37036 28804 37092 28806
rect 37116 28804 37172 28806
rect 37196 28804 37252 28806
rect 41956 28858 42012 28860
rect 42036 28858 42092 28860
rect 42116 28858 42172 28860
rect 42196 28858 42252 28860
rect 41956 28806 42002 28858
rect 42002 28806 42012 28858
rect 42036 28806 42066 28858
rect 42066 28806 42078 28858
rect 42078 28806 42092 28858
rect 42116 28806 42130 28858
rect 42130 28806 42142 28858
rect 42142 28806 42172 28858
rect 42196 28806 42206 28858
rect 42206 28806 42252 28858
rect 41956 28804 42012 28806
rect 42036 28804 42092 28806
rect 42116 28804 42172 28806
rect 42196 28804 42252 28806
rect 46956 28858 47012 28860
rect 47036 28858 47092 28860
rect 47116 28858 47172 28860
rect 47196 28858 47252 28860
rect 46956 28806 47002 28858
rect 47002 28806 47012 28858
rect 47036 28806 47066 28858
rect 47066 28806 47078 28858
rect 47078 28806 47092 28858
rect 47116 28806 47130 28858
rect 47130 28806 47142 28858
rect 47142 28806 47172 28858
rect 47196 28806 47206 28858
rect 47206 28806 47252 28858
rect 46956 28804 47012 28806
rect 47036 28804 47092 28806
rect 47116 28804 47172 28806
rect 47196 28804 47252 28806
rect 51956 28858 52012 28860
rect 52036 28858 52092 28860
rect 52116 28858 52172 28860
rect 52196 28858 52252 28860
rect 51956 28806 52002 28858
rect 52002 28806 52012 28858
rect 52036 28806 52066 28858
rect 52066 28806 52078 28858
rect 52078 28806 52092 28858
rect 52116 28806 52130 28858
rect 52130 28806 52142 28858
rect 52142 28806 52172 28858
rect 52196 28806 52206 28858
rect 52206 28806 52252 28858
rect 51956 28804 52012 28806
rect 52036 28804 52092 28806
rect 52116 28804 52172 28806
rect 52196 28804 52252 28806
rect 56956 28858 57012 28860
rect 57036 28858 57092 28860
rect 57116 28858 57172 28860
rect 57196 28858 57252 28860
rect 56956 28806 57002 28858
rect 57002 28806 57012 28858
rect 57036 28806 57066 28858
rect 57066 28806 57078 28858
rect 57078 28806 57092 28858
rect 57116 28806 57130 28858
rect 57130 28806 57142 28858
rect 57142 28806 57172 28858
rect 57196 28806 57206 28858
rect 57206 28806 57252 28858
rect 56956 28804 57012 28806
rect 57036 28804 57092 28806
rect 57116 28804 57172 28806
rect 57196 28804 57252 28806
rect 58530 28600 58586 28656
rect 2616 28314 2672 28316
rect 2696 28314 2752 28316
rect 2776 28314 2832 28316
rect 2856 28314 2912 28316
rect 2616 28262 2662 28314
rect 2662 28262 2672 28314
rect 2696 28262 2726 28314
rect 2726 28262 2738 28314
rect 2738 28262 2752 28314
rect 2776 28262 2790 28314
rect 2790 28262 2802 28314
rect 2802 28262 2832 28314
rect 2856 28262 2866 28314
rect 2866 28262 2912 28314
rect 2616 28260 2672 28262
rect 2696 28260 2752 28262
rect 2776 28260 2832 28262
rect 2856 28260 2912 28262
rect 7616 28314 7672 28316
rect 7696 28314 7752 28316
rect 7776 28314 7832 28316
rect 7856 28314 7912 28316
rect 7616 28262 7662 28314
rect 7662 28262 7672 28314
rect 7696 28262 7726 28314
rect 7726 28262 7738 28314
rect 7738 28262 7752 28314
rect 7776 28262 7790 28314
rect 7790 28262 7802 28314
rect 7802 28262 7832 28314
rect 7856 28262 7866 28314
rect 7866 28262 7912 28314
rect 7616 28260 7672 28262
rect 7696 28260 7752 28262
rect 7776 28260 7832 28262
rect 7856 28260 7912 28262
rect 12616 28314 12672 28316
rect 12696 28314 12752 28316
rect 12776 28314 12832 28316
rect 12856 28314 12912 28316
rect 12616 28262 12662 28314
rect 12662 28262 12672 28314
rect 12696 28262 12726 28314
rect 12726 28262 12738 28314
rect 12738 28262 12752 28314
rect 12776 28262 12790 28314
rect 12790 28262 12802 28314
rect 12802 28262 12832 28314
rect 12856 28262 12866 28314
rect 12866 28262 12912 28314
rect 12616 28260 12672 28262
rect 12696 28260 12752 28262
rect 12776 28260 12832 28262
rect 12856 28260 12912 28262
rect 17616 28314 17672 28316
rect 17696 28314 17752 28316
rect 17776 28314 17832 28316
rect 17856 28314 17912 28316
rect 17616 28262 17662 28314
rect 17662 28262 17672 28314
rect 17696 28262 17726 28314
rect 17726 28262 17738 28314
rect 17738 28262 17752 28314
rect 17776 28262 17790 28314
rect 17790 28262 17802 28314
rect 17802 28262 17832 28314
rect 17856 28262 17866 28314
rect 17866 28262 17912 28314
rect 17616 28260 17672 28262
rect 17696 28260 17752 28262
rect 17776 28260 17832 28262
rect 17856 28260 17912 28262
rect 22616 28314 22672 28316
rect 22696 28314 22752 28316
rect 22776 28314 22832 28316
rect 22856 28314 22912 28316
rect 22616 28262 22662 28314
rect 22662 28262 22672 28314
rect 22696 28262 22726 28314
rect 22726 28262 22738 28314
rect 22738 28262 22752 28314
rect 22776 28262 22790 28314
rect 22790 28262 22802 28314
rect 22802 28262 22832 28314
rect 22856 28262 22866 28314
rect 22866 28262 22912 28314
rect 22616 28260 22672 28262
rect 22696 28260 22752 28262
rect 22776 28260 22832 28262
rect 22856 28260 22912 28262
rect 27616 28314 27672 28316
rect 27696 28314 27752 28316
rect 27776 28314 27832 28316
rect 27856 28314 27912 28316
rect 27616 28262 27662 28314
rect 27662 28262 27672 28314
rect 27696 28262 27726 28314
rect 27726 28262 27738 28314
rect 27738 28262 27752 28314
rect 27776 28262 27790 28314
rect 27790 28262 27802 28314
rect 27802 28262 27832 28314
rect 27856 28262 27866 28314
rect 27866 28262 27912 28314
rect 27616 28260 27672 28262
rect 27696 28260 27752 28262
rect 27776 28260 27832 28262
rect 27856 28260 27912 28262
rect 32616 28314 32672 28316
rect 32696 28314 32752 28316
rect 32776 28314 32832 28316
rect 32856 28314 32912 28316
rect 32616 28262 32662 28314
rect 32662 28262 32672 28314
rect 32696 28262 32726 28314
rect 32726 28262 32738 28314
rect 32738 28262 32752 28314
rect 32776 28262 32790 28314
rect 32790 28262 32802 28314
rect 32802 28262 32832 28314
rect 32856 28262 32866 28314
rect 32866 28262 32912 28314
rect 32616 28260 32672 28262
rect 32696 28260 32752 28262
rect 32776 28260 32832 28262
rect 32856 28260 32912 28262
rect 37616 28314 37672 28316
rect 37696 28314 37752 28316
rect 37776 28314 37832 28316
rect 37856 28314 37912 28316
rect 37616 28262 37662 28314
rect 37662 28262 37672 28314
rect 37696 28262 37726 28314
rect 37726 28262 37738 28314
rect 37738 28262 37752 28314
rect 37776 28262 37790 28314
rect 37790 28262 37802 28314
rect 37802 28262 37832 28314
rect 37856 28262 37866 28314
rect 37866 28262 37912 28314
rect 37616 28260 37672 28262
rect 37696 28260 37752 28262
rect 37776 28260 37832 28262
rect 37856 28260 37912 28262
rect 42616 28314 42672 28316
rect 42696 28314 42752 28316
rect 42776 28314 42832 28316
rect 42856 28314 42912 28316
rect 42616 28262 42662 28314
rect 42662 28262 42672 28314
rect 42696 28262 42726 28314
rect 42726 28262 42738 28314
rect 42738 28262 42752 28314
rect 42776 28262 42790 28314
rect 42790 28262 42802 28314
rect 42802 28262 42832 28314
rect 42856 28262 42866 28314
rect 42866 28262 42912 28314
rect 42616 28260 42672 28262
rect 42696 28260 42752 28262
rect 42776 28260 42832 28262
rect 42856 28260 42912 28262
rect 47616 28314 47672 28316
rect 47696 28314 47752 28316
rect 47776 28314 47832 28316
rect 47856 28314 47912 28316
rect 47616 28262 47662 28314
rect 47662 28262 47672 28314
rect 47696 28262 47726 28314
rect 47726 28262 47738 28314
rect 47738 28262 47752 28314
rect 47776 28262 47790 28314
rect 47790 28262 47802 28314
rect 47802 28262 47832 28314
rect 47856 28262 47866 28314
rect 47866 28262 47912 28314
rect 47616 28260 47672 28262
rect 47696 28260 47752 28262
rect 47776 28260 47832 28262
rect 47856 28260 47912 28262
rect 52616 28314 52672 28316
rect 52696 28314 52752 28316
rect 52776 28314 52832 28316
rect 52856 28314 52912 28316
rect 52616 28262 52662 28314
rect 52662 28262 52672 28314
rect 52696 28262 52726 28314
rect 52726 28262 52738 28314
rect 52738 28262 52752 28314
rect 52776 28262 52790 28314
rect 52790 28262 52802 28314
rect 52802 28262 52832 28314
rect 52856 28262 52866 28314
rect 52866 28262 52912 28314
rect 52616 28260 52672 28262
rect 52696 28260 52752 28262
rect 52776 28260 52832 28262
rect 52856 28260 52912 28262
rect 57616 28314 57672 28316
rect 57696 28314 57752 28316
rect 57776 28314 57832 28316
rect 57856 28314 57912 28316
rect 57616 28262 57662 28314
rect 57662 28262 57672 28314
rect 57696 28262 57726 28314
rect 57726 28262 57738 28314
rect 57738 28262 57752 28314
rect 57776 28262 57790 28314
rect 57790 28262 57802 28314
rect 57802 28262 57832 28314
rect 57856 28262 57866 28314
rect 57866 28262 57912 28314
rect 57616 28260 57672 28262
rect 57696 28260 57752 28262
rect 57776 28260 57832 28262
rect 57856 28260 57912 28262
rect 58530 27820 58532 27840
rect 58532 27820 58584 27840
rect 58584 27820 58586 27840
rect 58530 27784 58586 27820
rect 1956 27770 2012 27772
rect 2036 27770 2092 27772
rect 2116 27770 2172 27772
rect 2196 27770 2252 27772
rect 1956 27718 2002 27770
rect 2002 27718 2012 27770
rect 2036 27718 2066 27770
rect 2066 27718 2078 27770
rect 2078 27718 2092 27770
rect 2116 27718 2130 27770
rect 2130 27718 2142 27770
rect 2142 27718 2172 27770
rect 2196 27718 2206 27770
rect 2206 27718 2252 27770
rect 1956 27716 2012 27718
rect 2036 27716 2092 27718
rect 2116 27716 2172 27718
rect 2196 27716 2252 27718
rect 6956 27770 7012 27772
rect 7036 27770 7092 27772
rect 7116 27770 7172 27772
rect 7196 27770 7252 27772
rect 6956 27718 7002 27770
rect 7002 27718 7012 27770
rect 7036 27718 7066 27770
rect 7066 27718 7078 27770
rect 7078 27718 7092 27770
rect 7116 27718 7130 27770
rect 7130 27718 7142 27770
rect 7142 27718 7172 27770
rect 7196 27718 7206 27770
rect 7206 27718 7252 27770
rect 6956 27716 7012 27718
rect 7036 27716 7092 27718
rect 7116 27716 7172 27718
rect 7196 27716 7252 27718
rect 11956 27770 12012 27772
rect 12036 27770 12092 27772
rect 12116 27770 12172 27772
rect 12196 27770 12252 27772
rect 11956 27718 12002 27770
rect 12002 27718 12012 27770
rect 12036 27718 12066 27770
rect 12066 27718 12078 27770
rect 12078 27718 12092 27770
rect 12116 27718 12130 27770
rect 12130 27718 12142 27770
rect 12142 27718 12172 27770
rect 12196 27718 12206 27770
rect 12206 27718 12252 27770
rect 11956 27716 12012 27718
rect 12036 27716 12092 27718
rect 12116 27716 12172 27718
rect 12196 27716 12252 27718
rect 16956 27770 17012 27772
rect 17036 27770 17092 27772
rect 17116 27770 17172 27772
rect 17196 27770 17252 27772
rect 16956 27718 17002 27770
rect 17002 27718 17012 27770
rect 17036 27718 17066 27770
rect 17066 27718 17078 27770
rect 17078 27718 17092 27770
rect 17116 27718 17130 27770
rect 17130 27718 17142 27770
rect 17142 27718 17172 27770
rect 17196 27718 17206 27770
rect 17206 27718 17252 27770
rect 16956 27716 17012 27718
rect 17036 27716 17092 27718
rect 17116 27716 17172 27718
rect 17196 27716 17252 27718
rect 21956 27770 22012 27772
rect 22036 27770 22092 27772
rect 22116 27770 22172 27772
rect 22196 27770 22252 27772
rect 21956 27718 22002 27770
rect 22002 27718 22012 27770
rect 22036 27718 22066 27770
rect 22066 27718 22078 27770
rect 22078 27718 22092 27770
rect 22116 27718 22130 27770
rect 22130 27718 22142 27770
rect 22142 27718 22172 27770
rect 22196 27718 22206 27770
rect 22206 27718 22252 27770
rect 21956 27716 22012 27718
rect 22036 27716 22092 27718
rect 22116 27716 22172 27718
rect 22196 27716 22252 27718
rect 26956 27770 27012 27772
rect 27036 27770 27092 27772
rect 27116 27770 27172 27772
rect 27196 27770 27252 27772
rect 26956 27718 27002 27770
rect 27002 27718 27012 27770
rect 27036 27718 27066 27770
rect 27066 27718 27078 27770
rect 27078 27718 27092 27770
rect 27116 27718 27130 27770
rect 27130 27718 27142 27770
rect 27142 27718 27172 27770
rect 27196 27718 27206 27770
rect 27206 27718 27252 27770
rect 26956 27716 27012 27718
rect 27036 27716 27092 27718
rect 27116 27716 27172 27718
rect 27196 27716 27252 27718
rect 31956 27770 32012 27772
rect 32036 27770 32092 27772
rect 32116 27770 32172 27772
rect 32196 27770 32252 27772
rect 31956 27718 32002 27770
rect 32002 27718 32012 27770
rect 32036 27718 32066 27770
rect 32066 27718 32078 27770
rect 32078 27718 32092 27770
rect 32116 27718 32130 27770
rect 32130 27718 32142 27770
rect 32142 27718 32172 27770
rect 32196 27718 32206 27770
rect 32206 27718 32252 27770
rect 31956 27716 32012 27718
rect 32036 27716 32092 27718
rect 32116 27716 32172 27718
rect 32196 27716 32252 27718
rect 36956 27770 37012 27772
rect 37036 27770 37092 27772
rect 37116 27770 37172 27772
rect 37196 27770 37252 27772
rect 36956 27718 37002 27770
rect 37002 27718 37012 27770
rect 37036 27718 37066 27770
rect 37066 27718 37078 27770
rect 37078 27718 37092 27770
rect 37116 27718 37130 27770
rect 37130 27718 37142 27770
rect 37142 27718 37172 27770
rect 37196 27718 37206 27770
rect 37206 27718 37252 27770
rect 36956 27716 37012 27718
rect 37036 27716 37092 27718
rect 37116 27716 37172 27718
rect 37196 27716 37252 27718
rect 41956 27770 42012 27772
rect 42036 27770 42092 27772
rect 42116 27770 42172 27772
rect 42196 27770 42252 27772
rect 41956 27718 42002 27770
rect 42002 27718 42012 27770
rect 42036 27718 42066 27770
rect 42066 27718 42078 27770
rect 42078 27718 42092 27770
rect 42116 27718 42130 27770
rect 42130 27718 42142 27770
rect 42142 27718 42172 27770
rect 42196 27718 42206 27770
rect 42206 27718 42252 27770
rect 41956 27716 42012 27718
rect 42036 27716 42092 27718
rect 42116 27716 42172 27718
rect 42196 27716 42252 27718
rect 46956 27770 47012 27772
rect 47036 27770 47092 27772
rect 47116 27770 47172 27772
rect 47196 27770 47252 27772
rect 46956 27718 47002 27770
rect 47002 27718 47012 27770
rect 47036 27718 47066 27770
rect 47066 27718 47078 27770
rect 47078 27718 47092 27770
rect 47116 27718 47130 27770
rect 47130 27718 47142 27770
rect 47142 27718 47172 27770
rect 47196 27718 47206 27770
rect 47206 27718 47252 27770
rect 46956 27716 47012 27718
rect 47036 27716 47092 27718
rect 47116 27716 47172 27718
rect 47196 27716 47252 27718
rect 51956 27770 52012 27772
rect 52036 27770 52092 27772
rect 52116 27770 52172 27772
rect 52196 27770 52252 27772
rect 51956 27718 52002 27770
rect 52002 27718 52012 27770
rect 52036 27718 52066 27770
rect 52066 27718 52078 27770
rect 52078 27718 52092 27770
rect 52116 27718 52130 27770
rect 52130 27718 52142 27770
rect 52142 27718 52172 27770
rect 52196 27718 52206 27770
rect 52206 27718 52252 27770
rect 51956 27716 52012 27718
rect 52036 27716 52092 27718
rect 52116 27716 52172 27718
rect 52196 27716 52252 27718
rect 56956 27770 57012 27772
rect 57036 27770 57092 27772
rect 57116 27770 57172 27772
rect 57196 27770 57252 27772
rect 56956 27718 57002 27770
rect 57002 27718 57012 27770
rect 57036 27718 57066 27770
rect 57066 27718 57078 27770
rect 57078 27718 57092 27770
rect 57116 27718 57130 27770
rect 57130 27718 57142 27770
rect 57142 27718 57172 27770
rect 57196 27718 57206 27770
rect 57206 27718 57252 27770
rect 56956 27716 57012 27718
rect 57036 27716 57092 27718
rect 57116 27716 57172 27718
rect 57196 27716 57252 27718
rect 2616 27226 2672 27228
rect 2696 27226 2752 27228
rect 2776 27226 2832 27228
rect 2856 27226 2912 27228
rect 2616 27174 2662 27226
rect 2662 27174 2672 27226
rect 2696 27174 2726 27226
rect 2726 27174 2738 27226
rect 2738 27174 2752 27226
rect 2776 27174 2790 27226
rect 2790 27174 2802 27226
rect 2802 27174 2832 27226
rect 2856 27174 2866 27226
rect 2866 27174 2912 27226
rect 2616 27172 2672 27174
rect 2696 27172 2752 27174
rect 2776 27172 2832 27174
rect 2856 27172 2912 27174
rect 7616 27226 7672 27228
rect 7696 27226 7752 27228
rect 7776 27226 7832 27228
rect 7856 27226 7912 27228
rect 7616 27174 7662 27226
rect 7662 27174 7672 27226
rect 7696 27174 7726 27226
rect 7726 27174 7738 27226
rect 7738 27174 7752 27226
rect 7776 27174 7790 27226
rect 7790 27174 7802 27226
rect 7802 27174 7832 27226
rect 7856 27174 7866 27226
rect 7866 27174 7912 27226
rect 7616 27172 7672 27174
rect 7696 27172 7752 27174
rect 7776 27172 7832 27174
rect 7856 27172 7912 27174
rect 12616 27226 12672 27228
rect 12696 27226 12752 27228
rect 12776 27226 12832 27228
rect 12856 27226 12912 27228
rect 12616 27174 12662 27226
rect 12662 27174 12672 27226
rect 12696 27174 12726 27226
rect 12726 27174 12738 27226
rect 12738 27174 12752 27226
rect 12776 27174 12790 27226
rect 12790 27174 12802 27226
rect 12802 27174 12832 27226
rect 12856 27174 12866 27226
rect 12866 27174 12912 27226
rect 12616 27172 12672 27174
rect 12696 27172 12752 27174
rect 12776 27172 12832 27174
rect 12856 27172 12912 27174
rect 17616 27226 17672 27228
rect 17696 27226 17752 27228
rect 17776 27226 17832 27228
rect 17856 27226 17912 27228
rect 17616 27174 17662 27226
rect 17662 27174 17672 27226
rect 17696 27174 17726 27226
rect 17726 27174 17738 27226
rect 17738 27174 17752 27226
rect 17776 27174 17790 27226
rect 17790 27174 17802 27226
rect 17802 27174 17832 27226
rect 17856 27174 17866 27226
rect 17866 27174 17912 27226
rect 17616 27172 17672 27174
rect 17696 27172 17752 27174
rect 17776 27172 17832 27174
rect 17856 27172 17912 27174
rect 22616 27226 22672 27228
rect 22696 27226 22752 27228
rect 22776 27226 22832 27228
rect 22856 27226 22912 27228
rect 22616 27174 22662 27226
rect 22662 27174 22672 27226
rect 22696 27174 22726 27226
rect 22726 27174 22738 27226
rect 22738 27174 22752 27226
rect 22776 27174 22790 27226
rect 22790 27174 22802 27226
rect 22802 27174 22832 27226
rect 22856 27174 22866 27226
rect 22866 27174 22912 27226
rect 22616 27172 22672 27174
rect 22696 27172 22752 27174
rect 22776 27172 22832 27174
rect 22856 27172 22912 27174
rect 27616 27226 27672 27228
rect 27696 27226 27752 27228
rect 27776 27226 27832 27228
rect 27856 27226 27912 27228
rect 27616 27174 27662 27226
rect 27662 27174 27672 27226
rect 27696 27174 27726 27226
rect 27726 27174 27738 27226
rect 27738 27174 27752 27226
rect 27776 27174 27790 27226
rect 27790 27174 27802 27226
rect 27802 27174 27832 27226
rect 27856 27174 27866 27226
rect 27866 27174 27912 27226
rect 27616 27172 27672 27174
rect 27696 27172 27752 27174
rect 27776 27172 27832 27174
rect 27856 27172 27912 27174
rect 32616 27226 32672 27228
rect 32696 27226 32752 27228
rect 32776 27226 32832 27228
rect 32856 27226 32912 27228
rect 32616 27174 32662 27226
rect 32662 27174 32672 27226
rect 32696 27174 32726 27226
rect 32726 27174 32738 27226
rect 32738 27174 32752 27226
rect 32776 27174 32790 27226
rect 32790 27174 32802 27226
rect 32802 27174 32832 27226
rect 32856 27174 32866 27226
rect 32866 27174 32912 27226
rect 32616 27172 32672 27174
rect 32696 27172 32752 27174
rect 32776 27172 32832 27174
rect 32856 27172 32912 27174
rect 37616 27226 37672 27228
rect 37696 27226 37752 27228
rect 37776 27226 37832 27228
rect 37856 27226 37912 27228
rect 37616 27174 37662 27226
rect 37662 27174 37672 27226
rect 37696 27174 37726 27226
rect 37726 27174 37738 27226
rect 37738 27174 37752 27226
rect 37776 27174 37790 27226
rect 37790 27174 37802 27226
rect 37802 27174 37832 27226
rect 37856 27174 37866 27226
rect 37866 27174 37912 27226
rect 37616 27172 37672 27174
rect 37696 27172 37752 27174
rect 37776 27172 37832 27174
rect 37856 27172 37912 27174
rect 42616 27226 42672 27228
rect 42696 27226 42752 27228
rect 42776 27226 42832 27228
rect 42856 27226 42912 27228
rect 42616 27174 42662 27226
rect 42662 27174 42672 27226
rect 42696 27174 42726 27226
rect 42726 27174 42738 27226
rect 42738 27174 42752 27226
rect 42776 27174 42790 27226
rect 42790 27174 42802 27226
rect 42802 27174 42832 27226
rect 42856 27174 42866 27226
rect 42866 27174 42912 27226
rect 42616 27172 42672 27174
rect 42696 27172 42752 27174
rect 42776 27172 42832 27174
rect 42856 27172 42912 27174
rect 47616 27226 47672 27228
rect 47696 27226 47752 27228
rect 47776 27226 47832 27228
rect 47856 27226 47912 27228
rect 47616 27174 47662 27226
rect 47662 27174 47672 27226
rect 47696 27174 47726 27226
rect 47726 27174 47738 27226
rect 47738 27174 47752 27226
rect 47776 27174 47790 27226
rect 47790 27174 47802 27226
rect 47802 27174 47832 27226
rect 47856 27174 47866 27226
rect 47866 27174 47912 27226
rect 47616 27172 47672 27174
rect 47696 27172 47752 27174
rect 47776 27172 47832 27174
rect 47856 27172 47912 27174
rect 52616 27226 52672 27228
rect 52696 27226 52752 27228
rect 52776 27226 52832 27228
rect 52856 27226 52912 27228
rect 52616 27174 52662 27226
rect 52662 27174 52672 27226
rect 52696 27174 52726 27226
rect 52726 27174 52738 27226
rect 52738 27174 52752 27226
rect 52776 27174 52790 27226
rect 52790 27174 52802 27226
rect 52802 27174 52832 27226
rect 52856 27174 52866 27226
rect 52866 27174 52912 27226
rect 52616 27172 52672 27174
rect 52696 27172 52752 27174
rect 52776 27172 52832 27174
rect 52856 27172 52912 27174
rect 57616 27226 57672 27228
rect 57696 27226 57752 27228
rect 57776 27226 57832 27228
rect 57856 27226 57912 27228
rect 57616 27174 57662 27226
rect 57662 27174 57672 27226
rect 57696 27174 57726 27226
rect 57726 27174 57738 27226
rect 57738 27174 57752 27226
rect 57776 27174 57790 27226
rect 57790 27174 57802 27226
rect 57802 27174 57832 27226
rect 57856 27174 57866 27226
rect 57866 27174 57912 27226
rect 57616 27172 57672 27174
rect 57696 27172 57752 27174
rect 57776 27172 57832 27174
rect 57856 27172 57912 27174
rect 58530 26968 58586 27024
rect 1956 26682 2012 26684
rect 2036 26682 2092 26684
rect 2116 26682 2172 26684
rect 2196 26682 2252 26684
rect 1956 26630 2002 26682
rect 2002 26630 2012 26682
rect 2036 26630 2066 26682
rect 2066 26630 2078 26682
rect 2078 26630 2092 26682
rect 2116 26630 2130 26682
rect 2130 26630 2142 26682
rect 2142 26630 2172 26682
rect 2196 26630 2206 26682
rect 2206 26630 2252 26682
rect 1956 26628 2012 26630
rect 2036 26628 2092 26630
rect 2116 26628 2172 26630
rect 2196 26628 2252 26630
rect 6956 26682 7012 26684
rect 7036 26682 7092 26684
rect 7116 26682 7172 26684
rect 7196 26682 7252 26684
rect 6956 26630 7002 26682
rect 7002 26630 7012 26682
rect 7036 26630 7066 26682
rect 7066 26630 7078 26682
rect 7078 26630 7092 26682
rect 7116 26630 7130 26682
rect 7130 26630 7142 26682
rect 7142 26630 7172 26682
rect 7196 26630 7206 26682
rect 7206 26630 7252 26682
rect 6956 26628 7012 26630
rect 7036 26628 7092 26630
rect 7116 26628 7172 26630
rect 7196 26628 7252 26630
rect 11956 26682 12012 26684
rect 12036 26682 12092 26684
rect 12116 26682 12172 26684
rect 12196 26682 12252 26684
rect 11956 26630 12002 26682
rect 12002 26630 12012 26682
rect 12036 26630 12066 26682
rect 12066 26630 12078 26682
rect 12078 26630 12092 26682
rect 12116 26630 12130 26682
rect 12130 26630 12142 26682
rect 12142 26630 12172 26682
rect 12196 26630 12206 26682
rect 12206 26630 12252 26682
rect 11956 26628 12012 26630
rect 12036 26628 12092 26630
rect 12116 26628 12172 26630
rect 12196 26628 12252 26630
rect 16956 26682 17012 26684
rect 17036 26682 17092 26684
rect 17116 26682 17172 26684
rect 17196 26682 17252 26684
rect 16956 26630 17002 26682
rect 17002 26630 17012 26682
rect 17036 26630 17066 26682
rect 17066 26630 17078 26682
rect 17078 26630 17092 26682
rect 17116 26630 17130 26682
rect 17130 26630 17142 26682
rect 17142 26630 17172 26682
rect 17196 26630 17206 26682
rect 17206 26630 17252 26682
rect 16956 26628 17012 26630
rect 17036 26628 17092 26630
rect 17116 26628 17172 26630
rect 17196 26628 17252 26630
rect 21956 26682 22012 26684
rect 22036 26682 22092 26684
rect 22116 26682 22172 26684
rect 22196 26682 22252 26684
rect 21956 26630 22002 26682
rect 22002 26630 22012 26682
rect 22036 26630 22066 26682
rect 22066 26630 22078 26682
rect 22078 26630 22092 26682
rect 22116 26630 22130 26682
rect 22130 26630 22142 26682
rect 22142 26630 22172 26682
rect 22196 26630 22206 26682
rect 22206 26630 22252 26682
rect 21956 26628 22012 26630
rect 22036 26628 22092 26630
rect 22116 26628 22172 26630
rect 22196 26628 22252 26630
rect 26956 26682 27012 26684
rect 27036 26682 27092 26684
rect 27116 26682 27172 26684
rect 27196 26682 27252 26684
rect 26956 26630 27002 26682
rect 27002 26630 27012 26682
rect 27036 26630 27066 26682
rect 27066 26630 27078 26682
rect 27078 26630 27092 26682
rect 27116 26630 27130 26682
rect 27130 26630 27142 26682
rect 27142 26630 27172 26682
rect 27196 26630 27206 26682
rect 27206 26630 27252 26682
rect 26956 26628 27012 26630
rect 27036 26628 27092 26630
rect 27116 26628 27172 26630
rect 27196 26628 27252 26630
rect 31956 26682 32012 26684
rect 32036 26682 32092 26684
rect 32116 26682 32172 26684
rect 32196 26682 32252 26684
rect 31956 26630 32002 26682
rect 32002 26630 32012 26682
rect 32036 26630 32066 26682
rect 32066 26630 32078 26682
rect 32078 26630 32092 26682
rect 32116 26630 32130 26682
rect 32130 26630 32142 26682
rect 32142 26630 32172 26682
rect 32196 26630 32206 26682
rect 32206 26630 32252 26682
rect 31956 26628 32012 26630
rect 32036 26628 32092 26630
rect 32116 26628 32172 26630
rect 32196 26628 32252 26630
rect 36956 26682 37012 26684
rect 37036 26682 37092 26684
rect 37116 26682 37172 26684
rect 37196 26682 37252 26684
rect 36956 26630 37002 26682
rect 37002 26630 37012 26682
rect 37036 26630 37066 26682
rect 37066 26630 37078 26682
rect 37078 26630 37092 26682
rect 37116 26630 37130 26682
rect 37130 26630 37142 26682
rect 37142 26630 37172 26682
rect 37196 26630 37206 26682
rect 37206 26630 37252 26682
rect 36956 26628 37012 26630
rect 37036 26628 37092 26630
rect 37116 26628 37172 26630
rect 37196 26628 37252 26630
rect 41956 26682 42012 26684
rect 42036 26682 42092 26684
rect 42116 26682 42172 26684
rect 42196 26682 42252 26684
rect 41956 26630 42002 26682
rect 42002 26630 42012 26682
rect 42036 26630 42066 26682
rect 42066 26630 42078 26682
rect 42078 26630 42092 26682
rect 42116 26630 42130 26682
rect 42130 26630 42142 26682
rect 42142 26630 42172 26682
rect 42196 26630 42206 26682
rect 42206 26630 42252 26682
rect 41956 26628 42012 26630
rect 42036 26628 42092 26630
rect 42116 26628 42172 26630
rect 42196 26628 42252 26630
rect 46956 26682 47012 26684
rect 47036 26682 47092 26684
rect 47116 26682 47172 26684
rect 47196 26682 47252 26684
rect 46956 26630 47002 26682
rect 47002 26630 47012 26682
rect 47036 26630 47066 26682
rect 47066 26630 47078 26682
rect 47078 26630 47092 26682
rect 47116 26630 47130 26682
rect 47130 26630 47142 26682
rect 47142 26630 47172 26682
rect 47196 26630 47206 26682
rect 47206 26630 47252 26682
rect 46956 26628 47012 26630
rect 47036 26628 47092 26630
rect 47116 26628 47172 26630
rect 47196 26628 47252 26630
rect 51956 26682 52012 26684
rect 52036 26682 52092 26684
rect 52116 26682 52172 26684
rect 52196 26682 52252 26684
rect 51956 26630 52002 26682
rect 52002 26630 52012 26682
rect 52036 26630 52066 26682
rect 52066 26630 52078 26682
rect 52078 26630 52092 26682
rect 52116 26630 52130 26682
rect 52130 26630 52142 26682
rect 52142 26630 52172 26682
rect 52196 26630 52206 26682
rect 52206 26630 52252 26682
rect 51956 26628 52012 26630
rect 52036 26628 52092 26630
rect 52116 26628 52172 26630
rect 52196 26628 52252 26630
rect 56956 26682 57012 26684
rect 57036 26682 57092 26684
rect 57116 26682 57172 26684
rect 57196 26682 57252 26684
rect 56956 26630 57002 26682
rect 57002 26630 57012 26682
rect 57036 26630 57066 26682
rect 57066 26630 57078 26682
rect 57078 26630 57092 26682
rect 57116 26630 57130 26682
rect 57130 26630 57142 26682
rect 57142 26630 57172 26682
rect 57196 26630 57206 26682
rect 57206 26630 57252 26682
rect 56956 26628 57012 26630
rect 57036 26628 57092 26630
rect 57116 26628 57172 26630
rect 57196 26628 57252 26630
rect 58346 26152 58402 26208
rect 2616 26138 2672 26140
rect 2696 26138 2752 26140
rect 2776 26138 2832 26140
rect 2856 26138 2912 26140
rect 2616 26086 2662 26138
rect 2662 26086 2672 26138
rect 2696 26086 2726 26138
rect 2726 26086 2738 26138
rect 2738 26086 2752 26138
rect 2776 26086 2790 26138
rect 2790 26086 2802 26138
rect 2802 26086 2832 26138
rect 2856 26086 2866 26138
rect 2866 26086 2912 26138
rect 2616 26084 2672 26086
rect 2696 26084 2752 26086
rect 2776 26084 2832 26086
rect 2856 26084 2912 26086
rect 7616 26138 7672 26140
rect 7696 26138 7752 26140
rect 7776 26138 7832 26140
rect 7856 26138 7912 26140
rect 7616 26086 7662 26138
rect 7662 26086 7672 26138
rect 7696 26086 7726 26138
rect 7726 26086 7738 26138
rect 7738 26086 7752 26138
rect 7776 26086 7790 26138
rect 7790 26086 7802 26138
rect 7802 26086 7832 26138
rect 7856 26086 7866 26138
rect 7866 26086 7912 26138
rect 7616 26084 7672 26086
rect 7696 26084 7752 26086
rect 7776 26084 7832 26086
rect 7856 26084 7912 26086
rect 12616 26138 12672 26140
rect 12696 26138 12752 26140
rect 12776 26138 12832 26140
rect 12856 26138 12912 26140
rect 12616 26086 12662 26138
rect 12662 26086 12672 26138
rect 12696 26086 12726 26138
rect 12726 26086 12738 26138
rect 12738 26086 12752 26138
rect 12776 26086 12790 26138
rect 12790 26086 12802 26138
rect 12802 26086 12832 26138
rect 12856 26086 12866 26138
rect 12866 26086 12912 26138
rect 12616 26084 12672 26086
rect 12696 26084 12752 26086
rect 12776 26084 12832 26086
rect 12856 26084 12912 26086
rect 17616 26138 17672 26140
rect 17696 26138 17752 26140
rect 17776 26138 17832 26140
rect 17856 26138 17912 26140
rect 17616 26086 17662 26138
rect 17662 26086 17672 26138
rect 17696 26086 17726 26138
rect 17726 26086 17738 26138
rect 17738 26086 17752 26138
rect 17776 26086 17790 26138
rect 17790 26086 17802 26138
rect 17802 26086 17832 26138
rect 17856 26086 17866 26138
rect 17866 26086 17912 26138
rect 17616 26084 17672 26086
rect 17696 26084 17752 26086
rect 17776 26084 17832 26086
rect 17856 26084 17912 26086
rect 22616 26138 22672 26140
rect 22696 26138 22752 26140
rect 22776 26138 22832 26140
rect 22856 26138 22912 26140
rect 22616 26086 22662 26138
rect 22662 26086 22672 26138
rect 22696 26086 22726 26138
rect 22726 26086 22738 26138
rect 22738 26086 22752 26138
rect 22776 26086 22790 26138
rect 22790 26086 22802 26138
rect 22802 26086 22832 26138
rect 22856 26086 22866 26138
rect 22866 26086 22912 26138
rect 22616 26084 22672 26086
rect 22696 26084 22752 26086
rect 22776 26084 22832 26086
rect 22856 26084 22912 26086
rect 27616 26138 27672 26140
rect 27696 26138 27752 26140
rect 27776 26138 27832 26140
rect 27856 26138 27912 26140
rect 27616 26086 27662 26138
rect 27662 26086 27672 26138
rect 27696 26086 27726 26138
rect 27726 26086 27738 26138
rect 27738 26086 27752 26138
rect 27776 26086 27790 26138
rect 27790 26086 27802 26138
rect 27802 26086 27832 26138
rect 27856 26086 27866 26138
rect 27866 26086 27912 26138
rect 27616 26084 27672 26086
rect 27696 26084 27752 26086
rect 27776 26084 27832 26086
rect 27856 26084 27912 26086
rect 32616 26138 32672 26140
rect 32696 26138 32752 26140
rect 32776 26138 32832 26140
rect 32856 26138 32912 26140
rect 32616 26086 32662 26138
rect 32662 26086 32672 26138
rect 32696 26086 32726 26138
rect 32726 26086 32738 26138
rect 32738 26086 32752 26138
rect 32776 26086 32790 26138
rect 32790 26086 32802 26138
rect 32802 26086 32832 26138
rect 32856 26086 32866 26138
rect 32866 26086 32912 26138
rect 32616 26084 32672 26086
rect 32696 26084 32752 26086
rect 32776 26084 32832 26086
rect 32856 26084 32912 26086
rect 37616 26138 37672 26140
rect 37696 26138 37752 26140
rect 37776 26138 37832 26140
rect 37856 26138 37912 26140
rect 37616 26086 37662 26138
rect 37662 26086 37672 26138
rect 37696 26086 37726 26138
rect 37726 26086 37738 26138
rect 37738 26086 37752 26138
rect 37776 26086 37790 26138
rect 37790 26086 37802 26138
rect 37802 26086 37832 26138
rect 37856 26086 37866 26138
rect 37866 26086 37912 26138
rect 37616 26084 37672 26086
rect 37696 26084 37752 26086
rect 37776 26084 37832 26086
rect 37856 26084 37912 26086
rect 42616 26138 42672 26140
rect 42696 26138 42752 26140
rect 42776 26138 42832 26140
rect 42856 26138 42912 26140
rect 42616 26086 42662 26138
rect 42662 26086 42672 26138
rect 42696 26086 42726 26138
rect 42726 26086 42738 26138
rect 42738 26086 42752 26138
rect 42776 26086 42790 26138
rect 42790 26086 42802 26138
rect 42802 26086 42832 26138
rect 42856 26086 42866 26138
rect 42866 26086 42912 26138
rect 42616 26084 42672 26086
rect 42696 26084 42752 26086
rect 42776 26084 42832 26086
rect 42856 26084 42912 26086
rect 47616 26138 47672 26140
rect 47696 26138 47752 26140
rect 47776 26138 47832 26140
rect 47856 26138 47912 26140
rect 47616 26086 47662 26138
rect 47662 26086 47672 26138
rect 47696 26086 47726 26138
rect 47726 26086 47738 26138
rect 47738 26086 47752 26138
rect 47776 26086 47790 26138
rect 47790 26086 47802 26138
rect 47802 26086 47832 26138
rect 47856 26086 47866 26138
rect 47866 26086 47912 26138
rect 47616 26084 47672 26086
rect 47696 26084 47752 26086
rect 47776 26084 47832 26086
rect 47856 26084 47912 26086
rect 52616 26138 52672 26140
rect 52696 26138 52752 26140
rect 52776 26138 52832 26140
rect 52856 26138 52912 26140
rect 52616 26086 52662 26138
rect 52662 26086 52672 26138
rect 52696 26086 52726 26138
rect 52726 26086 52738 26138
rect 52738 26086 52752 26138
rect 52776 26086 52790 26138
rect 52790 26086 52802 26138
rect 52802 26086 52832 26138
rect 52856 26086 52866 26138
rect 52866 26086 52912 26138
rect 52616 26084 52672 26086
rect 52696 26084 52752 26086
rect 52776 26084 52832 26086
rect 52856 26084 52912 26086
rect 57616 26138 57672 26140
rect 57696 26138 57752 26140
rect 57776 26138 57832 26140
rect 57856 26138 57912 26140
rect 57616 26086 57662 26138
rect 57662 26086 57672 26138
rect 57696 26086 57726 26138
rect 57726 26086 57738 26138
rect 57738 26086 57752 26138
rect 57776 26086 57790 26138
rect 57790 26086 57802 26138
rect 57802 26086 57832 26138
rect 57856 26086 57866 26138
rect 57866 26086 57912 26138
rect 57616 26084 57672 26086
rect 57696 26084 57752 26086
rect 57776 26084 57832 26086
rect 57856 26084 57912 26086
rect 1956 25594 2012 25596
rect 2036 25594 2092 25596
rect 2116 25594 2172 25596
rect 2196 25594 2252 25596
rect 1956 25542 2002 25594
rect 2002 25542 2012 25594
rect 2036 25542 2066 25594
rect 2066 25542 2078 25594
rect 2078 25542 2092 25594
rect 2116 25542 2130 25594
rect 2130 25542 2142 25594
rect 2142 25542 2172 25594
rect 2196 25542 2206 25594
rect 2206 25542 2252 25594
rect 1956 25540 2012 25542
rect 2036 25540 2092 25542
rect 2116 25540 2172 25542
rect 2196 25540 2252 25542
rect 6956 25594 7012 25596
rect 7036 25594 7092 25596
rect 7116 25594 7172 25596
rect 7196 25594 7252 25596
rect 6956 25542 7002 25594
rect 7002 25542 7012 25594
rect 7036 25542 7066 25594
rect 7066 25542 7078 25594
rect 7078 25542 7092 25594
rect 7116 25542 7130 25594
rect 7130 25542 7142 25594
rect 7142 25542 7172 25594
rect 7196 25542 7206 25594
rect 7206 25542 7252 25594
rect 6956 25540 7012 25542
rect 7036 25540 7092 25542
rect 7116 25540 7172 25542
rect 7196 25540 7252 25542
rect 11956 25594 12012 25596
rect 12036 25594 12092 25596
rect 12116 25594 12172 25596
rect 12196 25594 12252 25596
rect 11956 25542 12002 25594
rect 12002 25542 12012 25594
rect 12036 25542 12066 25594
rect 12066 25542 12078 25594
rect 12078 25542 12092 25594
rect 12116 25542 12130 25594
rect 12130 25542 12142 25594
rect 12142 25542 12172 25594
rect 12196 25542 12206 25594
rect 12206 25542 12252 25594
rect 11956 25540 12012 25542
rect 12036 25540 12092 25542
rect 12116 25540 12172 25542
rect 12196 25540 12252 25542
rect 16956 25594 17012 25596
rect 17036 25594 17092 25596
rect 17116 25594 17172 25596
rect 17196 25594 17252 25596
rect 16956 25542 17002 25594
rect 17002 25542 17012 25594
rect 17036 25542 17066 25594
rect 17066 25542 17078 25594
rect 17078 25542 17092 25594
rect 17116 25542 17130 25594
rect 17130 25542 17142 25594
rect 17142 25542 17172 25594
rect 17196 25542 17206 25594
rect 17206 25542 17252 25594
rect 16956 25540 17012 25542
rect 17036 25540 17092 25542
rect 17116 25540 17172 25542
rect 17196 25540 17252 25542
rect 21956 25594 22012 25596
rect 22036 25594 22092 25596
rect 22116 25594 22172 25596
rect 22196 25594 22252 25596
rect 21956 25542 22002 25594
rect 22002 25542 22012 25594
rect 22036 25542 22066 25594
rect 22066 25542 22078 25594
rect 22078 25542 22092 25594
rect 22116 25542 22130 25594
rect 22130 25542 22142 25594
rect 22142 25542 22172 25594
rect 22196 25542 22206 25594
rect 22206 25542 22252 25594
rect 21956 25540 22012 25542
rect 22036 25540 22092 25542
rect 22116 25540 22172 25542
rect 22196 25540 22252 25542
rect 26956 25594 27012 25596
rect 27036 25594 27092 25596
rect 27116 25594 27172 25596
rect 27196 25594 27252 25596
rect 26956 25542 27002 25594
rect 27002 25542 27012 25594
rect 27036 25542 27066 25594
rect 27066 25542 27078 25594
rect 27078 25542 27092 25594
rect 27116 25542 27130 25594
rect 27130 25542 27142 25594
rect 27142 25542 27172 25594
rect 27196 25542 27206 25594
rect 27206 25542 27252 25594
rect 26956 25540 27012 25542
rect 27036 25540 27092 25542
rect 27116 25540 27172 25542
rect 27196 25540 27252 25542
rect 31956 25594 32012 25596
rect 32036 25594 32092 25596
rect 32116 25594 32172 25596
rect 32196 25594 32252 25596
rect 31956 25542 32002 25594
rect 32002 25542 32012 25594
rect 32036 25542 32066 25594
rect 32066 25542 32078 25594
rect 32078 25542 32092 25594
rect 32116 25542 32130 25594
rect 32130 25542 32142 25594
rect 32142 25542 32172 25594
rect 32196 25542 32206 25594
rect 32206 25542 32252 25594
rect 31956 25540 32012 25542
rect 32036 25540 32092 25542
rect 32116 25540 32172 25542
rect 32196 25540 32252 25542
rect 36956 25594 37012 25596
rect 37036 25594 37092 25596
rect 37116 25594 37172 25596
rect 37196 25594 37252 25596
rect 36956 25542 37002 25594
rect 37002 25542 37012 25594
rect 37036 25542 37066 25594
rect 37066 25542 37078 25594
rect 37078 25542 37092 25594
rect 37116 25542 37130 25594
rect 37130 25542 37142 25594
rect 37142 25542 37172 25594
rect 37196 25542 37206 25594
rect 37206 25542 37252 25594
rect 36956 25540 37012 25542
rect 37036 25540 37092 25542
rect 37116 25540 37172 25542
rect 37196 25540 37252 25542
rect 41956 25594 42012 25596
rect 42036 25594 42092 25596
rect 42116 25594 42172 25596
rect 42196 25594 42252 25596
rect 41956 25542 42002 25594
rect 42002 25542 42012 25594
rect 42036 25542 42066 25594
rect 42066 25542 42078 25594
rect 42078 25542 42092 25594
rect 42116 25542 42130 25594
rect 42130 25542 42142 25594
rect 42142 25542 42172 25594
rect 42196 25542 42206 25594
rect 42206 25542 42252 25594
rect 41956 25540 42012 25542
rect 42036 25540 42092 25542
rect 42116 25540 42172 25542
rect 42196 25540 42252 25542
rect 46956 25594 47012 25596
rect 47036 25594 47092 25596
rect 47116 25594 47172 25596
rect 47196 25594 47252 25596
rect 46956 25542 47002 25594
rect 47002 25542 47012 25594
rect 47036 25542 47066 25594
rect 47066 25542 47078 25594
rect 47078 25542 47092 25594
rect 47116 25542 47130 25594
rect 47130 25542 47142 25594
rect 47142 25542 47172 25594
rect 47196 25542 47206 25594
rect 47206 25542 47252 25594
rect 46956 25540 47012 25542
rect 47036 25540 47092 25542
rect 47116 25540 47172 25542
rect 47196 25540 47252 25542
rect 51956 25594 52012 25596
rect 52036 25594 52092 25596
rect 52116 25594 52172 25596
rect 52196 25594 52252 25596
rect 51956 25542 52002 25594
rect 52002 25542 52012 25594
rect 52036 25542 52066 25594
rect 52066 25542 52078 25594
rect 52078 25542 52092 25594
rect 52116 25542 52130 25594
rect 52130 25542 52142 25594
rect 52142 25542 52172 25594
rect 52196 25542 52206 25594
rect 52206 25542 52252 25594
rect 51956 25540 52012 25542
rect 52036 25540 52092 25542
rect 52116 25540 52172 25542
rect 52196 25540 52252 25542
rect 56956 25594 57012 25596
rect 57036 25594 57092 25596
rect 57116 25594 57172 25596
rect 57196 25594 57252 25596
rect 56956 25542 57002 25594
rect 57002 25542 57012 25594
rect 57036 25542 57066 25594
rect 57066 25542 57078 25594
rect 57078 25542 57092 25594
rect 57116 25542 57130 25594
rect 57130 25542 57142 25594
rect 57142 25542 57172 25594
rect 57196 25542 57206 25594
rect 57206 25542 57252 25594
rect 56956 25540 57012 25542
rect 57036 25540 57092 25542
rect 57116 25540 57172 25542
rect 57196 25540 57252 25542
rect 58530 25336 58586 25392
rect 2616 25050 2672 25052
rect 2696 25050 2752 25052
rect 2776 25050 2832 25052
rect 2856 25050 2912 25052
rect 2616 24998 2662 25050
rect 2662 24998 2672 25050
rect 2696 24998 2726 25050
rect 2726 24998 2738 25050
rect 2738 24998 2752 25050
rect 2776 24998 2790 25050
rect 2790 24998 2802 25050
rect 2802 24998 2832 25050
rect 2856 24998 2866 25050
rect 2866 24998 2912 25050
rect 2616 24996 2672 24998
rect 2696 24996 2752 24998
rect 2776 24996 2832 24998
rect 2856 24996 2912 24998
rect 7616 25050 7672 25052
rect 7696 25050 7752 25052
rect 7776 25050 7832 25052
rect 7856 25050 7912 25052
rect 7616 24998 7662 25050
rect 7662 24998 7672 25050
rect 7696 24998 7726 25050
rect 7726 24998 7738 25050
rect 7738 24998 7752 25050
rect 7776 24998 7790 25050
rect 7790 24998 7802 25050
rect 7802 24998 7832 25050
rect 7856 24998 7866 25050
rect 7866 24998 7912 25050
rect 7616 24996 7672 24998
rect 7696 24996 7752 24998
rect 7776 24996 7832 24998
rect 7856 24996 7912 24998
rect 12616 25050 12672 25052
rect 12696 25050 12752 25052
rect 12776 25050 12832 25052
rect 12856 25050 12912 25052
rect 12616 24998 12662 25050
rect 12662 24998 12672 25050
rect 12696 24998 12726 25050
rect 12726 24998 12738 25050
rect 12738 24998 12752 25050
rect 12776 24998 12790 25050
rect 12790 24998 12802 25050
rect 12802 24998 12832 25050
rect 12856 24998 12866 25050
rect 12866 24998 12912 25050
rect 12616 24996 12672 24998
rect 12696 24996 12752 24998
rect 12776 24996 12832 24998
rect 12856 24996 12912 24998
rect 17616 25050 17672 25052
rect 17696 25050 17752 25052
rect 17776 25050 17832 25052
rect 17856 25050 17912 25052
rect 17616 24998 17662 25050
rect 17662 24998 17672 25050
rect 17696 24998 17726 25050
rect 17726 24998 17738 25050
rect 17738 24998 17752 25050
rect 17776 24998 17790 25050
rect 17790 24998 17802 25050
rect 17802 24998 17832 25050
rect 17856 24998 17866 25050
rect 17866 24998 17912 25050
rect 17616 24996 17672 24998
rect 17696 24996 17752 24998
rect 17776 24996 17832 24998
rect 17856 24996 17912 24998
rect 22616 25050 22672 25052
rect 22696 25050 22752 25052
rect 22776 25050 22832 25052
rect 22856 25050 22912 25052
rect 22616 24998 22662 25050
rect 22662 24998 22672 25050
rect 22696 24998 22726 25050
rect 22726 24998 22738 25050
rect 22738 24998 22752 25050
rect 22776 24998 22790 25050
rect 22790 24998 22802 25050
rect 22802 24998 22832 25050
rect 22856 24998 22866 25050
rect 22866 24998 22912 25050
rect 22616 24996 22672 24998
rect 22696 24996 22752 24998
rect 22776 24996 22832 24998
rect 22856 24996 22912 24998
rect 27616 25050 27672 25052
rect 27696 25050 27752 25052
rect 27776 25050 27832 25052
rect 27856 25050 27912 25052
rect 27616 24998 27662 25050
rect 27662 24998 27672 25050
rect 27696 24998 27726 25050
rect 27726 24998 27738 25050
rect 27738 24998 27752 25050
rect 27776 24998 27790 25050
rect 27790 24998 27802 25050
rect 27802 24998 27832 25050
rect 27856 24998 27866 25050
rect 27866 24998 27912 25050
rect 27616 24996 27672 24998
rect 27696 24996 27752 24998
rect 27776 24996 27832 24998
rect 27856 24996 27912 24998
rect 32616 25050 32672 25052
rect 32696 25050 32752 25052
rect 32776 25050 32832 25052
rect 32856 25050 32912 25052
rect 32616 24998 32662 25050
rect 32662 24998 32672 25050
rect 32696 24998 32726 25050
rect 32726 24998 32738 25050
rect 32738 24998 32752 25050
rect 32776 24998 32790 25050
rect 32790 24998 32802 25050
rect 32802 24998 32832 25050
rect 32856 24998 32866 25050
rect 32866 24998 32912 25050
rect 32616 24996 32672 24998
rect 32696 24996 32752 24998
rect 32776 24996 32832 24998
rect 32856 24996 32912 24998
rect 37616 25050 37672 25052
rect 37696 25050 37752 25052
rect 37776 25050 37832 25052
rect 37856 25050 37912 25052
rect 37616 24998 37662 25050
rect 37662 24998 37672 25050
rect 37696 24998 37726 25050
rect 37726 24998 37738 25050
rect 37738 24998 37752 25050
rect 37776 24998 37790 25050
rect 37790 24998 37802 25050
rect 37802 24998 37832 25050
rect 37856 24998 37866 25050
rect 37866 24998 37912 25050
rect 37616 24996 37672 24998
rect 37696 24996 37752 24998
rect 37776 24996 37832 24998
rect 37856 24996 37912 24998
rect 42616 25050 42672 25052
rect 42696 25050 42752 25052
rect 42776 25050 42832 25052
rect 42856 25050 42912 25052
rect 42616 24998 42662 25050
rect 42662 24998 42672 25050
rect 42696 24998 42726 25050
rect 42726 24998 42738 25050
rect 42738 24998 42752 25050
rect 42776 24998 42790 25050
rect 42790 24998 42802 25050
rect 42802 24998 42832 25050
rect 42856 24998 42866 25050
rect 42866 24998 42912 25050
rect 42616 24996 42672 24998
rect 42696 24996 42752 24998
rect 42776 24996 42832 24998
rect 42856 24996 42912 24998
rect 47616 25050 47672 25052
rect 47696 25050 47752 25052
rect 47776 25050 47832 25052
rect 47856 25050 47912 25052
rect 47616 24998 47662 25050
rect 47662 24998 47672 25050
rect 47696 24998 47726 25050
rect 47726 24998 47738 25050
rect 47738 24998 47752 25050
rect 47776 24998 47790 25050
rect 47790 24998 47802 25050
rect 47802 24998 47832 25050
rect 47856 24998 47866 25050
rect 47866 24998 47912 25050
rect 47616 24996 47672 24998
rect 47696 24996 47752 24998
rect 47776 24996 47832 24998
rect 47856 24996 47912 24998
rect 52616 25050 52672 25052
rect 52696 25050 52752 25052
rect 52776 25050 52832 25052
rect 52856 25050 52912 25052
rect 52616 24998 52662 25050
rect 52662 24998 52672 25050
rect 52696 24998 52726 25050
rect 52726 24998 52738 25050
rect 52738 24998 52752 25050
rect 52776 24998 52790 25050
rect 52790 24998 52802 25050
rect 52802 24998 52832 25050
rect 52856 24998 52866 25050
rect 52866 24998 52912 25050
rect 52616 24996 52672 24998
rect 52696 24996 52752 24998
rect 52776 24996 52832 24998
rect 52856 24996 52912 24998
rect 57616 25050 57672 25052
rect 57696 25050 57752 25052
rect 57776 25050 57832 25052
rect 57856 25050 57912 25052
rect 57616 24998 57662 25050
rect 57662 24998 57672 25050
rect 57696 24998 57726 25050
rect 57726 24998 57738 25050
rect 57738 24998 57752 25050
rect 57776 24998 57790 25050
rect 57790 24998 57802 25050
rect 57802 24998 57832 25050
rect 57856 24998 57866 25050
rect 57866 24998 57912 25050
rect 57616 24996 57672 24998
rect 57696 24996 57752 24998
rect 57776 24996 57832 24998
rect 57856 24996 57912 24998
rect 58530 24556 58532 24576
rect 58532 24556 58584 24576
rect 58584 24556 58586 24576
rect 58530 24520 58586 24556
rect 1956 24506 2012 24508
rect 2036 24506 2092 24508
rect 2116 24506 2172 24508
rect 2196 24506 2252 24508
rect 1956 24454 2002 24506
rect 2002 24454 2012 24506
rect 2036 24454 2066 24506
rect 2066 24454 2078 24506
rect 2078 24454 2092 24506
rect 2116 24454 2130 24506
rect 2130 24454 2142 24506
rect 2142 24454 2172 24506
rect 2196 24454 2206 24506
rect 2206 24454 2252 24506
rect 1956 24452 2012 24454
rect 2036 24452 2092 24454
rect 2116 24452 2172 24454
rect 2196 24452 2252 24454
rect 6956 24506 7012 24508
rect 7036 24506 7092 24508
rect 7116 24506 7172 24508
rect 7196 24506 7252 24508
rect 6956 24454 7002 24506
rect 7002 24454 7012 24506
rect 7036 24454 7066 24506
rect 7066 24454 7078 24506
rect 7078 24454 7092 24506
rect 7116 24454 7130 24506
rect 7130 24454 7142 24506
rect 7142 24454 7172 24506
rect 7196 24454 7206 24506
rect 7206 24454 7252 24506
rect 6956 24452 7012 24454
rect 7036 24452 7092 24454
rect 7116 24452 7172 24454
rect 7196 24452 7252 24454
rect 11956 24506 12012 24508
rect 12036 24506 12092 24508
rect 12116 24506 12172 24508
rect 12196 24506 12252 24508
rect 11956 24454 12002 24506
rect 12002 24454 12012 24506
rect 12036 24454 12066 24506
rect 12066 24454 12078 24506
rect 12078 24454 12092 24506
rect 12116 24454 12130 24506
rect 12130 24454 12142 24506
rect 12142 24454 12172 24506
rect 12196 24454 12206 24506
rect 12206 24454 12252 24506
rect 11956 24452 12012 24454
rect 12036 24452 12092 24454
rect 12116 24452 12172 24454
rect 12196 24452 12252 24454
rect 16956 24506 17012 24508
rect 17036 24506 17092 24508
rect 17116 24506 17172 24508
rect 17196 24506 17252 24508
rect 16956 24454 17002 24506
rect 17002 24454 17012 24506
rect 17036 24454 17066 24506
rect 17066 24454 17078 24506
rect 17078 24454 17092 24506
rect 17116 24454 17130 24506
rect 17130 24454 17142 24506
rect 17142 24454 17172 24506
rect 17196 24454 17206 24506
rect 17206 24454 17252 24506
rect 16956 24452 17012 24454
rect 17036 24452 17092 24454
rect 17116 24452 17172 24454
rect 17196 24452 17252 24454
rect 21956 24506 22012 24508
rect 22036 24506 22092 24508
rect 22116 24506 22172 24508
rect 22196 24506 22252 24508
rect 21956 24454 22002 24506
rect 22002 24454 22012 24506
rect 22036 24454 22066 24506
rect 22066 24454 22078 24506
rect 22078 24454 22092 24506
rect 22116 24454 22130 24506
rect 22130 24454 22142 24506
rect 22142 24454 22172 24506
rect 22196 24454 22206 24506
rect 22206 24454 22252 24506
rect 21956 24452 22012 24454
rect 22036 24452 22092 24454
rect 22116 24452 22172 24454
rect 22196 24452 22252 24454
rect 26956 24506 27012 24508
rect 27036 24506 27092 24508
rect 27116 24506 27172 24508
rect 27196 24506 27252 24508
rect 26956 24454 27002 24506
rect 27002 24454 27012 24506
rect 27036 24454 27066 24506
rect 27066 24454 27078 24506
rect 27078 24454 27092 24506
rect 27116 24454 27130 24506
rect 27130 24454 27142 24506
rect 27142 24454 27172 24506
rect 27196 24454 27206 24506
rect 27206 24454 27252 24506
rect 26956 24452 27012 24454
rect 27036 24452 27092 24454
rect 27116 24452 27172 24454
rect 27196 24452 27252 24454
rect 31956 24506 32012 24508
rect 32036 24506 32092 24508
rect 32116 24506 32172 24508
rect 32196 24506 32252 24508
rect 31956 24454 32002 24506
rect 32002 24454 32012 24506
rect 32036 24454 32066 24506
rect 32066 24454 32078 24506
rect 32078 24454 32092 24506
rect 32116 24454 32130 24506
rect 32130 24454 32142 24506
rect 32142 24454 32172 24506
rect 32196 24454 32206 24506
rect 32206 24454 32252 24506
rect 31956 24452 32012 24454
rect 32036 24452 32092 24454
rect 32116 24452 32172 24454
rect 32196 24452 32252 24454
rect 36956 24506 37012 24508
rect 37036 24506 37092 24508
rect 37116 24506 37172 24508
rect 37196 24506 37252 24508
rect 36956 24454 37002 24506
rect 37002 24454 37012 24506
rect 37036 24454 37066 24506
rect 37066 24454 37078 24506
rect 37078 24454 37092 24506
rect 37116 24454 37130 24506
rect 37130 24454 37142 24506
rect 37142 24454 37172 24506
rect 37196 24454 37206 24506
rect 37206 24454 37252 24506
rect 36956 24452 37012 24454
rect 37036 24452 37092 24454
rect 37116 24452 37172 24454
rect 37196 24452 37252 24454
rect 41956 24506 42012 24508
rect 42036 24506 42092 24508
rect 42116 24506 42172 24508
rect 42196 24506 42252 24508
rect 41956 24454 42002 24506
rect 42002 24454 42012 24506
rect 42036 24454 42066 24506
rect 42066 24454 42078 24506
rect 42078 24454 42092 24506
rect 42116 24454 42130 24506
rect 42130 24454 42142 24506
rect 42142 24454 42172 24506
rect 42196 24454 42206 24506
rect 42206 24454 42252 24506
rect 41956 24452 42012 24454
rect 42036 24452 42092 24454
rect 42116 24452 42172 24454
rect 42196 24452 42252 24454
rect 46956 24506 47012 24508
rect 47036 24506 47092 24508
rect 47116 24506 47172 24508
rect 47196 24506 47252 24508
rect 46956 24454 47002 24506
rect 47002 24454 47012 24506
rect 47036 24454 47066 24506
rect 47066 24454 47078 24506
rect 47078 24454 47092 24506
rect 47116 24454 47130 24506
rect 47130 24454 47142 24506
rect 47142 24454 47172 24506
rect 47196 24454 47206 24506
rect 47206 24454 47252 24506
rect 46956 24452 47012 24454
rect 47036 24452 47092 24454
rect 47116 24452 47172 24454
rect 47196 24452 47252 24454
rect 51956 24506 52012 24508
rect 52036 24506 52092 24508
rect 52116 24506 52172 24508
rect 52196 24506 52252 24508
rect 51956 24454 52002 24506
rect 52002 24454 52012 24506
rect 52036 24454 52066 24506
rect 52066 24454 52078 24506
rect 52078 24454 52092 24506
rect 52116 24454 52130 24506
rect 52130 24454 52142 24506
rect 52142 24454 52172 24506
rect 52196 24454 52206 24506
rect 52206 24454 52252 24506
rect 51956 24452 52012 24454
rect 52036 24452 52092 24454
rect 52116 24452 52172 24454
rect 52196 24452 52252 24454
rect 56956 24506 57012 24508
rect 57036 24506 57092 24508
rect 57116 24506 57172 24508
rect 57196 24506 57252 24508
rect 56956 24454 57002 24506
rect 57002 24454 57012 24506
rect 57036 24454 57066 24506
rect 57066 24454 57078 24506
rect 57078 24454 57092 24506
rect 57116 24454 57130 24506
rect 57130 24454 57142 24506
rect 57142 24454 57172 24506
rect 57196 24454 57206 24506
rect 57206 24454 57252 24506
rect 56956 24452 57012 24454
rect 57036 24452 57092 24454
rect 57116 24452 57172 24454
rect 57196 24452 57252 24454
rect 2616 23962 2672 23964
rect 2696 23962 2752 23964
rect 2776 23962 2832 23964
rect 2856 23962 2912 23964
rect 2616 23910 2662 23962
rect 2662 23910 2672 23962
rect 2696 23910 2726 23962
rect 2726 23910 2738 23962
rect 2738 23910 2752 23962
rect 2776 23910 2790 23962
rect 2790 23910 2802 23962
rect 2802 23910 2832 23962
rect 2856 23910 2866 23962
rect 2866 23910 2912 23962
rect 2616 23908 2672 23910
rect 2696 23908 2752 23910
rect 2776 23908 2832 23910
rect 2856 23908 2912 23910
rect 7616 23962 7672 23964
rect 7696 23962 7752 23964
rect 7776 23962 7832 23964
rect 7856 23962 7912 23964
rect 7616 23910 7662 23962
rect 7662 23910 7672 23962
rect 7696 23910 7726 23962
rect 7726 23910 7738 23962
rect 7738 23910 7752 23962
rect 7776 23910 7790 23962
rect 7790 23910 7802 23962
rect 7802 23910 7832 23962
rect 7856 23910 7866 23962
rect 7866 23910 7912 23962
rect 7616 23908 7672 23910
rect 7696 23908 7752 23910
rect 7776 23908 7832 23910
rect 7856 23908 7912 23910
rect 12616 23962 12672 23964
rect 12696 23962 12752 23964
rect 12776 23962 12832 23964
rect 12856 23962 12912 23964
rect 12616 23910 12662 23962
rect 12662 23910 12672 23962
rect 12696 23910 12726 23962
rect 12726 23910 12738 23962
rect 12738 23910 12752 23962
rect 12776 23910 12790 23962
rect 12790 23910 12802 23962
rect 12802 23910 12832 23962
rect 12856 23910 12866 23962
rect 12866 23910 12912 23962
rect 12616 23908 12672 23910
rect 12696 23908 12752 23910
rect 12776 23908 12832 23910
rect 12856 23908 12912 23910
rect 17616 23962 17672 23964
rect 17696 23962 17752 23964
rect 17776 23962 17832 23964
rect 17856 23962 17912 23964
rect 17616 23910 17662 23962
rect 17662 23910 17672 23962
rect 17696 23910 17726 23962
rect 17726 23910 17738 23962
rect 17738 23910 17752 23962
rect 17776 23910 17790 23962
rect 17790 23910 17802 23962
rect 17802 23910 17832 23962
rect 17856 23910 17866 23962
rect 17866 23910 17912 23962
rect 17616 23908 17672 23910
rect 17696 23908 17752 23910
rect 17776 23908 17832 23910
rect 17856 23908 17912 23910
rect 22616 23962 22672 23964
rect 22696 23962 22752 23964
rect 22776 23962 22832 23964
rect 22856 23962 22912 23964
rect 22616 23910 22662 23962
rect 22662 23910 22672 23962
rect 22696 23910 22726 23962
rect 22726 23910 22738 23962
rect 22738 23910 22752 23962
rect 22776 23910 22790 23962
rect 22790 23910 22802 23962
rect 22802 23910 22832 23962
rect 22856 23910 22866 23962
rect 22866 23910 22912 23962
rect 22616 23908 22672 23910
rect 22696 23908 22752 23910
rect 22776 23908 22832 23910
rect 22856 23908 22912 23910
rect 27616 23962 27672 23964
rect 27696 23962 27752 23964
rect 27776 23962 27832 23964
rect 27856 23962 27912 23964
rect 27616 23910 27662 23962
rect 27662 23910 27672 23962
rect 27696 23910 27726 23962
rect 27726 23910 27738 23962
rect 27738 23910 27752 23962
rect 27776 23910 27790 23962
rect 27790 23910 27802 23962
rect 27802 23910 27832 23962
rect 27856 23910 27866 23962
rect 27866 23910 27912 23962
rect 27616 23908 27672 23910
rect 27696 23908 27752 23910
rect 27776 23908 27832 23910
rect 27856 23908 27912 23910
rect 32616 23962 32672 23964
rect 32696 23962 32752 23964
rect 32776 23962 32832 23964
rect 32856 23962 32912 23964
rect 32616 23910 32662 23962
rect 32662 23910 32672 23962
rect 32696 23910 32726 23962
rect 32726 23910 32738 23962
rect 32738 23910 32752 23962
rect 32776 23910 32790 23962
rect 32790 23910 32802 23962
rect 32802 23910 32832 23962
rect 32856 23910 32866 23962
rect 32866 23910 32912 23962
rect 32616 23908 32672 23910
rect 32696 23908 32752 23910
rect 32776 23908 32832 23910
rect 32856 23908 32912 23910
rect 37616 23962 37672 23964
rect 37696 23962 37752 23964
rect 37776 23962 37832 23964
rect 37856 23962 37912 23964
rect 37616 23910 37662 23962
rect 37662 23910 37672 23962
rect 37696 23910 37726 23962
rect 37726 23910 37738 23962
rect 37738 23910 37752 23962
rect 37776 23910 37790 23962
rect 37790 23910 37802 23962
rect 37802 23910 37832 23962
rect 37856 23910 37866 23962
rect 37866 23910 37912 23962
rect 37616 23908 37672 23910
rect 37696 23908 37752 23910
rect 37776 23908 37832 23910
rect 37856 23908 37912 23910
rect 42616 23962 42672 23964
rect 42696 23962 42752 23964
rect 42776 23962 42832 23964
rect 42856 23962 42912 23964
rect 42616 23910 42662 23962
rect 42662 23910 42672 23962
rect 42696 23910 42726 23962
rect 42726 23910 42738 23962
rect 42738 23910 42752 23962
rect 42776 23910 42790 23962
rect 42790 23910 42802 23962
rect 42802 23910 42832 23962
rect 42856 23910 42866 23962
rect 42866 23910 42912 23962
rect 42616 23908 42672 23910
rect 42696 23908 42752 23910
rect 42776 23908 42832 23910
rect 42856 23908 42912 23910
rect 47616 23962 47672 23964
rect 47696 23962 47752 23964
rect 47776 23962 47832 23964
rect 47856 23962 47912 23964
rect 47616 23910 47662 23962
rect 47662 23910 47672 23962
rect 47696 23910 47726 23962
rect 47726 23910 47738 23962
rect 47738 23910 47752 23962
rect 47776 23910 47790 23962
rect 47790 23910 47802 23962
rect 47802 23910 47832 23962
rect 47856 23910 47866 23962
rect 47866 23910 47912 23962
rect 47616 23908 47672 23910
rect 47696 23908 47752 23910
rect 47776 23908 47832 23910
rect 47856 23908 47912 23910
rect 52616 23962 52672 23964
rect 52696 23962 52752 23964
rect 52776 23962 52832 23964
rect 52856 23962 52912 23964
rect 52616 23910 52662 23962
rect 52662 23910 52672 23962
rect 52696 23910 52726 23962
rect 52726 23910 52738 23962
rect 52738 23910 52752 23962
rect 52776 23910 52790 23962
rect 52790 23910 52802 23962
rect 52802 23910 52832 23962
rect 52856 23910 52866 23962
rect 52866 23910 52912 23962
rect 52616 23908 52672 23910
rect 52696 23908 52752 23910
rect 52776 23908 52832 23910
rect 52856 23908 52912 23910
rect 57616 23962 57672 23964
rect 57696 23962 57752 23964
rect 57776 23962 57832 23964
rect 57856 23962 57912 23964
rect 57616 23910 57662 23962
rect 57662 23910 57672 23962
rect 57696 23910 57726 23962
rect 57726 23910 57738 23962
rect 57738 23910 57752 23962
rect 57776 23910 57790 23962
rect 57790 23910 57802 23962
rect 57802 23910 57832 23962
rect 57856 23910 57866 23962
rect 57866 23910 57912 23962
rect 57616 23908 57672 23910
rect 57696 23908 57752 23910
rect 57776 23908 57832 23910
rect 57856 23908 57912 23910
rect 58530 23704 58586 23760
rect 1956 23418 2012 23420
rect 2036 23418 2092 23420
rect 2116 23418 2172 23420
rect 2196 23418 2252 23420
rect 1956 23366 2002 23418
rect 2002 23366 2012 23418
rect 2036 23366 2066 23418
rect 2066 23366 2078 23418
rect 2078 23366 2092 23418
rect 2116 23366 2130 23418
rect 2130 23366 2142 23418
rect 2142 23366 2172 23418
rect 2196 23366 2206 23418
rect 2206 23366 2252 23418
rect 1956 23364 2012 23366
rect 2036 23364 2092 23366
rect 2116 23364 2172 23366
rect 2196 23364 2252 23366
rect 6956 23418 7012 23420
rect 7036 23418 7092 23420
rect 7116 23418 7172 23420
rect 7196 23418 7252 23420
rect 6956 23366 7002 23418
rect 7002 23366 7012 23418
rect 7036 23366 7066 23418
rect 7066 23366 7078 23418
rect 7078 23366 7092 23418
rect 7116 23366 7130 23418
rect 7130 23366 7142 23418
rect 7142 23366 7172 23418
rect 7196 23366 7206 23418
rect 7206 23366 7252 23418
rect 6956 23364 7012 23366
rect 7036 23364 7092 23366
rect 7116 23364 7172 23366
rect 7196 23364 7252 23366
rect 11956 23418 12012 23420
rect 12036 23418 12092 23420
rect 12116 23418 12172 23420
rect 12196 23418 12252 23420
rect 11956 23366 12002 23418
rect 12002 23366 12012 23418
rect 12036 23366 12066 23418
rect 12066 23366 12078 23418
rect 12078 23366 12092 23418
rect 12116 23366 12130 23418
rect 12130 23366 12142 23418
rect 12142 23366 12172 23418
rect 12196 23366 12206 23418
rect 12206 23366 12252 23418
rect 11956 23364 12012 23366
rect 12036 23364 12092 23366
rect 12116 23364 12172 23366
rect 12196 23364 12252 23366
rect 16956 23418 17012 23420
rect 17036 23418 17092 23420
rect 17116 23418 17172 23420
rect 17196 23418 17252 23420
rect 16956 23366 17002 23418
rect 17002 23366 17012 23418
rect 17036 23366 17066 23418
rect 17066 23366 17078 23418
rect 17078 23366 17092 23418
rect 17116 23366 17130 23418
rect 17130 23366 17142 23418
rect 17142 23366 17172 23418
rect 17196 23366 17206 23418
rect 17206 23366 17252 23418
rect 16956 23364 17012 23366
rect 17036 23364 17092 23366
rect 17116 23364 17172 23366
rect 17196 23364 17252 23366
rect 21956 23418 22012 23420
rect 22036 23418 22092 23420
rect 22116 23418 22172 23420
rect 22196 23418 22252 23420
rect 21956 23366 22002 23418
rect 22002 23366 22012 23418
rect 22036 23366 22066 23418
rect 22066 23366 22078 23418
rect 22078 23366 22092 23418
rect 22116 23366 22130 23418
rect 22130 23366 22142 23418
rect 22142 23366 22172 23418
rect 22196 23366 22206 23418
rect 22206 23366 22252 23418
rect 21956 23364 22012 23366
rect 22036 23364 22092 23366
rect 22116 23364 22172 23366
rect 22196 23364 22252 23366
rect 26956 23418 27012 23420
rect 27036 23418 27092 23420
rect 27116 23418 27172 23420
rect 27196 23418 27252 23420
rect 26956 23366 27002 23418
rect 27002 23366 27012 23418
rect 27036 23366 27066 23418
rect 27066 23366 27078 23418
rect 27078 23366 27092 23418
rect 27116 23366 27130 23418
rect 27130 23366 27142 23418
rect 27142 23366 27172 23418
rect 27196 23366 27206 23418
rect 27206 23366 27252 23418
rect 26956 23364 27012 23366
rect 27036 23364 27092 23366
rect 27116 23364 27172 23366
rect 27196 23364 27252 23366
rect 31956 23418 32012 23420
rect 32036 23418 32092 23420
rect 32116 23418 32172 23420
rect 32196 23418 32252 23420
rect 31956 23366 32002 23418
rect 32002 23366 32012 23418
rect 32036 23366 32066 23418
rect 32066 23366 32078 23418
rect 32078 23366 32092 23418
rect 32116 23366 32130 23418
rect 32130 23366 32142 23418
rect 32142 23366 32172 23418
rect 32196 23366 32206 23418
rect 32206 23366 32252 23418
rect 31956 23364 32012 23366
rect 32036 23364 32092 23366
rect 32116 23364 32172 23366
rect 32196 23364 32252 23366
rect 36956 23418 37012 23420
rect 37036 23418 37092 23420
rect 37116 23418 37172 23420
rect 37196 23418 37252 23420
rect 36956 23366 37002 23418
rect 37002 23366 37012 23418
rect 37036 23366 37066 23418
rect 37066 23366 37078 23418
rect 37078 23366 37092 23418
rect 37116 23366 37130 23418
rect 37130 23366 37142 23418
rect 37142 23366 37172 23418
rect 37196 23366 37206 23418
rect 37206 23366 37252 23418
rect 36956 23364 37012 23366
rect 37036 23364 37092 23366
rect 37116 23364 37172 23366
rect 37196 23364 37252 23366
rect 41956 23418 42012 23420
rect 42036 23418 42092 23420
rect 42116 23418 42172 23420
rect 42196 23418 42252 23420
rect 41956 23366 42002 23418
rect 42002 23366 42012 23418
rect 42036 23366 42066 23418
rect 42066 23366 42078 23418
rect 42078 23366 42092 23418
rect 42116 23366 42130 23418
rect 42130 23366 42142 23418
rect 42142 23366 42172 23418
rect 42196 23366 42206 23418
rect 42206 23366 42252 23418
rect 41956 23364 42012 23366
rect 42036 23364 42092 23366
rect 42116 23364 42172 23366
rect 42196 23364 42252 23366
rect 46956 23418 47012 23420
rect 47036 23418 47092 23420
rect 47116 23418 47172 23420
rect 47196 23418 47252 23420
rect 46956 23366 47002 23418
rect 47002 23366 47012 23418
rect 47036 23366 47066 23418
rect 47066 23366 47078 23418
rect 47078 23366 47092 23418
rect 47116 23366 47130 23418
rect 47130 23366 47142 23418
rect 47142 23366 47172 23418
rect 47196 23366 47206 23418
rect 47206 23366 47252 23418
rect 46956 23364 47012 23366
rect 47036 23364 47092 23366
rect 47116 23364 47172 23366
rect 47196 23364 47252 23366
rect 51956 23418 52012 23420
rect 52036 23418 52092 23420
rect 52116 23418 52172 23420
rect 52196 23418 52252 23420
rect 51956 23366 52002 23418
rect 52002 23366 52012 23418
rect 52036 23366 52066 23418
rect 52066 23366 52078 23418
rect 52078 23366 52092 23418
rect 52116 23366 52130 23418
rect 52130 23366 52142 23418
rect 52142 23366 52172 23418
rect 52196 23366 52206 23418
rect 52206 23366 52252 23418
rect 51956 23364 52012 23366
rect 52036 23364 52092 23366
rect 52116 23364 52172 23366
rect 52196 23364 52252 23366
rect 56956 23418 57012 23420
rect 57036 23418 57092 23420
rect 57116 23418 57172 23420
rect 57196 23418 57252 23420
rect 56956 23366 57002 23418
rect 57002 23366 57012 23418
rect 57036 23366 57066 23418
rect 57066 23366 57078 23418
rect 57078 23366 57092 23418
rect 57116 23366 57130 23418
rect 57130 23366 57142 23418
rect 57142 23366 57172 23418
rect 57196 23366 57206 23418
rect 57206 23366 57252 23418
rect 56956 23364 57012 23366
rect 57036 23364 57092 23366
rect 57116 23364 57172 23366
rect 57196 23364 57252 23366
rect 58530 22888 58586 22944
rect 2616 22874 2672 22876
rect 2696 22874 2752 22876
rect 2776 22874 2832 22876
rect 2856 22874 2912 22876
rect 2616 22822 2662 22874
rect 2662 22822 2672 22874
rect 2696 22822 2726 22874
rect 2726 22822 2738 22874
rect 2738 22822 2752 22874
rect 2776 22822 2790 22874
rect 2790 22822 2802 22874
rect 2802 22822 2832 22874
rect 2856 22822 2866 22874
rect 2866 22822 2912 22874
rect 2616 22820 2672 22822
rect 2696 22820 2752 22822
rect 2776 22820 2832 22822
rect 2856 22820 2912 22822
rect 7616 22874 7672 22876
rect 7696 22874 7752 22876
rect 7776 22874 7832 22876
rect 7856 22874 7912 22876
rect 7616 22822 7662 22874
rect 7662 22822 7672 22874
rect 7696 22822 7726 22874
rect 7726 22822 7738 22874
rect 7738 22822 7752 22874
rect 7776 22822 7790 22874
rect 7790 22822 7802 22874
rect 7802 22822 7832 22874
rect 7856 22822 7866 22874
rect 7866 22822 7912 22874
rect 7616 22820 7672 22822
rect 7696 22820 7752 22822
rect 7776 22820 7832 22822
rect 7856 22820 7912 22822
rect 12616 22874 12672 22876
rect 12696 22874 12752 22876
rect 12776 22874 12832 22876
rect 12856 22874 12912 22876
rect 12616 22822 12662 22874
rect 12662 22822 12672 22874
rect 12696 22822 12726 22874
rect 12726 22822 12738 22874
rect 12738 22822 12752 22874
rect 12776 22822 12790 22874
rect 12790 22822 12802 22874
rect 12802 22822 12832 22874
rect 12856 22822 12866 22874
rect 12866 22822 12912 22874
rect 12616 22820 12672 22822
rect 12696 22820 12752 22822
rect 12776 22820 12832 22822
rect 12856 22820 12912 22822
rect 17616 22874 17672 22876
rect 17696 22874 17752 22876
rect 17776 22874 17832 22876
rect 17856 22874 17912 22876
rect 17616 22822 17662 22874
rect 17662 22822 17672 22874
rect 17696 22822 17726 22874
rect 17726 22822 17738 22874
rect 17738 22822 17752 22874
rect 17776 22822 17790 22874
rect 17790 22822 17802 22874
rect 17802 22822 17832 22874
rect 17856 22822 17866 22874
rect 17866 22822 17912 22874
rect 17616 22820 17672 22822
rect 17696 22820 17752 22822
rect 17776 22820 17832 22822
rect 17856 22820 17912 22822
rect 22616 22874 22672 22876
rect 22696 22874 22752 22876
rect 22776 22874 22832 22876
rect 22856 22874 22912 22876
rect 22616 22822 22662 22874
rect 22662 22822 22672 22874
rect 22696 22822 22726 22874
rect 22726 22822 22738 22874
rect 22738 22822 22752 22874
rect 22776 22822 22790 22874
rect 22790 22822 22802 22874
rect 22802 22822 22832 22874
rect 22856 22822 22866 22874
rect 22866 22822 22912 22874
rect 22616 22820 22672 22822
rect 22696 22820 22752 22822
rect 22776 22820 22832 22822
rect 22856 22820 22912 22822
rect 27616 22874 27672 22876
rect 27696 22874 27752 22876
rect 27776 22874 27832 22876
rect 27856 22874 27912 22876
rect 27616 22822 27662 22874
rect 27662 22822 27672 22874
rect 27696 22822 27726 22874
rect 27726 22822 27738 22874
rect 27738 22822 27752 22874
rect 27776 22822 27790 22874
rect 27790 22822 27802 22874
rect 27802 22822 27832 22874
rect 27856 22822 27866 22874
rect 27866 22822 27912 22874
rect 27616 22820 27672 22822
rect 27696 22820 27752 22822
rect 27776 22820 27832 22822
rect 27856 22820 27912 22822
rect 32616 22874 32672 22876
rect 32696 22874 32752 22876
rect 32776 22874 32832 22876
rect 32856 22874 32912 22876
rect 32616 22822 32662 22874
rect 32662 22822 32672 22874
rect 32696 22822 32726 22874
rect 32726 22822 32738 22874
rect 32738 22822 32752 22874
rect 32776 22822 32790 22874
rect 32790 22822 32802 22874
rect 32802 22822 32832 22874
rect 32856 22822 32866 22874
rect 32866 22822 32912 22874
rect 32616 22820 32672 22822
rect 32696 22820 32752 22822
rect 32776 22820 32832 22822
rect 32856 22820 32912 22822
rect 37616 22874 37672 22876
rect 37696 22874 37752 22876
rect 37776 22874 37832 22876
rect 37856 22874 37912 22876
rect 37616 22822 37662 22874
rect 37662 22822 37672 22874
rect 37696 22822 37726 22874
rect 37726 22822 37738 22874
rect 37738 22822 37752 22874
rect 37776 22822 37790 22874
rect 37790 22822 37802 22874
rect 37802 22822 37832 22874
rect 37856 22822 37866 22874
rect 37866 22822 37912 22874
rect 37616 22820 37672 22822
rect 37696 22820 37752 22822
rect 37776 22820 37832 22822
rect 37856 22820 37912 22822
rect 42616 22874 42672 22876
rect 42696 22874 42752 22876
rect 42776 22874 42832 22876
rect 42856 22874 42912 22876
rect 42616 22822 42662 22874
rect 42662 22822 42672 22874
rect 42696 22822 42726 22874
rect 42726 22822 42738 22874
rect 42738 22822 42752 22874
rect 42776 22822 42790 22874
rect 42790 22822 42802 22874
rect 42802 22822 42832 22874
rect 42856 22822 42866 22874
rect 42866 22822 42912 22874
rect 42616 22820 42672 22822
rect 42696 22820 42752 22822
rect 42776 22820 42832 22822
rect 42856 22820 42912 22822
rect 47616 22874 47672 22876
rect 47696 22874 47752 22876
rect 47776 22874 47832 22876
rect 47856 22874 47912 22876
rect 47616 22822 47662 22874
rect 47662 22822 47672 22874
rect 47696 22822 47726 22874
rect 47726 22822 47738 22874
rect 47738 22822 47752 22874
rect 47776 22822 47790 22874
rect 47790 22822 47802 22874
rect 47802 22822 47832 22874
rect 47856 22822 47866 22874
rect 47866 22822 47912 22874
rect 47616 22820 47672 22822
rect 47696 22820 47752 22822
rect 47776 22820 47832 22822
rect 47856 22820 47912 22822
rect 52616 22874 52672 22876
rect 52696 22874 52752 22876
rect 52776 22874 52832 22876
rect 52856 22874 52912 22876
rect 52616 22822 52662 22874
rect 52662 22822 52672 22874
rect 52696 22822 52726 22874
rect 52726 22822 52738 22874
rect 52738 22822 52752 22874
rect 52776 22822 52790 22874
rect 52790 22822 52802 22874
rect 52802 22822 52832 22874
rect 52856 22822 52866 22874
rect 52866 22822 52912 22874
rect 52616 22820 52672 22822
rect 52696 22820 52752 22822
rect 52776 22820 52832 22822
rect 52856 22820 52912 22822
rect 57616 22874 57672 22876
rect 57696 22874 57752 22876
rect 57776 22874 57832 22876
rect 57856 22874 57912 22876
rect 57616 22822 57662 22874
rect 57662 22822 57672 22874
rect 57696 22822 57726 22874
rect 57726 22822 57738 22874
rect 57738 22822 57752 22874
rect 57776 22822 57790 22874
rect 57790 22822 57802 22874
rect 57802 22822 57832 22874
rect 57856 22822 57866 22874
rect 57866 22822 57912 22874
rect 57616 22820 57672 22822
rect 57696 22820 57752 22822
rect 57776 22820 57832 22822
rect 57856 22820 57912 22822
rect 1956 22330 2012 22332
rect 2036 22330 2092 22332
rect 2116 22330 2172 22332
rect 2196 22330 2252 22332
rect 1956 22278 2002 22330
rect 2002 22278 2012 22330
rect 2036 22278 2066 22330
rect 2066 22278 2078 22330
rect 2078 22278 2092 22330
rect 2116 22278 2130 22330
rect 2130 22278 2142 22330
rect 2142 22278 2172 22330
rect 2196 22278 2206 22330
rect 2206 22278 2252 22330
rect 1956 22276 2012 22278
rect 2036 22276 2092 22278
rect 2116 22276 2172 22278
rect 2196 22276 2252 22278
rect 6956 22330 7012 22332
rect 7036 22330 7092 22332
rect 7116 22330 7172 22332
rect 7196 22330 7252 22332
rect 6956 22278 7002 22330
rect 7002 22278 7012 22330
rect 7036 22278 7066 22330
rect 7066 22278 7078 22330
rect 7078 22278 7092 22330
rect 7116 22278 7130 22330
rect 7130 22278 7142 22330
rect 7142 22278 7172 22330
rect 7196 22278 7206 22330
rect 7206 22278 7252 22330
rect 6956 22276 7012 22278
rect 7036 22276 7092 22278
rect 7116 22276 7172 22278
rect 7196 22276 7252 22278
rect 11956 22330 12012 22332
rect 12036 22330 12092 22332
rect 12116 22330 12172 22332
rect 12196 22330 12252 22332
rect 11956 22278 12002 22330
rect 12002 22278 12012 22330
rect 12036 22278 12066 22330
rect 12066 22278 12078 22330
rect 12078 22278 12092 22330
rect 12116 22278 12130 22330
rect 12130 22278 12142 22330
rect 12142 22278 12172 22330
rect 12196 22278 12206 22330
rect 12206 22278 12252 22330
rect 11956 22276 12012 22278
rect 12036 22276 12092 22278
rect 12116 22276 12172 22278
rect 12196 22276 12252 22278
rect 16956 22330 17012 22332
rect 17036 22330 17092 22332
rect 17116 22330 17172 22332
rect 17196 22330 17252 22332
rect 16956 22278 17002 22330
rect 17002 22278 17012 22330
rect 17036 22278 17066 22330
rect 17066 22278 17078 22330
rect 17078 22278 17092 22330
rect 17116 22278 17130 22330
rect 17130 22278 17142 22330
rect 17142 22278 17172 22330
rect 17196 22278 17206 22330
rect 17206 22278 17252 22330
rect 16956 22276 17012 22278
rect 17036 22276 17092 22278
rect 17116 22276 17172 22278
rect 17196 22276 17252 22278
rect 21956 22330 22012 22332
rect 22036 22330 22092 22332
rect 22116 22330 22172 22332
rect 22196 22330 22252 22332
rect 21956 22278 22002 22330
rect 22002 22278 22012 22330
rect 22036 22278 22066 22330
rect 22066 22278 22078 22330
rect 22078 22278 22092 22330
rect 22116 22278 22130 22330
rect 22130 22278 22142 22330
rect 22142 22278 22172 22330
rect 22196 22278 22206 22330
rect 22206 22278 22252 22330
rect 21956 22276 22012 22278
rect 22036 22276 22092 22278
rect 22116 22276 22172 22278
rect 22196 22276 22252 22278
rect 26956 22330 27012 22332
rect 27036 22330 27092 22332
rect 27116 22330 27172 22332
rect 27196 22330 27252 22332
rect 26956 22278 27002 22330
rect 27002 22278 27012 22330
rect 27036 22278 27066 22330
rect 27066 22278 27078 22330
rect 27078 22278 27092 22330
rect 27116 22278 27130 22330
rect 27130 22278 27142 22330
rect 27142 22278 27172 22330
rect 27196 22278 27206 22330
rect 27206 22278 27252 22330
rect 26956 22276 27012 22278
rect 27036 22276 27092 22278
rect 27116 22276 27172 22278
rect 27196 22276 27252 22278
rect 31956 22330 32012 22332
rect 32036 22330 32092 22332
rect 32116 22330 32172 22332
rect 32196 22330 32252 22332
rect 31956 22278 32002 22330
rect 32002 22278 32012 22330
rect 32036 22278 32066 22330
rect 32066 22278 32078 22330
rect 32078 22278 32092 22330
rect 32116 22278 32130 22330
rect 32130 22278 32142 22330
rect 32142 22278 32172 22330
rect 32196 22278 32206 22330
rect 32206 22278 32252 22330
rect 31956 22276 32012 22278
rect 32036 22276 32092 22278
rect 32116 22276 32172 22278
rect 32196 22276 32252 22278
rect 36956 22330 37012 22332
rect 37036 22330 37092 22332
rect 37116 22330 37172 22332
rect 37196 22330 37252 22332
rect 36956 22278 37002 22330
rect 37002 22278 37012 22330
rect 37036 22278 37066 22330
rect 37066 22278 37078 22330
rect 37078 22278 37092 22330
rect 37116 22278 37130 22330
rect 37130 22278 37142 22330
rect 37142 22278 37172 22330
rect 37196 22278 37206 22330
rect 37206 22278 37252 22330
rect 36956 22276 37012 22278
rect 37036 22276 37092 22278
rect 37116 22276 37172 22278
rect 37196 22276 37252 22278
rect 41956 22330 42012 22332
rect 42036 22330 42092 22332
rect 42116 22330 42172 22332
rect 42196 22330 42252 22332
rect 41956 22278 42002 22330
rect 42002 22278 42012 22330
rect 42036 22278 42066 22330
rect 42066 22278 42078 22330
rect 42078 22278 42092 22330
rect 42116 22278 42130 22330
rect 42130 22278 42142 22330
rect 42142 22278 42172 22330
rect 42196 22278 42206 22330
rect 42206 22278 42252 22330
rect 41956 22276 42012 22278
rect 42036 22276 42092 22278
rect 42116 22276 42172 22278
rect 42196 22276 42252 22278
rect 46956 22330 47012 22332
rect 47036 22330 47092 22332
rect 47116 22330 47172 22332
rect 47196 22330 47252 22332
rect 46956 22278 47002 22330
rect 47002 22278 47012 22330
rect 47036 22278 47066 22330
rect 47066 22278 47078 22330
rect 47078 22278 47092 22330
rect 47116 22278 47130 22330
rect 47130 22278 47142 22330
rect 47142 22278 47172 22330
rect 47196 22278 47206 22330
rect 47206 22278 47252 22330
rect 46956 22276 47012 22278
rect 47036 22276 47092 22278
rect 47116 22276 47172 22278
rect 47196 22276 47252 22278
rect 51956 22330 52012 22332
rect 52036 22330 52092 22332
rect 52116 22330 52172 22332
rect 52196 22330 52252 22332
rect 51956 22278 52002 22330
rect 52002 22278 52012 22330
rect 52036 22278 52066 22330
rect 52066 22278 52078 22330
rect 52078 22278 52092 22330
rect 52116 22278 52130 22330
rect 52130 22278 52142 22330
rect 52142 22278 52172 22330
rect 52196 22278 52206 22330
rect 52206 22278 52252 22330
rect 51956 22276 52012 22278
rect 52036 22276 52092 22278
rect 52116 22276 52172 22278
rect 52196 22276 52252 22278
rect 56956 22330 57012 22332
rect 57036 22330 57092 22332
rect 57116 22330 57172 22332
rect 57196 22330 57252 22332
rect 56956 22278 57002 22330
rect 57002 22278 57012 22330
rect 57036 22278 57066 22330
rect 57066 22278 57078 22330
rect 57078 22278 57092 22330
rect 57116 22278 57130 22330
rect 57130 22278 57142 22330
rect 57142 22278 57172 22330
rect 57196 22278 57206 22330
rect 57206 22278 57252 22330
rect 56956 22276 57012 22278
rect 57036 22276 57092 22278
rect 57116 22276 57172 22278
rect 57196 22276 57252 22278
rect 58530 22072 58586 22128
rect 2616 21786 2672 21788
rect 2696 21786 2752 21788
rect 2776 21786 2832 21788
rect 2856 21786 2912 21788
rect 2616 21734 2662 21786
rect 2662 21734 2672 21786
rect 2696 21734 2726 21786
rect 2726 21734 2738 21786
rect 2738 21734 2752 21786
rect 2776 21734 2790 21786
rect 2790 21734 2802 21786
rect 2802 21734 2832 21786
rect 2856 21734 2866 21786
rect 2866 21734 2912 21786
rect 2616 21732 2672 21734
rect 2696 21732 2752 21734
rect 2776 21732 2832 21734
rect 2856 21732 2912 21734
rect 7616 21786 7672 21788
rect 7696 21786 7752 21788
rect 7776 21786 7832 21788
rect 7856 21786 7912 21788
rect 7616 21734 7662 21786
rect 7662 21734 7672 21786
rect 7696 21734 7726 21786
rect 7726 21734 7738 21786
rect 7738 21734 7752 21786
rect 7776 21734 7790 21786
rect 7790 21734 7802 21786
rect 7802 21734 7832 21786
rect 7856 21734 7866 21786
rect 7866 21734 7912 21786
rect 7616 21732 7672 21734
rect 7696 21732 7752 21734
rect 7776 21732 7832 21734
rect 7856 21732 7912 21734
rect 12616 21786 12672 21788
rect 12696 21786 12752 21788
rect 12776 21786 12832 21788
rect 12856 21786 12912 21788
rect 12616 21734 12662 21786
rect 12662 21734 12672 21786
rect 12696 21734 12726 21786
rect 12726 21734 12738 21786
rect 12738 21734 12752 21786
rect 12776 21734 12790 21786
rect 12790 21734 12802 21786
rect 12802 21734 12832 21786
rect 12856 21734 12866 21786
rect 12866 21734 12912 21786
rect 12616 21732 12672 21734
rect 12696 21732 12752 21734
rect 12776 21732 12832 21734
rect 12856 21732 12912 21734
rect 17616 21786 17672 21788
rect 17696 21786 17752 21788
rect 17776 21786 17832 21788
rect 17856 21786 17912 21788
rect 17616 21734 17662 21786
rect 17662 21734 17672 21786
rect 17696 21734 17726 21786
rect 17726 21734 17738 21786
rect 17738 21734 17752 21786
rect 17776 21734 17790 21786
rect 17790 21734 17802 21786
rect 17802 21734 17832 21786
rect 17856 21734 17866 21786
rect 17866 21734 17912 21786
rect 17616 21732 17672 21734
rect 17696 21732 17752 21734
rect 17776 21732 17832 21734
rect 17856 21732 17912 21734
rect 22616 21786 22672 21788
rect 22696 21786 22752 21788
rect 22776 21786 22832 21788
rect 22856 21786 22912 21788
rect 22616 21734 22662 21786
rect 22662 21734 22672 21786
rect 22696 21734 22726 21786
rect 22726 21734 22738 21786
rect 22738 21734 22752 21786
rect 22776 21734 22790 21786
rect 22790 21734 22802 21786
rect 22802 21734 22832 21786
rect 22856 21734 22866 21786
rect 22866 21734 22912 21786
rect 22616 21732 22672 21734
rect 22696 21732 22752 21734
rect 22776 21732 22832 21734
rect 22856 21732 22912 21734
rect 27616 21786 27672 21788
rect 27696 21786 27752 21788
rect 27776 21786 27832 21788
rect 27856 21786 27912 21788
rect 27616 21734 27662 21786
rect 27662 21734 27672 21786
rect 27696 21734 27726 21786
rect 27726 21734 27738 21786
rect 27738 21734 27752 21786
rect 27776 21734 27790 21786
rect 27790 21734 27802 21786
rect 27802 21734 27832 21786
rect 27856 21734 27866 21786
rect 27866 21734 27912 21786
rect 27616 21732 27672 21734
rect 27696 21732 27752 21734
rect 27776 21732 27832 21734
rect 27856 21732 27912 21734
rect 32616 21786 32672 21788
rect 32696 21786 32752 21788
rect 32776 21786 32832 21788
rect 32856 21786 32912 21788
rect 32616 21734 32662 21786
rect 32662 21734 32672 21786
rect 32696 21734 32726 21786
rect 32726 21734 32738 21786
rect 32738 21734 32752 21786
rect 32776 21734 32790 21786
rect 32790 21734 32802 21786
rect 32802 21734 32832 21786
rect 32856 21734 32866 21786
rect 32866 21734 32912 21786
rect 32616 21732 32672 21734
rect 32696 21732 32752 21734
rect 32776 21732 32832 21734
rect 32856 21732 32912 21734
rect 37616 21786 37672 21788
rect 37696 21786 37752 21788
rect 37776 21786 37832 21788
rect 37856 21786 37912 21788
rect 37616 21734 37662 21786
rect 37662 21734 37672 21786
rect 37696 21734 37726 21786
rect 37726 21734 37738 21786
rect 37738 21734 37752 21786
rect 37776 21734 37790 21786
rect 37790 21734 37802 21786
rect 37802 21734 37832 21786
rect 37856 21734 37866 21786
rect 37866 21734 37912 21786
rect 37616 21732 37672 21734
rect 37696 21732 37752 21734
rect 37776 21732 37832 21734
rect 37856 21732 37912 21734
rect 42616 21786 42672 21788
rect 42696 21786 42752 21788
rect 42776 21786 42832 21788
rect 42856 21786 42912 21788
rect 42616 21734 42662 21786
rect 42662 21734 42672 21786
rect 42696 21734 42726 21786
rect 42726 21734 42738 21786
rect 42738 21734 42752 21786
rect 42776 21734 42790 21786
rect 42790 21734 42802 21786
rect 42802 21734 42832 21786
rect 42856 21734 42866 21786
rect 42866 21734 42912 21786
rect 42616 21732 42672 21734
rect 42696 21732 42752 21734
rect 42776 21732 42832 21734
rect 42856 21732 42912 21734
rect 47616 21786 47672 21788
rect 47696 21786 47752 21788
rect 47776 21786 47832 21788
rect 47856 21786 47912 21788
rect 47616 21734 47662 21786
rect 47662 21734 47672 21786
rect 47696 21734 47726 21786
rect 47726 21734 47738 21786
rect 47738 21734 47752 21786
rect 47776 21734 47790 21786
rect 47790 21734 47802 21786
rect 47802 21734 47832 21786
rect 47856 21734 47866 21786
rect 47866 21734 47912 21786
rect 47616 21732 47672 21734
rect 47696 21732 47752 21734
rect 47776 21732 47832 21734
rect 47856 21732 47912 21734
rect 52616 21786 52672 21788
rect 52696 21786 52752 21788
rect 52776 21786 52832 21788
rect 52856 21786 52912 21788
rect 52616 21734 52662 21786
rect 52662 21734 52672 21786
rect 52696 21734 52726 21786
rect 52726 21734 52738 21786
rect 52738 21734 52752 21786
rect 52776 21734 52790 21786
rect 52790 21734 52802 21786
rect 52802 21734 52832 21786
rect 52856 21734 52866 21786
rect 52866 21734 52912 21786
rect 52616 21732 52672 21734
rect 52696 21732 52752 21734
rect 52776 21732 52832 21734
rect 52856 21732 52912 21734
rect 57616 21786 57672 21788
rect 57696 21786 57752 21788
rect 57776 21786 57832 21788
rect 57856 21786 57912 21788
rect 57616 21734 57662 21786
rect 57662 21734 57672 21786
rect 57696 21734 57726 21786
rect 57726 21734 57738 21786
rect 57738 21734 57752 21786
rect 57776 21734 57790 21786
rect 57790 21734 57802 21786
rect 57802 21734 57832 21786
rect 57856 21734 57866 21786
rect 57866 21734 57912 21786
rect 57616 21732 57672 21734
rect 57696 21732 57752 21734
rect 57776 21732 57832 21734
rect 57856 21732 57912 21734
rect 58530 21292 58532 21312
rect 58532 21292 58584 21312
rect 58584 21292 58586 21312
rect 58530 21256 58586 21292
rect 1956 21242 2012 21244
rect 2036 21242 2092 21244
rect 2116 21242 2172 21244
rect 2196 21242 2252 21244
rect 1956 21190 2002 21242
rect 2002 21190 2012 21242
rect 2036 21190 2066 21242
rect 2066 21190 2078 21242
rect 2078 21190 2092 21242
rect 2116 21190 2130 21242
rect 2130 21190 2142 21242
rect 2142 21190 2172 21242
rect 2196 21190 2206 21242
rect 2206 21190 2252 21242
rect 1956 21188 2012 21190
rect 2036 21188 2092 21190
rect 2116 21188 2172 21190
rect 2196 21188 2252 21190
rect 6956 21242 7012 21244
rect 7036 21242 7092 21244
rect 7116 21242 7172 21244
rect 7196 21242 7252 21244
rect 6956 21190 7002 21242
rect 7002 21190 7012 21242
rect 7036 21190 7066 21242
rect 7066 21190 7078 21242
rect 7078 21190 7092 21242
rect 7116 21190 7130 21242
rect 7130 21190 7142 21242
rect 7142 21190 7172 21242
rect 7196 21190 7206 21242
rect 7206 21190 7252 21242
rect 6956 21188 7012 21190
rect 7036 21188 7092 21190
rect 7116 21188 7172 21190
rect 7196 21188 7252 21190
rect 11956 21242 12012 21244
rect 12036 21242 12092 21244
rect 12116 21242 12172 21244
rect 12196 21242 12252 21244
rect 11956 21190 12002 21242
rect 12002 21190 12012 21242
rect 12036 21190 12066 21242
rect 12066 21190 12078 21242
rect 12078 21190 12092 21242
rect 12116 21190 12130 21242
rect 12130 21190 12142 21242
rect 12142 21190 12172 21242
rect 12196 21190 12206 21242
rect 12206 21190 12252 21242
rect 11956 21188 12012 21190
rect 12036 21188 12092 21190
rect 12116 21188 12172 21190
rect 12196 21188 12252 21190
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 17002 21242
rect 17002 21190 17012 21242
rect 17036 21190 17066 21242
rect 17066 21190 17078 21242
rect 17078 21190 17092 21242
rect 17116 21190 17130 21242
rect 17130 21190 17142 21242
rect 17142 21190 17172 21242
rect 17196 21190 17206 21242
rect 17206 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 21956 21242 22012 21244
rect 22036 21242 22092 21244
rect 22116 21242 22172 21244
rect 22196 21242 22252 21244
rect 21956 21190 22002 21242
rect 22002 21190 22012 21242
rect 22036 21190 22066 21242
rect 22066 21190 22078 21242
rect 22078 21190 22092 21242
rect 22116 21190 22130 21242
rect 22130 21190 22142 21242
rect 22142 21190 22172 21242
rect 22196 21190 22206 21242
rect 22206 21190 22252 21242
rect 21956 21188 22012 21190
rect 22036 21188 22092 21190
rect 22116 21188 22172 21190
rect 22196 21188 22252 21190
rect 26956 21242 27012 21244
rect 27036 21242 27092 21244
rect 27116 21242 27172 21244
rect 27196 21242 27252 21244
rect 26956 21190 27002 21242
rect 27002 21190 27012 21242
rect 27036 21190 27066 21242
rect 27066 21190 27078 21242
rect 27078 21190 27092 21242
rect 27116 21190 27130 21242
rect 27130 21190 27142 21242
rect 27142 21190 27172 21242
rect 27196 21190 27206 21242
rect 27206 21190 27252 21242
rect 26956 21188 27012 21190
rect 27036 21188 27092 21190
rect 27116 21188 27172 21190
rect 27196 21188 27252 21190
rect 31956 21242 32012 21244
rect 32036 21242 32092 21244
rect 32116 21242 32172 21244
rect 32196 21242 32252 21244
rect 31956 21190 32002 21242
rect 32002 21190 32012 21242
rect 32036 21190 32066 21242
rect 32066 21190 32078 21242
rect 32078 21190 32092 21242
rect 32116 21190 32130 21242
rect 32130 21190 32142 21242
rect 32142 21190 32172 21242
rect 32196 21190 32206 21242
rect 32206 21190 32252 21242
rect 31956 21188 32012 21190
rect 32036 21188 32092 21190
rect 32116 21188 32172 21190
rect 32196 21188 32252 21190
rect 36956 21242 37012 21244
rect 37036 21242 37092 21244
rect 37116 21242 37172 21244
rect 37196 21242 37252 21244
rect 36956 21190 37002 21242
rect 37002 21190 37012 21242
rect 37036 21190 37066 21242
rect 37066 21190 37078 21242
rect 37078 21190 37092 21242
rect 37116 21190 37130 21242
rect 37130 21190 37142 21242
rect 37142 21190 37172 21242
rect 37196 21190 37206 21242
rect 37206 21190 37252 21242
rect 36956 21188 37012 21190
rect 37036 21188 37092 21190
rect 37116 21188 37172 21190
rect 37196 21188 37252 21190
rect 41956 21242 42012 21244
rect 42036 21242 42092 21244
rect 42116 21242 42172 21244
rect 42196 21242 42252 21244
rect 41956 21190 42002 21242
rect 42002 21190 42012 21242
rect 42036 21190 42066 21242
rect 42066 21190 42078 21242
rect 42078 21190 42092 21242
rect 42116 21190 42130 21242
rect 42130 21190 42142 21242
rect 42142 21190 42172 21242
rect 42196 21190 42206 21242
rect 42206 21190 42252 21242
rect 41956 21188 42012 21190
rect 42036 21188 42092 21190
rect 42116 21188 42172 21190
rect 42196 21188 42252 21190
rect 46956 21242 47012 21244
rect 47036 21242 47092 21244
rect 47116 21242 47172 21244
rect 47196 21242 47252 21244
rect 46956 21190 47002 21242
rect 47002 21190 47012 21242
rect 47036 21190 47066 21242
rect 47066 21190 47078 21242
rect 47078 21190 47092 21242
rect 47116 21190 47130 21242
rect 47130 21190 47142 21242
rect 47142 21190 47172 21242
rect 47196 21190 47206 21242
rect 47206 21190 47252 21242
rect 46956 21188 47012 21190
rect 47036 21188 47092 21190
rect 47116 21188 47172 21190
rect 47196 21188 47252 21190
rect 51956 21242 52012 21244
rect 52036 21242 52092 21244
rect 52116 21242 52172 21244
rect 52196 21242 52252 21244
rect 51956 21190 52002 21242
rect 52002 21190 52012 21242
rect 52036 21190 52066 21242
rect 52066 21190 52078 21242
rect 52078 21190 52092 21242
rect 52116 21190 52130 21242
rect 52130 21190 52142 21242
rect 52142 21190 52172 21242
rect 52196 21190 52206 21242
rect 52206 21190 52252 21242
rect 51956 21188 52012 21190
rect 52036 21188 52092 21190
rect 52116 21188 52172 21190
rect 52196 21188 52252 21190
rect 56956 21242 57012 21244
rect 57036 21242 57092 21244
rect 57116 21242 57172 21244
rect 57196 21242 57252 21244
rect 56956 21190 57002 21242
rect 57002 21190 57012 21242
rect 57036 21190 57066 21242
rect 57066 21190 57078 21242
rect 57078 21190 57092 21242
rect 57116 21190 57130 21242
rect 57130 21190 57142 21242
rect 57142 21190 57172 21242
rect 57196 21190 57206 21242
rect 57206 21190 57252 21242
rect 56956 21188 57012 21190
rect 57036 21188 57092 21190
rect 57116 21188 57172 21190
rect 57196 21188 57252 21190
rect 2616 20698 2672 20700
rect 2696 20698 2752 20700
rect 2776 20698 2832 20700
rect 2856 20698 2912 20700
rect 2616 20646 2662 20698
rect 2662 20646 2672 20698
rect 2696 20646 2726 20698
rect 2726 20646 2738 20698
rect 2738 20646 2752 20698
rect 2776 20646 2790 20698
rect 2790 20646 2802 20698
rect 2802 20646 2832 20698
rect 2856 20646 2866 20698
rect 2866 20646 2912 20698
rect 2616 20644 2672 20646
rect 2696 20644 2752 20646
rect 2776 20644 2832 20646
rect 2856 20644 2912 20646
rect 7616 20698 7672 20700
rect 7696 20698 7752 20700
rect 7776 20698 7832 20700
rect 7856 20698 7912 20700
rect 7616 20646 7662 20698
rect 7662 20646 7672 20698
rect 7696 20646 7726 20698
rect 7726 20646 7738 20698
rect 7738 20646 7752 20698
rect 7776 20646 7790 20698
rect 7790 20646 7802 20698
rect 7802 20646 7832 20698
rect 7856 20646 7866 20698
rect 7866 20646 7912 20698
rect 7616 20644 7672 20646
rect 7696 20644 7752 20646
rect 7776 20644 7832 20646
rect 7856 20644 7912 20646
rect 12616 20698 12672 20700
rect 12696 20698 12752 20700
rect 12776 20698 12832 20700
rect 12856 20698 12912 20700
rect 12616 20646 12662 20698
rect 12662 20646 12672 20698
rect 12696 20646 12726 20698
rect 12726 20646 12738 20698
rect 12738 20646 12752 20698
rect 12776 20646 12790 20698
rect 12790 20646 12802 20698
rect 12802 20646 12832 20698
rect 12856 20646 12866 20698
rect 12866 20646 12912 20698
rect 12616 20644 12672 20646
rect 12696 20644 12752 20646
rect 12776 20644 12832 20646
rect 12856 20644 12912 20646
rect 17616 20698 17672 20700
rect 17696 20698 17752 20700
rect 17776 20698 17832 20700
rect 17856 20698 17912 20700
rect 17616 20646 17662 20698
rect 17662 20646 17672 20698
rect 17696 20646 17726 20698
rect 17726 20646 17738 20698
rect 17738 20646 17752 20698
rect 17776 20646 17790 20698
rect 17790 20646 17802 20698
rect 17802 20646 17832 20698
rect 17856 20646 17866 20698
rect 17866 20646 17912 20698
rect 17616 20644 17672 20646
rect 17696 20644 17752 20646
rect 17776 20644 17832 20646
rect 17856 20644 17912 20646
rect 22616 20698 22672 20700
rect 22696 20698 22752 20700
rect 22776 20698 22832 20700
rect 22856 20698 22912 20700
rect 22616 20646 22662 20698
rect 22662 20646 22672 20698
rect 22696 20646 22726 20698
rect 22726 20646 22738 20698
rect 22738 20646 22752 20698
rect 22776 20646 22790 20698
rect 22790 20646 22802 20698
rect 22802 20646 22832 20698
rect 22856 20646 22866 20698
rect 22866 20646 22912 20698
rect 22616 20644 22672 20646
rect 22696 20644 22752 20646
rect 22776 20644 22832 20646
rect 22856 20644 22912 20646
rect 27616 20698 27672 20700
rect 27696 20698 27752 20700
rect 27776 20698 27832 20700
rect 27856 20698 27912 20700
rect 27616 20646 27662 20698
rect 27662 20646 27672 20698
rect 27696 20646 27726 20698
rect 27726 20646 27738 20698
rect 27738 20646 27752 20698
rect 27776 20646 27790 20698
rect 27790 20646 27802 20698
rect 27802 20646 27832 20698
rect 27856 20646 27866 20698
rect 27866 20646 27912 20698
rect 27616 20644 27672 20646
rect 27696 20644 27752 20646
rect 27776 20644 27832 20646
rect 27856 20644 27912 20646
rect 32616 20698 32672 20700
rect 32696 20698 32752 20700
rect 32776 20698 32832 20700
rect 32856 20698 32912 20700
rect 32616 20646 32662 20698
rect 32662 20646 32672 20698
rect 32696 20646 32726 20698
rect 32726 20646 32738 20698
rect 32738 20646 32752 20698
rect 32776 20646 32790 20698
rect 32790 20646 32802 20698
rect 32802 20646 32832 20698
rect 32856 20646 32866 20698
rect 32866 20646 32912 20698
rect 32616 20644 32672 20646
rect 32696 20644 32752 20646
rect 32776 20644 32832 20646
rect 32856 20644 32912 20646
rect 37616 20698 37672 20700
rect 37696 20698 37752 20700
rect 37776 20698 37832 20700
rect 37856 20698 37912 20700
rect 37616 20646 37662 20698
rect 37662 20646 37672 20698
rect 37696 20646 37726 20698
rect 37726 20646 37738 20698
rect 37738 20646 37752 20698
rect 37776 20646 37790 20698
rect 37790 20646 37802 20698
rect 37802 20646 37832 20698
rect 37856 20646 37866 20698
rect 37866 20646 37912 20698
rect 37616 20644 37672 20646
rect 37696 20644 37752 20646
rect 37776 20644 37832 20646
rect 37856 20644 37912 20646
rect 42616 20698 42672 20700
rect 42696 20698 42752 20700
rect 42776 20698 42832 20700
rect 42856 20698 42912 20700
rect 42616 20646 42662 20698
rect 42662 20646 42672 20698
rect 42696 20646 42726 20698
rect 42726 20646 42738 20698
rect 42738 20646 42752 20698
rect 42776 20646 42790 20698
rect 42790 20646 42802 20698
rect 42802 20646 42832 20698
rect 42856 20646 42866 20698
rect 42866 20646 42912 20698
rect 42616 20644 42672 20646
rect 42696 20644 42752 20646
rect 42776 20644 42832 20646
rect 42856 20644 42912 20646
rect 47616 20698 47672 20700
rect 47696 20698 47752 20700
rect 47776 20698 47832 20700
rect 47856 20698 47912 20700
rect 47616 20646 47662 20698
rect 47662 20646 47672 20698
rect 47696 20646 47726 20698
rect 47726 20646 47738 20698
rect 47738 20646 47752 20698
rect 47776 20646 47790 20698
rect 47790 20646 47802 20698
rect 47802 20646 47832 20698
rect 47856 20646 47866 20698
rect 47866 20646 47912 20698
rect 47616 20644 47672 20646
rect 47696 20644 47752 20646
rect 47776 20644 47832 20646
rect 47856 20644 47912 20646
rect 52616 20698 52672 20700
rect 52696 20698 52752 20700
rect 52776 20698 52832 20700
rect 52856 20698 52912 20700
rect 52616 20646 52662 20698
rect 52662 20646 52672 20698
rect 52696 20646 52726 20698
rect 52726 20646 52738 20698
rect 52738 20646 52752 20698
rect 52776 20646 52790 20698
rect 52790 20646 52802 20698
rect 52802 20646 52832 20698
rect 52856 20646 52866 20698
rect 52866 20646 52912 20698
rect 52616 20644 52672 20646
rect 52696 20644 52752 20646
rect 52776 20644 52832 20646
rect 52856 20644 52912 20646
rect 57616 20698 57672 20700
rect 57696 20698 57752 20700
rect 57776 20698 57832 20700
rect 57856 20698 57912 20700
rect 57616 20646 57662 20698
rect 57662 20646 57672 20698
rect 57696 20646 57726 20698
rect 57726 20646 57738 20698
rect 57738 20646 57752 20698
rect 57776 20646 57790 20698
rect 57790 20646 57802 20698
rect 57802 20646 57832 20698
rect 57856 20646 57866 20698
rect 57866 20646 57912 20698
rect 57616 20644 57672 20646
rect 57696 20644 57752 20646
rect 57776 20644 57832 20646
rect 57856 20644 57912 20646
rect 58530 20440 58586 20496
rect 1956 20154 2012 20156
rect 2036 20154 2092 20156
rect 2116 20154 2172 20156
rect 2196 20154 2252 20156
rect 1956 20102 2002 20154
rect 2002 20102 2012 20154
rect 2036 20102 2066 20154
rect 2066 20102 2078 20154
rect 2078 20102 2092 20154
rect 2116 20102 2130 20154
rect 2130 20102 2142 20154
rect 2142 20102 2172 20154
rect 2196 20102 2206 20154
rect 2206 20102 2252 20154
rect 1956 20100 2012 20102
rect 2036 20100 2092 20102
rect 2116 20100 2172 20102
rect 2196 20100 2252 20102
rect 6956 20154 7012 20156
rect 7036 20154 7092 20156
rect 7116 20154 7172 20156
rect 7196 20154 7252 20156
rect 6956 20102 7002 20154
rect 7002 20102 7012 20154
rect 7036 20102 7066 20154
rect 7066 20102 7078 20154
rect 7078 20102 7092 20154
rect 7116 20102 7130 20154
rect 7130 20102 7142 20154
rect 7142 20102 7172 20154
rect 7196 20102 7206 20154
rect 7206 20102 7252 20154
rect 6956 20100 7012 20102
rect 7036 20100 7092 20102
rect 7116 20100 7172 20102
rect 7196 20100 7252 20102
rect 11956 20154 12012 20156
rect 12036 20154 12092 20156
rect 12116 20154 12172 20156
rect 12196 20154 12252 20156
rect 11956 20102 12002 20154
rect 12002 20102 12012 20154
rect 12036 20102 12066 20154
rect 12066 20102 12078 20154
rect 12078 20102 12092 20154
rect 12116 20102 12130 20154
rect 12130 20102 12142 20154
rect 12142 20102 12172 20154
rect 12196 20102 12206 20154
rect 12206 20102 12252 20154
rect 11956 20100 12012 20102
rect 12036 20100 12092 20102
rect 12116 20100 12172 20102
rect 12196 20100 12252 20102
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 17002 20154
rect 17002 20102 17012 20154
rect 17036 20102 17066 20154
rect 17066 20102 17078 20154
rect 17078 20102 17092 20154
rect 17116 20102 17130 20154
rect 17130 20102 17142 20154
rect 17142 20102 17172 20154
rect 17196 20102 17206 20154
rect 17206 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 21956 20154 22012 20156
rect 22036 20154 22092 20156
rect 22116 20154 22172 20156
rect 22196 20154 22252 20156
rect 21956 20102 22002 20154
rect 22002 20102 22012 20154
rect 22036 20102 22066 20154
rect 22066 20102 22078 20154
rect 22078 20102 22092 20154
rect 22116 20102 22130 20154
rect 22130 20102 22142 20154
rect 22142 20102 22172 20154
rect 22196 20102 22206 20154
rect 22206 20102 22252 20154
rect 21956 20100 22012 20102
rect 22036 20100 22092 20102
rect 22116 20100 22172 20102
rect 22196 20100 22252 20102
rect 26956 20154 27012 20156
rect 27036 20154 27092 20156
rect 27116 20154 27172 20156
rect 27196 20154 27252 20156
rect 26956 20102 27002 20154
rect 27002 20102 27012 20154
rect 27036 20102 27066 20154
rect 27066 20102 27078 20154
rect 27078 20102 27092 20154
rect 27116 20102 27130 20154
rect 27130 20102 27142 20154
rect 27142 20102 27172 20154
rect 27196 20102 27206 20154
rect 27206 20102 27252 20154
rect 26956 20100 27012 20102
rect 27036 20100 27092 20102
rect 27116 20100 27172 20102
rect 27196 20100 27252 20102
rect 31956 20154 32012 20156
rect 32036 20154 32092 20156
rect 32116 20154 32172 20156
rect 32196 20154 32252 20156
rect 31956 20102 32002 20154
rect 32002 20102 32012 20154
rect 32036 20102 32066 20154
rect 32066 20102 32078 20154
rect 32078 20102 32092 20154
rect 32116 20102 32130 20154
rect 32130 20102 32142 20154
rect 32142 20102 32172 20154
rect 32196 20102 32206 20154
rect 32206 20102 32252 20154
rect 31956 20100 32012 20102
rect 32036 20100 32092 20102
rect 32116 20100 32172 20102
rect 32196 20100 32252 20102
rect 36956 20154 37012 20156
rect 37036 20154 37092 20156
rect 37116 20154 37172 20156
rect 37196 20154 37252 20156
rect 36956 20102 37002 20154
rect 37002 20102 37012 20154
rect 37036 20102 37066 20154
rect 37066 20102 37078 20154
rect 37078 20102 37092 20154
rect 37116 20102 37130 20154
rect 37130 20102 37142 20154
rect 37142 20102 37172 20154
rect 37196 20102 37206 20154
rect 37206 20102 37252 20154
rect 36956 20100 37012 20102
rect 37036 20100 37092 20102
rect 37116 20100 37172 20102
rect 37196 20100 37252 20102
rect 41956 20154 42012 20156
rect 42036 20154 42092 20156
rect 42116 20154 42172 20156
rect 42196 20154 42252 20156
rect 41956 20102 42002 20154
rect 42002 20102 42012 20154
rect 42036 20102 42066 20154
rect 42066 20102 42078 20154
rect 42078 20102 42092 20154
rect 42116 20102 42130 20154
rect 42130 20102 42142 20154
rect 42142 20102 42172 20154
rect 42196 20102 42206 20154
rect 42206 20102 42252 20154
rect 41956 20100 42012 20102
rect 42036 20100 42092 20102
rect 42116 20100 42172 20102
rect 42196 20100 42252 20102
rect 46956 20154 47012 20156
rect 47036 20154 47092 20156
rect 47116 20154 47172 20156
rect 47196 20154 47252 20156
rect 46956 20102 47002 20154
rect 47002 20102 47012 20154
rect 47036 20102 47066 20154
rect 47066 20102 47078 20154
rect 47078 20102 47092 20154
rect 47116 20102 47130 20154
rect 47130 20102 47142 20154
rect 47142 20102 47172 20154
rect 47196 20102 47206 20154
rect 47206 20102 47252 20154
rect 46956 20100 47012 20102
rect 47036 20100 47092 20102
rect 47116 20100 47172 20102
rect 47196 20100 47252 20102
rect 51956 20154 52012 20156
rect 52036 20154 52092 20156
rect 52116 20154 52172 20156
rect 52196 20154 52252 20156
rect 51956 20102 52002 20154
rect 52002 20102 52012 20154
rect 52036 20102 52066 20154
rect 52066 20102 52078 20154
rect 52078 20102 52092 20154
rect 52116 20102 52130 20154
rect 52130 20102 52142 20154
rect 52142 20102 52172 20154
rect 52196 20102 52206 20154
rect 52206 20102 52252 20154
rect 51956 20100 52012 20102
rect 52036 20100 52092 20102
rect 52116 20100 52172 20102
rect 52196 20100 52252 20102
rect 56956 20154 57012 20156
rect 57036 20154 57092 20156
rect 57116 20154 57172 20156
rect 57196 20154 57252 20156
rect 56956 20102 57002 20154
rect 57002 20102 57012 20154
rect 57036 20102 57066 20154
rect 57066 20102 57078 20154
rect 57078 20102 57092 20154
rect 57116 20102 57130 20154
rect 57130 20102 57142 20154
rect 57142 20102 57172 20154
rect 57196 20102 57206 20154
rect 57206 20102 57252 20154
rect 56956 20100 57012 20102
rect 57036 20100 57092 20102
rect 57116 20100 57172 20102
rect 57196 20100 57252 20102
rect 58530 19624 58586 19680
rect 2616 19610 2672 19612
rect 2696 19610 2752 19612
rect 2776 19610 2832 19612
rect 2856 19610 2912 19612
rect 2616 19558 2662 19610
rect 2662 19558 2672 19610
rect 2696 19558 2726 19610
rect 2726 19558 2738 19610
rect 2738 19558 2752 19610
rect 2776 19558 2790 19610
rect 2790 19558 2802 19610
rect 2802 19558 2832 19610
rect 2856 19558 2866 19610
rect 2866 19558 2912 19610
rect 2616 19556 2672 19558
rect 2696 19556 2752 19558
rect 2776 19556 2832 19558
rect 2856 19556 2912 19558
rect 7616 19610 7672 19612
rect 7696 19610 7752 19612
rect 7776 19610 7832 19612
rect 7856 19610 7912 19612
rect 7616 19558 7662 19610
rect 7662 19558 7672 19610
rect 7696 19558 7726 19610
rect 7726 19558 7738 19610
rect 7738 19558 7752 19610
rect 7776 19558 7790 19610
rect 7790 19558 7802 19610
rect 7802 19558 7832 19610
rect 7856 19558 7866 19610
rect 7866 19558 7912 19610
rect 7616 19556 7672 19558
rect 7696 19556 7752 19558
rect 7776 19556 7832 19558
rect 7856 19556 7912 19558
rect 12616 19610 12672 19612
rect 12696 19610 12752 19612
rect 12776 19610 12832 19612
rect 12856 19610 12912 19612
rect 12616 19558 12662 19610
rect 12662 19558 12672 19610
rect 12696 19558 12726 19610
rect 12726 19558 12738 19610
rect 12738 19558 12752 19610
rect 12776 19558 12790 19610
rect 12790 19558 12802 19610
rect 12802 19558 12832 19610
rect 12856 19558 12866 19610
rect 12866 19558 12912 19610
rect 12616 19556 12672 19558
rect 12696 19556 12752 19558
rect 12776 19556 12832 19558
rect 12856 19556 12912 19558
rect 17616 19610 17672 19612
rect 17696 19610 17752 19612
rect 17776 19610 17832 19612
rect 17856 19610 17912 19612
rect 17616 19558 17662 19610
rect 17662 19558 17672 19610
rect 17696 19558 17726 19610
rect 17726 19558 17738 19610
rect 17738 19558 17752 19610
rect 17776 19558 17790 19610
rect 17790 19558 17802 19610
rect 17802 19558 17832 19610
rect 17856 19558 17866 19610
rect 17866 19558 17912 19610
rect 17616 19556 17672 19558
rect 17696 19556 17752 19558
rect 17776 19556 17832 19558
rect 17856 19556 17912 19558
rect 22616 19610 22672 19612
rect 22696 19610 22752 19612
rect 22776 19610 22832 19612
rect 22856 19610 22912 19612
rect 22616 19558 22662 19610
rect 22662 19558 22672 19610
rect 22696 19558 22726 19610
rect 22726 19558 22738 19610
rect 22738 19558 22752 19610
rect 22776 19558 22790 19610
rect 22790 19558 22802 19610
rect 22802 19558 22832 19610
rect 22856 19558 22866 19610
rect 22866 19558 22912 19610
rect 22616 19556 22672 19558
rect 22696 19556 22752 19558
rect 22776 19556 22832 19558
rect 22856 19556 22912 19558
rect 27616 19610 27672 19612
rect 27696 19610 27752 19612
rect 27776 19610 27832 19612
rect 27856 19610 27912 19612
rect 27616 19558 27662 19610
rect 27662 19558 27672 19610
rect 27696 19558 27726 19610
rect 27726 19558 27738 19610
rect 27738 19558 27752 19610
rect 27776 19558 27790 19610
rect 27790 19558 27802 19610
rect 27802 19558 27832 19610
rect 27856 19558 27866 19610
rect 27866 19558 27912 19610
rect 27616 19556 27672 19558
rect 27696 19556 27752 19558
rect 27776 19556 27832 19558
rect 27856 19556 27912 19558
rect 32616 19610 32672 19612
rect 32696 19610 32752 19612
rect 32776 19610 32832 19612
rect 32856 19610 32912 19612
rect 32616 19558 32662 19610
rect 32662 19558 32672 19610
rect 32696 19558 32726 19610
rect 32726 19558 32738 19610
rect 32738 19558 32752 19610
rect 32776 19558 32790 19610
rect 32790 19558 32802 19610
rect 32802 19558 32832 19610
rect 32856 19558 32866 19610
rect 32866 19558 32912 19610
rect 32616 19556 32672 19558
rect 32696 19556 32752 19558
rect 32776 19556 32832 19558
rect 32856 19556 32912 19558
rect 37616 19610 37672 19612
rect 37696 19610 37752 19612
rect 37776 19610 37832 19612
rect 37856 19610 37912 19612
rect 37616 19558 37662 19610
rect 37662 19558 37672 19610
rect 37696 19558 37726 19610
rect 37726 19558 37738 19610
rect 37738 19558 37752 19610
rect 37776 19558 37790 19610
rect 37790 19558 37802 19610
rect 37802 19558 37832 19610
rect 37856 19558 37866 19610
rect 37866 19558 37912 19610
rect 37616 19556 37672 19558
rect 37696 19556 37752 19558
rect 37776 19556 37832 19558
rect 37856 19556 37912 19558
rect 42616 19610 42672 19612
rect 42696 19610 42752 19612
rect 42776 19610 42832 19612
rect 42856 19610 42912 19612
rect 42616 19558 42662 19610
rect 42662 19558 42672 19610
rect 42696 19558 42726 19610
rect 42726 19558 42738 19610
rect 42738 19558 42752 19610
rect 42776 19558 42790 19610
rect 42790 19558 42802 19610
rect 42802 19558 42832 19610
rect 42856 19558 42866 19610
rect 42866 19558 42912 19610
rect 42616 19556 42672 19558
rect 42696 19556 42752 19558
rect 42776 19556 42832 19558
rect 42856 19556 42912 19558
rect 47616 19610 47672 19612
rect 47696 19610 47752 19612
rect 47776 19610 47832 19612
rect 47856 19610 47912 19612
rect 47616 19558 47662 19610
rect 47662 19558 47672 19610
rect 47696 19558 47726 19610
rect 47726 19558 47738 19610
rect 47738 19558 47752 19610
rect 47776 19558 47790 19610
rect 47790 19558 47802 19610
rect 47802 19558 47832 19610
rect 47856 19558 47866 19610
rect 47866 19558 47912 19610
rect 47616 19556 47672 19558
rect 47696 19556 47752 19558
rect 47776 19556 47832 19558
rect 47856 19556 47912 19558
rect 52616 19610 52672 19612
rect 52696 19610 52752 19612
rect 52776 19610 52832 19612
rect 52856 19610 52912 19612
rect 52616 19558 52662 19610
rect 52662 19558 52672 19610
rect 52696 19558 52726 19610
rect 52726 19558 52738 19610
rect 52738 19558 52752 19610
rect 52776 19558 52790 19610
rect 52790 19558 52802 19610
rect 52802 19558 52832 19610
rect 52856 19558 52866 19610
rect 52866 19558 52912 19610
rect 52616 19556 52672 19558
rect 52696 19556 52752 19558
rect 52776 19556 52832 19558
rect 52856 19556 52912 19558
rect 57616 19610 57672 19612
rect 57696 19610 57752 19612
rect 57776 19610 57832 19612
rect 57856 19610 57912 19612
rect 57616 19558 57662 19610
rect 57662 19558 57672 19610
rect 57696 19558 57726 19610
rect 57726 19558 57738 19610
rect 57738 19558 57752 19610
rect 57776 19558 57790 19610
rect 57790 19558 57802 19610
rect 57802 19558 57832 19610
rect 57856 19558 57866 19610
rect 57866 19558 57912 19610
rect 57616 19556 57672 19558
rect 57696 19556 57752 19558
rect 57776 19556 57832 19558
rect 57856 19556 57912 19558
rect 1956 19066 2012 19068
rect 2036 19066 2092 19068
rect 2116 19066 2172 19068
rect 2196 19066 2252 19068
rect 1956 19014 2002 19066
rect 2002 19014 2012 19066
rect 2036 19014 2066 19066
rect 2066 19014 2078 19066
rect 2078 19014 2092 19066
rect 2116 19014 2130 19066
rect 2130 19014 2142 19066
rect 2142 19014 2172 19066
rect 2196 19014 2206 19066
rect 2206 19014 2252 19066
rect 1956 19012 2012 19014
rect 2036 19012 2092 19014
rect 2116 19012 2172 19014
rect 2196 19012 2252 19014
rect 6956 19066 7012 19068
rect 7036 19066 7092 19068
rect 7116 19066 7172 19068
rect 7196 19066 7252 19068
rect 6956 19014 7002 19066
rect 7002 19014 7012 19066
rect 7036 19014 7066 19066
rect 7066 19014 7078 19066
rect 7078 19014 7092 19066
rect 7116 19014 7130 19066
rect 7130 19014 7142 19066
rect 7142 19014 7172 19066
rect 7196 19014 7206 19066
rect 7206 19014 7252 19066
rect 6956 19012 7012 19014
rect 7036 19012 7092 19014
rect 7116 19012 7172 19014
rect 7196 19012 7252 19014
rect 11956 19066 12012 19068
rect 12036 19066 12092 19068
rect 12116 19066 12172 19068
rect 12196 19066 12252 19068
rect 11956 19014 12002 19066
rect 12002 19014 12012 19066
rect 12036 19014 12066 19066
rect 12066 19014 12078 19066
rect 12078 19014 12092 19066
rect 12116 19014 12130 19066
rect 12130 19014 12142 19066
rect 12142 19014 12172 19066
rect 12196 19014 12206 19066
rect 12206 19014 12252 19066
rect 11956 19012 12012 19014
rect 12036 19012 12092 19014
rect 12116 19012 12172 19014
rect 12196 19012 12252 19014
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 17002 19066
rect 17002 19014 17012 19066
rect 17036 19014 17066 19066
rect 17066 19014 17078 19066
rect 17078 19014 17092 19066
rect 17116 19014 17130 19066
rect 17130 19014 17142 19066
rect 17142 19014 17172 19066
rect 17196 19014 17206 19066
rect 17206 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 21956 19066 22012 19068
rect 22036 19066 22092 19068
rect 22116 19066 22172 19068
rect 22196 19066 22252 19068
rect 21956 19014 22002 19066
rect 22002 19014 22012 19066
rect 22036 19014 22066 19066
rect 22066 19014 22078 19066
rect 22078 19014 22092 19066
rect 22116 19014 22130 19066
rect 22130 19014 22142 19066
rect 22142 19014 22172 19066
rect 22196 19014 22206 19066
rect 22206 19014 22252 19066
rect 21956 19012 22012 19014
rect 22036 19012 22092 19014
rect 22116 19012 22172 19014
rect 22196 19012 22252 19014
rect 26956 19066 27012 19068
rect 27036 19066 27092 19068
rect 27116 19066 27172 19068
rect 27196 19066 27252 19068
rect 26956 19014 27002 19066
rect 27002 19014 27012 19066
rect 27036 19014 27066 19066
rect 27066 19014 27078 19066
rect 27078 19014 27092 19066
rect 27116 19014 27130 19066
rect 27130 19014 27142 19066
rect 27142 19014 27172 19066
rect 27196 19014 27206 19066
rect 27206 19014 27252 19066
rect 26956 19012 27012 19014
rect 27036 19012 27092 19014
rect 27116 19012 27172 19014
rect 27196 19012 27252 19014
rect 31956 19066 32012 19068
rect 32036 19066 32092 19068
rect 32116 19066 32172 19068
rect 32196 19066 32252 19068
rect 31956 19014 32002 19066
rect 32002 19014 32012 19066
rect 32036 19014 32066 19066
rect 32066 19014 32078 19066
rect 32078 19014 32092 19066
rect 32116 19014 32130 19066
rect 32130 19014 32142 19066
rect 32142 19014 32172 19066
rect 32196 19014 32206 19066
rect 32206 19014 32252 19066
rect 31956 19012 32012 19014
rect 32036 19012 32092 19014
rect 32116 19012 32172 19014
rect 32196 19012 32252 19014
rect 36956 19066 37012 19068
rect 37036 19066 37092 19068
rect 37116 19066 37172 19068
rect 37196 19066 37252 19068
rect 36956 19014 37002 19066
rect 37002 19014 37012 19066
rect 37036 19014 37066 19066
rect 37066 19014 37078 19066
rect 37078 19014 37092 19066
rect 37116 19014 37130 19066
rect 37130 19014 37142 19066
rect 37142 19014 37172 19066
rect 37196 19014 37206 19066
rect 37206 19014 37252 19066
rect 36956 19012 37012 19014
rect 37036 19012 37092 19014
rect 37116 19012 37172 19014
rect 37196 19012 37252 19014
rect 41956 19066 42012 19068
rect 42036 19066 42092 19068
rect 42116 19066 42172 19068
rect 42196 19066 42252 19068
rect 41956 19014 42002 19066
rect 42002 19014 42012 19066
rect 42036 19014 42066 19066
rect 42066 19014 42078 19066
rect 42078 19014 42092 19066
rect 42116 19014 42130 19066
rect 42130 19014 42142 19066
rect 42142 19014 42172 19066
rect 42196 19014 42206 19066
rect 42206 19014 42252 19066
rect 41956 19012 42012 19014
rect 42036 19012 42092 19014
rect 42116 19012 42172 19014
rect 42196 19012 42252 19014
rect 46956 19066 47012 19068
rect 47036 19066 47092 19068
rect 47116 19066 47172 19068
rect 47196 19066 47252 19068
rect 46956 19014 47002 19066
rect 47002 19014 47012 19066
rect 47036 19014 47066 19066
rect 47066 19014 47078 19066
rect 47078 19014 47092 19066
rect 47116 19014 47130 19066
rect 47130 19014 47142 19066
rect 47142 19014 47172 19066
rect 47196 19014 47206 19066
rect 47206 19014 47252 19066
rect 46956 19012 47012 19014
rect 47036 19012 47092 19014
rect 47116 19012 47172 19014
rect 47196 19012 47252 19014
rect 51956 19066 52012 19068
rect 52036 19066 52092 19068
rect 52116 19066 52172 19068
rect 52196 19066 52252 19068
rect 51956 19014 52002 19066
rect 52002 19014 52012 19066
rect 52036 19014 52066 19066
rect 52066 19014 52078 19066
rect 52078 19014 52092 19066
rect 52116 19014 52130 19066
rect 52130 19014 52142 19066
rect 52142 19014 52172 19066
rect 52196 19014 52206 19066
rect 52206 19014 52252 19066
rect 51956 19012 52012 19014
rect 52036 19012 52092 19014
rect 52116 19012 52172 19014
rect 52196 19012 52252 19014
rect 56956 19066 57012 19068
rect 57036 19066 57092 19068
rect 57116 19066 57172 19068
rect 57196 19066 57252 19068
rect 56956 19014 57002 19066
rect 57002 19014 57012 19066
rect 57036 19014 57066 19066
rect 57066 19014 57078 19066
rect 57078 19014 57092 19066
rect 57116 19014 57130 19066
rect 57130 19014 57142 19066
rect 57142 19014 57172 19066
rect 57196 19014 57206 19066
rect 57206 19014 57252 19066
rect 56956 19012 57012 19014
rect 57036 19012 57092 19014
rect 57116 19012 57172 19014
rect 57196 19012 57252 19014
rect 58530 18808 58586 18864
rect 2616 18522 2672 18524
rect 2696 18522 2752 18524
rect 2776 18522 2832 18524
rect 2856 18522 2912 18524
rect 2616 18470 2662 18522
rect 2662 18470 2672 18522
rect 2696 18470 2726 18522
rect 2726 18470 2738 18522
rect 2738 18470 2752 18522
rect 2776 18470 2790 18522
rect 2790 18470 2802 18522
rect 2802 18470 2832 18522
rect 2856 18470 2866 18522
rect 2866 18470 2912 18522
rect 2616 18468 2672 18470
rect 2696 18468 2752 18470
rect 2776 18468 2832 18470
rect 2856 18468 2912 18470
rect 7616 18522 7672 18524
rect 7696 18522 7752 18524
rect 7776 18522 7832 18524
rect 7856 18522 7912 18524
rect 7616 18470 7662 18522
rect 7662 18470 7672 18522
rect 7696 18470 7726 18522
rect 7726 18470 7738 18522
rect 7738 18470 7752 18522
rect 7776 18470 7790 18522
rect 7790 18470 7802 18522
rect 7802 18470 7832 18522
rect 7856 18470 7866 18522
rect 7866 18470 7912 18522
rect 7616 18468 7672 18470
rect 7696 18468 7752 18470
rect 7776 18468 7832 18470
rect 7856 18468 7912 18470
rect 12616 18522 12672 18524
rect 12696 18522 12752 18524
rect 12776 18522 12832 18524
rect 12856 18522 12912 18524
rect 12616 18470 12662 18522
rect 12662 18470 12672 18522
rect 12696 18470 12726 18522
rect 12726 18470 12738 18522
rect 12738 18470 12752 18522
rect 12776 18470 12790 18522
rect 12790 18470 12802 18522
rect 12802 18470 12832 18522
rect 12856 18470 12866 18522
rect 12866 18470 12912 18522
rect 12616 18468 12672 18470
rect 12696 18468 12752 18470
rect 12776 18468 12832 18470
rect 12856 18468 12912 18470
rect 17616 18522 17672 18524
rect 17696 18522 17752 18524
rect 17776 18522 17832 18524
rect 17856 18522 17912 18524
rect 17616 18470 17662 18522
rect 17662 18470 17672 18522
rect 17696 18470 17726 18522
rect 17726 18470 17738 18522
rect 17738 18470 17752 18522
rect 17776 18470 17790 18522
rect 17790 18470 17802 18522
rect 17802 18470 17832 18522
rect 17856 18470 17866 18522
rect 17866 18470 17912 18522
rect 17616 18468 17672 18470
rect 17696 18468 17752 18470
rect 17776 18468 17832 18470
rect 17856 18468 17912 18470
rect 22616 18522 22672 18524
rect 22696 18522 22752 18524
rect 22776 18522 22832 18524
rect 22856 18522 22912 18524
rect 22616 18470 22662 18522
rect 22662 18470 22672 18522
rect 22696 18470 22726 18522
rect 22726 18470 22738 18522
rect 22738 18470 22752 18522
rect 22776 18470 22790 18522
rect 22790 18470 22802 18522
rect 22802 18470 22832 18522
rect 22856 18470 22866 18522
rect 22866 18470 22912 18522
rect 22616 18468 22672 18470
rect 22696 18468 22752 18470
rect 22776 18468 22832 18470
rect 22856 18468 22912 18470
rect 27616 18522 27672 18524
rect 27696 18522 27752 18524
rect 27776 18522 27832 18524
rect 27856 18522 27912 18524
rect 27616 18470 27662 18522
rect 27662 18470 27672 18522
rect 27696 18470 27726 18522
rect 27726 18470 27738 18522
rect 27738 18470 27752 18522
rect 27776 18470 27790 18522
rect 27790 18470 27802 18522
rect 27802 18470 27832 18522
rect 27856 18470 27866 18522
rect 27866 18470 27912 18522
rect 27616 18468 27672 18470
rect 27696 18468 27752 18470
rect 27776 18468 27832 18470
rect 27856 18468 27912 18470
rect 32616 18522 32672 18524
rect 32696 18522 32752 18524
rect 32776 18522 32832 18524
rect 32856 18522 32912 18524
rect 32616 18470 32662 18522
rect 32662 18470 32672 18522
rect 32696 18470 32726 18522
rect 32726 18470 32738 18522
rect 32738 18470 32752 18522
rect 32776 18470 32790 18522
rect 32790 18470 32802 18522
rect 32802 18470 32832 18522
rect 32856 18470 32866 18522
rect 32866 18470 32912 18522
rect 32616 18468 32672 18470
rect 32696 18468 32752 18470
rect 32776 18468 32832 18470
rect 32856 18468 32912 18470
rect 37616 18522 37672 18524
rect 37696 18522 37752 18524
rect 37776 18522 37832 18524
rect 37856 18522 37912 18524
rect 37616 18470 37662 18522
rect 37662 18470 37672 18522
rect 37696 18470 37726 18522
rect 37726 18470 37738 18522
rect 37738 18470 37752 18522
rect 37776 18470 37790 18522
rect 37790 18470 37802 18522
rect 37802 18470 37832 18522
rect 37856 18470 37866 18522
rect 37866 18470 37912 18522
rect 37616 18468 37672 18470
rect 37696 18468 37752 18470
rect 37776 18468 37832 18470
rect 37856 18468 37912 18470
rect 42616 18522 42672 18524
rect 42696 18522 42752 18524
rect 42776 18522 42832 18524
rect 42856 18522 42912 18524
rect 42616 18470 42662 18522
rect 42662 18470 42672 18522
rect 42696 18470 42726 18522
rect 42726 18470 42738 18522
rect 42738 18470 42752 18522
rect 42776 18470 42790 18522
rect 42790 18470 42802 18522
rect 42802 18470 42832 18522
rect 42856 18470 42866 18522
rect 42866 18470 42912 18522
rect 42616 18468 42672 18470
rect 42696 18468 42752 18470
rect 42776 18468 42832 18470
rect 42856 18468 42912 18470
rect 47616 18522 47672 18524
rect 47696 18522 47752 18524
rect 47776 18522 47832 18524
rect 47856 18522 47912 18524
rect 47616 18470 47662 18522
rect 47662 18470 47672 18522
rect 47696 18470 47726 18522
rect 47726 18470 47738 18522
rect 47738 18470 47752 18522
rect 47776 18470 47790 18522
rect 47790 18470 47802 18522
rect 47802 18470 47832 18522
rect 47856 18470 47866 18522
rect 47866 18470 47912 18522
rect 47616 18468 47672 18470
rect 47696 18468 47752 18470
rect 47776 18468 47832 18470
rect 47856 18468 47912 18470
rect 52616 18522 52672 18524
rect 52696 18522 52752 18524
rect 52776 18522 52832 18524
rect 52856 18522 52912 18524
rect 52616 18470 52662 18522
rect 52662 18470 52672 18522
rect 52696 18470 52726 18522
rect 52726 18470 52738 18522
rect 52738 18470 52752 18522
rect 52776 18470 52790 18522
rect 52790 18470 52802 18522
rect 52802 18470 52832 18522
rect 52856 18470 52866 18522
rect 52866 18470 52912 18522
rect 52616 18468 52672 18470
rect 52696 18468 52752 18470
rect 52776 18468 52832 18470
rect 52856 18468 52912 18470
rect 57616 18522 57672 18524
rect 57696 18522 57752 18524
rect 57776 18522 57832 18524
rect 57856 18522 57912 18524
rect 57616 18470 57662 18522
rect 57662 18470 57672 18522
rect 57696 18470 57726 18522
rect 57726 18470 57738 18522
rect 57738 18470 57752 18522
rect 57776 18470 57790 18522
rect 57790 18470 57802 18522
rect 57802 18470 57832 18522
rect 57856 18470 57866 18522
rect 57866 18470 57912 18522
rect 57616 18468 57672 18470
rect 57696 18468 57752 18470
rect 57776 18468 57832 18470
rect 57856 18468 57912 18470
rect 58530 18028 58532 18048
rect 58532 18028 58584 18048
rect 58584 18028 58586 18048
rect 58530 17992 58586 18028
rect 1956 17978 2012 17980
rect 2036 17978 2092 17980
rect 2116 17978 2172 17980
rect 2196 17978 2252 17980
rect 1956 17926 2002 17978
rect 2002 17926 2012 17978
rect 2036 17926 2066 17978
rect 2066 17926 2078 17978
rect 2078 17926 2092 17978
rect 2116 17926 2130 17978
rect 2130 17926 2142 17978
rect 2142 17926 2172 17978
rect 2196 17926 2206 17978
rect 2206 17926 2252 17978
rect 1956 17924 2012 17926
rect 2036 17924 2092 17926
rect 2116 17924 2172 17926
rect 2196 17924 2252 17926
rect 6956 17978 7012 17980
rect 7036 17978 7092 17980
rect 7116 17978 7172 17980
rect 7196 17978 7252 17980
rect 6956 17926 7002 17978
rect 7002 17926 7012 17978
rect 7036 17926 7066 17978
rect 7066 17926 7078 17978
rect 7078 17926 7092 17978
rect 7116 17926 7130 17978
rect 7130 17926 7142 17978
rect 7142 17926 7172 17978
rect 7196 17926 7206 17978
rect 7206 17926 7252 17978
rect 6956 17924 7012 17926
rect 7036 17924 7092 17926
rect 7116 17924 7172 17926
rect 7196 17924 7252 17926
rect 11956 17978 12012 17980
rect 12036 17978 12092 17980
rect 12116 17978 12172 17980
rect 12196 17978 12252 17980
rect 11956 17926 12002 17978
rect 12002 17926 12012 17978
rect 12036 17926 12066 17978
rect 12066 17926 12078 17978
rect 12078 17926 12092 17978
rect 12116 17926 12130 17978
rect 12130 17926 12142 17978
rect 12142 17926 12172 17978
rect 12196 17926 12206 17978
rect 12206 17926 12252 17978
rect 11956 17924 12012 17926
rect 12036 17924 12092 17926
rect 12116 17924 12172 17926
rect 12196 17924 12252 17926
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 17002 17978
rect 17002 17926 17012 17978
rect 17036 17926 17066 17978
rect 17066 17926 17078 17978
rect 17078 17926 17092 17978
rect 17116 17926 17130 17978
rect 17130 17926 17142 17978
rect 17142 17926 17172 17978
rect 17196 17926 17206 17978
rect 17206 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 21956 17978 22012 17980
rect 22036 17978 22092 17980
rect 22116 17978 22172 17980
rect 22196 17978 22252 17980
rect 21956 17926 22002 17978
rect 22002 17926 22012 17978
rect 22036 17926 22066 17978
rect 22066 17926 22078 17978
rect 22078 17926 22092 17978
rect 22116 17926 22130 17978
rect 22130 17926 22142 17978
rect 22142 17926 22172 17978
rect 22196 17926 22206 17978
rect 22206 17926 22252 17978
rect 21956 17924 22012 17926
rect 22036 17924 22092 17926
rect 22116 17924 22172 17926
rect 22196 17924 22252 17926
rect 26956 17978 27012 17980
rect 27036 17978 27092 17980
rect 27116 17978 27172 17980
rect 27196 17978 27252 17980
rect 26956 17926 27002 17978
rect 27002 17926 27012 17978
rect 27036 17926 27066 17978
rect 27066 17926 27078 17978
rect 27078 17926 27092 17978
rect 27116 17926 27130 17978
rect 27130 17926 27142 17978
rect 27142 17926 27172 17978
rect 27196 17926 27206 17978
rect 27206 17926 27252 17978
rect 26956 17924 27012 17926
rect 27036 17924 27092 17926
rect 27116 17924 27172 17926
rect 27196 17924 27252 17926
rect 31956 17978 32012 17980
rect 32036 17978 32092 17980
rect 32116 17978 32172 17980
rect 32196 17978 32252 17980
rect 31956 17926 32002 17978
rect 32002 17926 32012 17978
rect 32036 17926 32066 17978
rect 32066 17926 32078 17978
rect 32078 17926 32092 17978
rect 32116 17926 32130 17978
rect 32130 17926 32142 17978
rect 32142 17926 32172 17978
rect 32196 17926 32206 17978
rect 32206 17926 32252 17978
rect 31956 17924 32012 17926
rect 32036 17924 32092 17926
rect 32116 17924 32172 17926
rect 32196 17924 32252 17926
rect 36956 17978 37012 17980
rect 37036 17978 37092 17980
rect 37116 17978 37172 17980
rect 37196 17978 37252 17980
rect 36956 17926 37002 17978
rect 37002 17926 37012 17978
rect 37036 17926 37066 17978
rect 37066 17926 37078 17978
rect 37078 17926 37092 17978
rect 37116 17926 37130 17978
rect 37130 17926 37142 17978
rect 37142 17926 37172 17978
rect 37196 17926 37206 17978
rect 37206 17926 37252 17978
rect 36956 17924 37012 17926
rect 37036 17924 37092 17926
rect 37116 17924 37172 17926
rect 37196 17924 37252 17926
rect 41956 17978 42012 17980
rect 42036 17978 42092 17980
rect 42116 17978 42172 17980
rect 42196 17978 42252 17980
rect 41956 17926 42002 17978
rect 42002 17926 42012 17978
rect 42036 17926 42066 17978
rect 42066 17926 42078 17978
rect 42078 17926 42092 17978
rect 42116 17926 42130 17978
rect 42130 17926 42142 17978
rect 42142 17926 42172 17978
rect 42196 17926 42206 17978
rect 42206 17926 42252 17978
rect 41956 17924 42012 17926
rect 42036 17924 42092 17926
rect 42116 17924 42172 17926
rect 42196 17924 42252 17926
rect 46956 17978 47012 17980
rect 47036 17978 47092 17980
rect 47116 17978 47172 17980
rect 47196 17978 47252 17980
rect 46956 17926 47002 17978
rect 47002 17926 47012 17978
rect 47036 17926 47066 17978
rect 47066 17926 47078 17978
rect 47078 17926 47092 17978
rect 47116 17926 47130 17978
rect 47130 17926 47142 17978
rect 47142 17926 47172 17978
rect 47196 17926 47206 17978
rect 47206 17926 47252 17978
rect 46956 17924 47012 17926
rect 47036 17924 47092 17926
rect 47116 17924 47172 17926
rect 47196 17924 47252 17926
rect 51956 17978 52012 17980
rect 52036 17978 52092 17980
rect 52116 17978 52172 17980
rect 52196 17978 52252 17980
rect 51956 17926 52002 17978
rect 52002 17926 52012 17978
rect 52036 17926 52066 17978
rect 52066 17926 52078 17978
rect 52078 17926 52092 17978
rect 52116 17926 52130 17978
rect 52130 17926 52142 17978
rect 52142 17926 52172 17978
rect 52196 17926 52206 17978
rect 52206 17926 52252 17978
rect 51956 17924 52012 17926
rect 52036 17924 52092 17926
rect 52116 17924 52172 17926
rect 52196 17924 52252 17926
rect 56956 17978 57012 17980
rect 57036 17978 57092 17980
rect 57116 17978 57172 17980
rect 57196 17978 57252 17980
rect 56956 17926 57002 17978
rect 57002 17926 57012 17978
rect 57036 17926 57066 17978
rect 57066 17926 57078 17978
rect 57078 17926 57092 17978
rect 57116 17926 57130 17978
rect 57130 17926 57142 17978
rect 57142 17926 57172 17978
rect 57196 17926 57206 17978
rect 57206 17926 57252 17978
rect 56956 17924 57012 17926
rect 57036 17924 57092 17926
rect 57116 17924 57172 17926
rect 57196 17924 57252 17926
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 22616 17434 22672 17436
rect 22696 17434 22752 17436
rect 22776 17434 22832 17436
rect 22856 17434 22912 17436
rect 22616 17382 22662 17434
rect 22662 17382 22672 17434
rect 22696 17382 22726 17434
rect 22726 17382 22738 17434
rect 22738 17382 22752 17434
rect 22776 17382 22790 17434
rect 22790 17382 22802 17434
rect 22802 17382 22832 17434
rect 22856 17382 22866 17434
rect 22866 17382 22912 17434
rect 22616 17380 22672 17382
rect 22696 17380 22752 17382
rect 22776 17380 22832 17382
rect 22856 17380 22912 17382
rect 27616 17434 27672 17436
rect 27696 17434 27752 17436
rect 27776 17434 27832 17436
rect 27856 17434 27912 17436
rect 27616 17382 27662 17434
rect 27662 17382 27672 17434
rect 27696 17382 27726 17434
rect 27726 17382 27738 17434
rect 27738 17382 27752 17434
rect 27776 17382 27790 17434
rect 27790 17382 27802 17434
rect 27802 17382 27832 17434
rect 27856 17382 27866 17434
rect 27866 17382 27912 17434
rect 27616 17380 27672 17382
rect 27696 17380 27752 17382
rect 27776 17380 27832 17382
rect 27856 17380 27912 17382
rect 32616 17434 32672 17436
rect 32696 17434 32752 17436
rect 32776 17434 32832 17436
rect 32856 17434 32912 17436
rect 32616 17382 32662 17434
rect 32662 17382 32672 17434
rect 32696 17382 32726 17434
rect 32726 17382 32738 17434
rect 32738 17382 32752 17434
rect 32776 17382 32790 17434
rect 32790 17382 32802 17434
rect 32802 17382 32832 17434
rect 32856 17382 32866 17434
rect 32866 17382 32912 17434
rect 32616 17380 32672 17382
rect 32696 17380 32752 17382
rect 32776 17380 32832 17382
rect 32856 17380 32912 17382
rect 37616 17434 37672 17436
rect 37696 17434 37752 17436
rect 37776 17434 37832 17436
rect 37856 17434 37912 17436
rect 37616 17382 37662 17434
rect 37662 17382 37672 17434
rect 37696 17382 37726 17434
rect 37726 17382 37738 17434
rect 37738 17382 37752 17434
rect 37776 17382 37790 17434
rect 37790 17382 37802 17434
rect 37802 17382 37832 17434
rect 37856 17382 37866 17434
rect 37866 17382 37912 17434
rect 37616 17380 37672 17382
rect 37696 17380 37752 17382
rect 37776 17380 37832 17382
rect 37856 17380 37912 17382
rect 42616 17434 42672 17436
rect 42696 17434 42752 17436
rect 42776 17434 42832 17436
rect 42856 17434 42912 17436
rect 42616 17382 42662 17434
rect 42662 17382 42672 17434
rect 42696 17382 42726 17434
rect 42726 17382 42738 17434
rect 42738 17382 42752 17434
rect 42776 17382 42790 17434
rect 42790 17382 42802 17434
rect 42802 17382 42832 17434
rect 42856 17382 42866 17434
rect 42866 17382 42912 17434
rect 42616 17380 42672 17382
rect 42696 17380 42752 17382
rect 42776 17380 42832 17382
rect 42856 17380 42912 17382
rect 47616 17434 47672 17436
rect 47696 17434 47752 17436
rect 47776 17434 47832 17436
rect 47856 17434 47912 17436
rect 47616 17382 47662 17434
rect 47662 17382 47672 17434
rect 47696 17382 47726 17434
rect 47726 17382 47738 17434
rect 47738 17382 47752 17434
rect 47776 17382 47790 17434
rect 47790 17382 47802 17434
rect 47802 17382 47832 17434
rect 47856 17382 47866 17434
rect 47866 17382 47912 17434
rect 47616 17380 47672 17382
rect 47696 17380 47752 17382
rect 47776 17380 47832 17382
rect 47856 17380 47912 17382
rect 52616 17434 52672 17436
rect 52696 17434 52752 17436
rect 52776 17434 52832 17436
rect 52856 17434 52912 17436
rect 52616 17382 52662 17434
rect 52662 17382 52672 17434
rect 52696 17382 52726 17434
rect 52726 17382 52738 17434
rect 52738 17382 52752 17434
rect 52776 17382 52790 17434
rect 52790 17382 52802 17434
rect 52802 17382 52832 17434
rect 52856 17382 52866 17434
rect 52866 17382 52912 17434
rect 52616 17380 52672 17382
rect 52696 17380 52752 17382
rect 52776 17380 52832 17382
rect 52856 17380 52912 17382
rect 57616 17434 57672 17436
rect 57696 17434 57752 17436
rect 57776 17434 57832 17436
rect 57856 17434 57912 17436
rect 57616 17382 57662 17434
rect 57662 17382 57672 17434
rect 57696 17382 57726 17434
rect 57726 17382 57738 17434
rect 57738 17382 57752 17434
rect 57776 17382 57790 17434
rect 57790 17382 57802 17434
rect 57802 17382 57832 17434
rect 57856 17382 57866 17434
rect 57866 17382 57912 17434
rect 57616 17380 57672 17382
rect 57696 17380 57752 17382
rect 57776 17380 57832 17382
rect 57856 17380 57912 17382
rect 58530 17176 58586 17232
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 21956 16890 22012 16892
rect 22036 16890 22092 16892
rect 22116 16890 22172 16892
rect 22196 16890 22252 16892
rect 21956 16838 22002 16890
rect 22002 16838 22012 16890
rect 22036 16838 22066 16890
rect 22066 16838 22078 16890
rect 22078 16838 22092 16890
rect 22116 16838 22130 16890
rect 22130 16838 22142 16890
rect 22142 16838 22172 16890
rect 22196 16838 22206 16890
rect 22206 16838 22252 16890
rect 21956 16836 22012 16838
rect 22036 16836 22092 16838
rect 22116 16836 22172 16838
rect 22196 16836 22252 16838
rect 26956 16890 27012 16892
rect 27036 16890 27092 16892
rect 27116 16890 27172 16892
rect 27196 16890 27252 16892
rect 26956 16838 27002 16890
rect 27002 16838 27012 16890
rect 27036 16838 27066 16890
rect 27066 16838 27078 16890
rect 27078 16838 27092 16890
rect 27116 16838 27130 16890
rect 27130 16838 27142 16890
rect 27142 16838 27172 16890
rect 27196 16838 27206 16890
rect 27206 16838 27252 16890
rect 26956 16836 27012 16838
rect 27036 16836 27092 16838
rect 27116 16836 27172 16838
rect 27196 16836 27252 16838
rect 31956 16890 32012 16892
rect 32036 16890 32092 16892
rect 32116 16890 32172 16892
rect 32196 16890 32252 16892
rect 31956 16838 32002 16890
rect 32002 16838 32012 16890
rect 32036 16838 32066 16890
rect 32066 16838 32078 16890
rect 32078 16838 32092 16890
rect 32116 16838 32130 16890
rect 32130 16838 32142 16890
rect 32142 16838 32172 16890
rect 32196 16838 32206 16890
rect 32206 16838 32252 16890
rect 31956 16836 32012 16838
rect 32036 16836 32092 16838
rect 32116 16836 32172 16838
rect 32196 16836 32252 16838
rect 36956 16890 37012 16892
rect 37036 16890 37092 16892
rect 37116 16890 37172 16892
rect 37196 16890 37252 16892
rect 36956 16838 37002 16890
rect 37002 16838 37012 16890
rect 37036 16838 37066 16890
rect 37066 16838 37078 16890
rect 37078 16838 37092 16890
rect 37116 16838 37130 16890
rect 37130 16838 37142 16890
rect 37142 16838 37172 16890
rect 37196 16838 37206 16890
rect 37206 16838 37252 16890
rect 36956 16836 37012 16838
rect 37036 16836 37092 16838
rect 37116 16836 37172 16838
rect 37196 16836 37252 16838
rect 41956 16890 42012 16892
rect 42036 16890 42092 16892
rect 42116 16890 42172 16892
rect 42196 16890 42252 16892
rect 41956 16838 42002 16890
rect 42002 16838 42012 16890
rect 42036 16838 42066 16890
rect 42066 16838 42078 16890
rect 42078 16838 42092 16890
rect 42116 16838 42130 16890
rect 42130 16838 42142 16890
rect 42142 16838 42172 16890
rect 42196 16838 42206 16890
rect 42206 16838 42252 16890
rect 41956 16836 42012 16838
rect 42036 16836 42092 16838
rect 42116 16836 42172 16838
rect 42196 16836 42252 16838
rect 46956 16890 47012 16892
rect 47036 16890 47092 16892
rect 47116 16890 47172 16892
rect 47196 16890 47252 16892
rect 46956 16838 47002 16890
rect 47002 16838 47012 16890
rect 47036 16838 47066 16890
rect 47066 16838 47078 16890
rect 47078 16838 47092 16890
rect 47116 16838 47130 16890
rect 47130 16838 47142 16890
rect 47142 16838 47172 16890
rect 47196 16838 47206 16890
rect 47206 16838 47252 16890
rect 46956 16836 47012 16838
rect 47036 16836 47092 16838
rect 47116 16836 47172 16838
rect 47196 16836 47252 16838
rect 51956 16890 52012 16892
rect 52036 16890 52092 16892
rect 52116 16890 52172 16892
rect 52196 16890 52252 16892
rect 51956 16838 52002 16890
rect 52002 16838 52012 16890
rect 52036 16838 52066 16890
rect 52066 16838 52078 16890
rect 52078 16838 52092 16890
rect 52116 16838 52130 16890
rect 52130 16838 52142 16890
rect 52142 16838 52172 16890
rect 52196 16838 52206 16890
rect 52206 16838 52252 16890
rect 51956 16836 52012 16838
rect 52036 16836 52092 16838
rect 52116 16836 52172 16838
rect 52196 16836 52252 16838
rect 56956 16890 57012 16892
rect 57036 16890 57092 16892
rect 57116 16890 57172 16892
rect 57196 16890 57252 16892
rect 56956 16838 57002 16890
rect 57002 16838 57012 16890
rect 57036 16838 57066 16890
rect 57066 16838 57078 16890
rect 57078 16838 57092 16890
rect 57116 16838 57130 16890
rect 57130 16838 57142 16890
rect 57142 16838 57172 16890
rect 57196 16838 57206 16890
rect 57206 16838 57252 16890
rect 56956 16836 57012 16838
rect 57036 16836 57092 16838
rect 57116 16836 57172 16838
rect 57196 16836 57252 16838
rect 57886 16496 57942 16552
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 22616 16346 22672 16348
rect 22696 16346 22752 16348
rect 22776 16346 22832 16348
rect 22856 16346 22912 16348
rect 22616 16294 22662 16346
rect 22662 16294 22672 16346
rect 22696 16294 22726 16346
rect 22726 16294 22738 16346
rect 22738 16294 22752 16346
rect 22776 16294 22790 16346
rect 22790 16294 22802 16346
rect 22802 16294 22832 16346
rect 22856 16294 22866 16346
rect 22866 16294 22912 16346
rect 22616 16292 22672 16294
rect 22696 16292 22752 16294
rect 22776 16292 22832 16294
rect 22856 16292 22912 16294
rect 27616 16346 27672 16348
rect 27696 16346 27752 16348
rect 27776 16346 27832 16348
rect 27856 16346 27912 16348
rect 27616 16294 27662 16346
rect 27662 16294 27672 16346
rect 27696 16294 27726 16346
rect 27726 16294 27738 16346
rect 27738 16294 27752 16346
rect 27776 16294 27790 16346
rect 27790 16294 27802 16346
rect 27802 16294 27832 16346
rect 27856 16294 27866 16346
rect 27866 16294 27912 16346
rect 27616 16292 27672 16294
rect 27696 16292 27752 16294
rect 27776 16292 27832 16294
rect 27856 16292 27912 16294
rect 32616 16346 32672 16348
rect 32696 16346 32752 16348
rect 32776 16346 32832 16348
rect 32856 16346 32912 16348
rect 32616 16294 32662 16346
rect 32662 16294 32672 16346
rect 32696 16294 32726 16346
rect 32726 16294 32738 16346
rect 32738 16294 32752 16346
rect 32776 16294 32790 16346
rect 32790 16294 32802 16346
rect 32802 16294 32832 16346
rect 32856 16294 32866 16346
rect 32866 16294 32912 16346
rect 32616 16292 32672 16294
rect 32696 16292 32752 16294
rect 32776 16292 32832 16294
rect 32856 16292 32912 16294
rect 37616 16346 37672 16348
rect 37696 16346 37752 16348
rect 37776 16346 37832 16348
rect 37856 16346 37912 16348
rect 37616 16294 37662 16346
rect 37662 16294 37672 16346
rect 37696 16294 37726 16346
rect 37726 16294 37738 16346
rect 37738 16294 37752 16346
rect 37776 16294 37790 16346
rect 37790 16294 37802 16346
rect 37802 16294 37832 16346
rect 37856 16294 37866 16346
rect 37866 16294 37912 16346
rect 37616 16292 37672 16294
rect 37696 16292 37752 16294
rect 37776 16292 37832 16294
rect 37856 16292 37912 16294
rect 42616 16346 42672 16348
rect 42696 16346 42752 16348
rect 42776 16346 42832 16348
rect 42856 16346 42912 16348
rect 42616 16294 42662 16346
rect 42662 16294 42672 16346
rect 42696 16294 42726 16346
rect 42726 16294 42738 16346
rect 42738 16294 42752 16346
rect 42776 16294 42790 16346
rect 42790 16294 42802 16346
rect 42802 16294 42832 16346
rect 42856 16294 42866 16346
rect 42866 16294 42912 16346
rect 42616 16292 42672 16294
rect 42696 16292 42752 16294
rect 42776 16292 42832 16294
rect 42856 16292 42912 16294
rect 47616 16346 47672 16348
rect 47696 16346 47752 16348
rect 47776 16346 47832 16348
rect 47856 16346 47912 16348
rect 47616 16294 47662 16346
rect 47662 16294 47672 16346
rect 47696 16294 47726 16346
rect 47726 16294 47738 16346
rect 47738 16294 47752 16346
rect 47776 16294 47790 16346
rect 47790 16294 47802 16346
rect 47802 16294 47832 16346
rect 47856 16294 47866 16346
rect 47866 16294 47912 16346
rect 47616 16292 47672 16294
rect 47696 16292 47752 16294
rect 47776 16292 47832 16294
rect 47856 16292 47912 16294
rect 52616 16346 52672 16348
rect 52696 16346 52752 16348
rect 52776 16346 52832 16348
rect 52856 16346 52912 16348
rect 52616 16294 52662 16346
rect 52662 16294 52672 16346
rect 52696 16294 52726 16346
rect 52726 16294 52738 16346
rect 52738 16294 52752 16346
rect 52776 16294 52790 16346
rect 52790 16294 52802 16346
rect 52802 16294 52832 16346
rect 52856 16294 52866 16346
rect 52866 16294 52912 16346
rect 52616 16292 52672 16294
rect 52696 16292 52752 16294
rect 52776 16292 52832 16294
rect 52856 16292 52912 16294
rect 57616 16346 57672 16348
rect 57696 16346 57752 16348
rect 57776 16346 57832 16348
rect 57856 16346 57912 16348
rect 57616 16294 57662 16346
rect 57662 16294 57672 16346
rect 57696 16294 57726 16346
rect 57726 16294 57738 16346
rect 57738 16294 57752 16346
rect 57776 16294 57790 16346
rect 57790 16294 57802 16346
rect 57802 16294 57832 16346
rect 57856 16294 57866 16346
rect 57866 16294 57912 16346
rect 57616 16292 57672 16294
rect 57696 16292 57752 16294
rect 57776 16292 57832 16294
rect 57856 16292 57912 16294
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 21956 15802 22012 15804
rect 22036 15802 22092 15804
rect 22116 15802 22172 15804
rect 22196 15802 22252 15804
rect 21956 15750 22002 15802
rect 22002 15750 22012 15802
rect 22036 15750 22066 15802
rect 22066 15750 22078 15802
rect 22078 15750 22092 15802
rect 22116 15750 22130 15802
rect 22130 15750 22142 15802
rect 22142 15750 22172 15802
rect 22196 15750 22206 15802
rect 22206 15750 22252 15802
rect 21956 15748 22012 15750
rect 22036 15748 22092 15750
rect 22116 15748 22172 15750
rect 22196 15748 22252 15750
rect 26956 15802 27012 15804
rect 27036 15802 27092 15804
rect 27116 15802 27172 15804
rect 27196 15802 27252 15804
rect 26956 15750 27002 15802
rect 27002 15750 27012 15802
rect 27036 15750 27066 15802
rect 27066 15750 27078 15802
rect 27078 15750 27092 15802
rect 27116 15750 27130 15802
rect 27130 15750 27142 15802
rect 27142 15750 27172 15802
rect 27196 15750 27206 15802
rect 27206 15750 27252 15802
rect 26956 15748 27012 15750
rect 27036 15748 27092 15750
rect 27116 15748 27172 15750
rect 27196 15748 27252 15750
rect 31956 15802 32012 15804
rect 32036 15802 32092 15804
rect 32116 15802 32172 15804
rect 32196 15802 32252 15804
rect 31956 15750 32002 15802
rect 32002 15750 32012 15802
rect 32036 15750 32066 15802
rect 32066 15750 32078 15802
rect 32078 15750 32092 15802
rect 32116 15750 32130 15802
rect 32130 15750 32142 15802
rect 32142 15750 32172 15802
rect 32196 15750 32206 15802
rect 32206 15750 32252 15802
rect 31956 15748 32012 15750
rect 32036 15748 32092 15750
rect 32116 15748 32172 15750
rect 32196 15748 32252 15750
rect 36956 15802 37012 15804
rect 37036 15802 37092 15804
rect 37116 15802 37172 15804
rect 37196 15802 37252 15804
rect 36956 15750 37002 15802
rect 37002 15750 37012 15802
rect 37036 15750 37066 15802
rect 37066 15750 37078 15802
rect 37078 15750 37092 15802
rect 37116 15750 37130 15802
rect 37130 15750 37142 15802
rect 37142 15750 37172 15802
rect 37196 15750 37206 15802
rect 37206 15750 37252 15802
rect 36956 15748 37012 15750
rect 37036 15748 37092 15750
rect 37116 15748 37172 15750
rect 37196 15748 37252 15750
rect 41956 15802 42012 15804
rect 42036 15802 42092 15804
rect 42116 15802 42172 15804
rect 42196 15802 42252 15804
rect 41956 15750 42002 15802
rect 42002 15750 42012 15802
rect 42036 15750 42066 15802
rect 42066 15750 42078 15802
rect 42078 15750 42092 15802
rect 42116 15750 42130 15802
rect 42130 15750 42142 15802
rect 42142 15750 42172 15802
rect 42196 15750 42206 15802
rect 42206 15750 42252 15802
rect 41956 15748 42012 15750
rect 42036 15748 42092 15750
rect 42116 15748 42172 15750
rect 42196 15748 42252 15750
rect 46956 15802 47012 15804
rect 47036 15802 47092 15804
rect 47116 15802 47172 15804
rect 47196 15802 47252 15804
rect 46956 15750 47002 15802
rect 47002 15750 47012 15802
rect 47036 15750 47066 15802
rect 47066 15750 47078 15802
rect 47078 15750 47092 15802
rect 47116 15750 47130 15802
rect 47130 15750 47142 15802
rect 47142 15750 47172 15802
rect 47196 15750 47206 15802
rect 47206 15750 47252 15802
rect 46956 15748 47012 15750
rect 47036 15748 47092 15750
rect 47116 15748 47172 15750
rect 47196 15748 47252 15750
rect 51956 15802 52012 15804
rect 52036 15802 52092 15804
rect 52116 15802 52172 15804
rect 52196 15802 52252 15804
rect 51956 15750 52002 15802
rect 52002 15750 52012 15802
rect 52036 15750 52066 15802
rect 52066 15750 52078 15802
rect 52078 15750 52092 15802
rect 52116 15750 52130 15802
rect 52130 15750 52142 15802
rect 52142 15750 52172 15802
rect 52196 15750 52206 15802
rect 52206 15750 52252 15802
rect 51956 15748 52012 15750
rect 52036 15748 52092 15750
rect 52116 15748 52172 15750
rect 52196 15748 52252 15750
rect 56956 15802 57012 15804
rect 57036 15802 57092 15804
rect 57116 15802 57172 15804
rect 57196 15802 57252 15804
rect 56956 15750 57002 15802
rect 57002 15750 57012 15802
rect 57036 15750 57066 15802
rect 57066 15750 57078 15802
rect 57078 15750 57092 15802
rect 57116 15750 57130 15802
rect 57130 15750 57142 15802
rect 57142 15750 57172 15802
rect 57196 15750 57206 15802
rect 57206 15750 57252 15802
rect 56956 15748 57012 15750
rect 57036 15748 57092 15750
rect 57116 15748 57172 15750
rect 57196 15748 57252 15750
rect 58530 15544 58586 15600
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 22616 15258 22672 15260
rect 22696 15258 22752 15260
rect 22776 15258 22832 15260
rect 22856 15258 22912 15260
rect 22616 15206 22662 15258
rect 22662 15206 22672 15258
rect 22696 15206 22726 15258
rect 22726 15206 22738 15258
rect 22738 15206 22752 15258
rect 22776 15206 22790 15258
rect 22790 15206 22802 15258
rect 22802 15206 22832 15258
rect 22856 15206 22866 15258
rect 22866 15206 22912 15258
rect 22616 15204 22672 15206
rect 22696 15204 22752 15206
rect 22776 15204 22832 15206
rect 22856 15204 22912 15206
rect 27616 15258 27672 15260
rect 27696 15258 27752 15260
rect 27776 15258 27832 15260
rect 27856 15258 27912 15260
rect 27616 15206 27662 15258
rect 27662 15206 27672 15258
rect 27696 15206 27726 15258
rect 27726 15206 27738 15258
rect 27738 15206 27752 15258
rect 27776 15206 27790 15258
rect 27790 15206 27802 15258
rect 27802 15206 27832 15258
rect 27856 15206 27866 15258
rect 27866 15206 27912 15258
rect 27616 15204 27672 15206
rect 27696 15204 27752 15206
rect 27776 15204 27832 15206
rect 27856 15204 27912 15206
rect 32616 15258 32672 15260
rect 32696 15258 32752 15260
rect 32776 15258 32832 15260
rect 32856 15258 32912 15260
rect 32616 15206 32662 15258
rect 32662 15206 32672 15258
rect 32696 15206 32726 15258
rect 32726 15206 32738 15258
rect 32738 15206 32752 15258
rect 32776 15206 32790 15258
rect 32790 15206 32802 15258
rect 32802 15206 32832 15258
rect 32856 15206 32866 15258
rect 32866 15206 32912 15258
rect 32616 15204 32672 15206
rect 32696 15204 32752 15206
rect 32776 15204 32832 15206
rect 32856 15204 32912 15206
rect 37616 15258 37672 15260
rect 37696 15258 37752 15260
rect 37776 15258 37832 15260
rect 37856 15258 37912 15260
rect 37616 15206 37662 15258
rect 37662 15206 37672 15258
rect 37696 15206 37726 15258
rect 37726 15206 37738 15258
rect 37738 15206 37752 15258
rect 37776 15206 37790 15258
rect 37790 15206 37802 15258
rect 37802 15206 37832 15258
rect 37856 15206 37866 15258
rect 37866 15206 37912 15258
rect 37616 15204 37672 15206
rect 37696 15204 37752 15206
rect 37776 15204 37832 15206
rect 37856 15204 37912 15206
rect 42616 15258 42672 15260
rect 42696 15258 42752 15260
rect 42776 15258 42832 15260
rect 42856 15258 42912 15260
rect 42616 15206 42662 15258
rect 42662 15206 42672 15258
rect 42696 15206 42726 15258
rect 42726 15206 42738 15258
rect 42738 15206 42752 15258
rect 42776 15206 42790 15258
rect 42790 15206 42802 15258
rect 42802 15206 42832 15258
rect 42856 15206 42866 15258
rect 42866 15206 42912 15258
rect 42616 15204 42672 15206
rect 42696 15204 42752 15206
rect 42776 15204 42832 15206
rect 42856 15204 42912 15206
rect 47616 15258 47672 15260
rect 47696 15258 47752 15260
rect 47776 15258 47832 15260
rect 47856 15258 47912 15260
rect 47616 15206 47662 15258
rect 47662 15206 47672 15258
rect 47696 15206 47726 15258
rect 47726 15206 47738 15258
rect 47738 15206 47752 15258
rect 47776 15206 47790 15258
rect 47790 15206 47802 15258
rect 47802 15206 47832 15258
rect 47856 15206 47866 15258
rect 47866 15206 47912 15258
rect 47616 15204 47672 15206
rect 47696 15204 47752 15206
rect 47776 15204 47832 15206
rect 47856 15204 47912 15206
rect 52616 15258 52672 15260
rect 52696 15258 52752 15260
rect 52776 15258 52832 15260
rect 52856 15258 52912 15260
rect 52616 15206 52662 15258
rect 52662 15206 52672 15258
rect 52696 15206 52726 15258
rect 52726 15206 52738 15258
rect 52738 15206 52752 15258
rect 52776 15206 52790 15258
rect 52790 15206 52802 15258
rect 52802 15206 52832 15258
rect 52856 15206 52866 15258
rect 52866 15206 52912 15258
rect 52616 15204 52672 15206
rect 52696 15204 52752 15206
rect 52776 15204 52832 15206
rect 52856 15204 52912 15206
rect 57616 15258 57672 15260
rect 57696 15258 57752 15260
rect 57776 15258 57832 15260
rect 57856 15258 57912 15260
rect 57616 15206 57662 15258
rect 57662 15206 57672 15258
rect 57696 15206 57726 15258
rect 57726 15206 57738 15258
rect 57738 15206 57752 15258
rect 57776 15206 57790 15258
rect 57790 15206 57802 15258
rect 57802 15206 57832 15258
rect 57856 15206 57866 15258
rect 57866 15206 57912 15258
rect 57616 15204 57672 15206
rect 57696 15204 57752 15206
rect 57776 15204 57832 15206
rect 57856 15204 57912 15206
rect 58530 14764 58532 14784
rect 58532 14764 58584 14784
rect 58584 14764 58586 14784
rect 58530 14728 58586 14764
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 21956 14714 22012 14716
rect 22036 14714 22092 14716
rect 22116 14714 22172 14716
rect 22196 14714 22252 14716
rect 21956 14662 22002 14714
rect 22002 14662 22012 14714
rect 22036 14662 22066 14714
rect 22066 14662 22078 14714
rect 22078 14662 22092 14714
rect 22116 14662 22130 14714
rect 22130 14662 22142 14714
rect 22142 14662 22172 14714
rect 22196 14662 22206 14714
rect 22206 14662 22252 14714
rect 21956 14660 22012 14662
rect 22036 14660 22092 14662
rect 22116 14660 22172 14662
rect 22196 14660 22252 14662
rect 26956 14714 27012 14716
rect 27036 14714 27092 14716
rect 27116 14714 27172 14716
rect 27196 14714 27252 14716
rect 26956 14662 27002 14714
rect 27002 14662 27012 14714
rect 27036 14662 27066 14714
rect 27066 14662 27078 14714
rect 27078 14662 27092 14714
rect 27116 14662 27130 14714
rect 27130 14662 27142 14714
rect 27142 14662 27172 14714
rect 27196 14662 27206 14714
rect 27206 14662 27252 14714
rect 26956 14660 27012 14662
rect 27036 14660 27092 14662
rect 27116 14660 27172 14662
rect 27196 14660 27252 14662
rect 31956 14714 32012 14716
rect 32036 14714 32092 14716
rect 32116 14714 32172 14716
rect 32196 14714 32252 14716
rect 31956 14662 32002 14714
rect 32002 14662 32012 14714
rect 32036 14662 32066 14714
rect 32066 14662 32078 14714
rect 32078 14662 32092 14714
rect 32116 14662 32130 14714
rect 32130 14662 32142 14714
rect 32142 14662 32172 14714
rect 32196 14662 32206 14714
rect 32206 14662 32252 14714
rect 31956 14660 32012 14662
rect 32036 14660 32092 14662
rect 32116 14660 32172 14662
rect 32196 14660 32252 14662
rect 36956 14714 37012 14716
rect 37036 14714 37092 14716
rect 37116 14714 37172 14716
rect 37196 14714 37252 14716
rect 36956 14662 37002 14714
rect 37002 14662 37012 14714
rect 37036 14662 37066 14714
rect 37066 14662 37078 14714
rect 37078 14662 37092 14714
rect 37116 14662 37130 14714
rect 37130 14662 37142 14714
rect 37142 14662 37172 14714
rect 37196 14662 37206 14714
rect 37206 14662 37252 14714
rect 36956 14660 37012 14662
rect 37036 14660 37092 14662
rect 37116 14660 37172 14662
rect 37196 14660 37252 14662
rect 41956 14714 42012 14716
rect 42036 14714 42092 14716
rect 42116 14714 42172 14716
rect 42196 14714 42252 14716
rect 41956 14662 42002 14714
rect 42002 14662 42012 14714
rect 42036 14662 42066 14714
rect 42066 14662 42078 14714
rect 42078 14662 42092 14714
rect 42116 14662 42130 14714
rect 42130 14662 42142 14714
rect 42142 14662 42172 14714
rect 42196 14662 42206 14714
rect 42206 14662 42252 14714
rect 41956 14660 42012 14662
rect 42036 14660 42092 14662
rect 42116 14660 42172 14662
rect 42196 14660 42252 14662
rect 46956 14714 47012 14716
rect 47036 14714 47092 14716
rect 47116 14714 47172 14716
rect 47196 14714 47252 14716
rect 46956 14662 47002 14714
rect 47002 14662 47012 14714
rect 47036 14662 47066 14714
rect 47066 14662 47078 14714
rect 47078 14662 47092 14714
rect 47116 14662 47130 14714
rect 47130 14662 47142 14714
rect 47142 14662 47172 14714
rect 47196 14662 47206 14714
rect 47206 14662 47252 14714
rect 46956 14660 47012 14662
rect 47036 14660 47092 14662
rect 47116 14660 47172 14662
rect 47196 14660 47252 14662
rect 51956 14714 52012 14716
rect 52036 14714 52092 14716
rect 52116 14714 52172 14716
rect 52196 14714 52252 14716
rect 51956 14662 52002 14714
rect 52002 14662 52012 14714
rect 52036 14662 52066 14714
rect 52066 14662 52078 14714
rect 52078 14662 52092 14714
rect 52116 14662 52130 14714
rect 52130 14662 52142 14714
rect 52142 14662 52172 14714
rect 52196 14662 52206 14714
rect 52206 14662 52252 14714
rect 51956 14660 52012 14662
rect 52036 14660 52092 14662
rect 52116 14660 52172 14662
rect 52196 14660 52252 14662
rect 56956 14714 57012 14716
rect 57036 14714 57092 14716
rect 57116 14714 57172 14716
rect 57196 14714 57252 14716
rect 56956 14662 57002 14714
rect 57002 14662 57012 14714
rect 57036 14662 57066 14714
rect 57066 14662 57078 14714
rect 57078 14662 57092 14714
rect 57116 14662 57130 14714
rect 57130 14662 57142 14714
rect 57142 14662 57172 14714
rect 57196 14662 57206 14714
rect 57206 14662 57252 14714
rect 56956 14660 57012 14662
rect 57036 14660 57092 14662
rect 57116 14660 57172 14662
rect 57196 14660 57252 14662
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 22616 14170 22672 14172
rect 22696 14170 22752 14172
rect 22776 14170 22832 14172
rect 22856 14170 22912 14172
rect 22616 14118 22662 14170
rect 22662 14118 22672 14170
rect 22696 14118 22726 14170
rect 22726 14118 22738 14170
rect 22738 14118 22752 14170
rect 22776 14118 22790 14170
rect 22790 14118 22802 14170
rect 22802 14118 22832 14170
rect 22856 14118 22866 14170
rect 22866 14118 22912 14170
rect 22616 14116 22672 14118
rect 22696 14116 22752 14118
rect 22776 14116 22832 14118
rect 22856 14116 22912 14118
rect 27616 14170 27672 14172
rect 27696 14170 27752 14172
rect 27776 14170 27832 14172
rect 27856 14170 27912 14172
rect 27616 14118 27662 14170
rect 27662 14118 27672 14170
rect 27696 14118 27726 14170
rect 27726 14118 27738 14170
rect 27738 14118 27752 14170
rect 27776 14118 27790 14170
rect 27790 14118 27802 14170
rect 27802 14118 27832 14170
rect 27856 14118 27866 14170
rect 27866 14118 27912 14170
rect 27616 14116 27672 14118
rect 27696 14116 27752 14118
rect 27776 14116 27832 14118
rect 27856 14116 27912 14118
rect 32616 14170 32672 14172
rect 32696 14170 32752 14172
rect 32776 14170 32832 14172
rect 32856 14170 32912 14172
rect 32616 14118 32662 14170
rect 32662 14118 32672 14170
rect 32696 14118 32726 14170
rect 32726 14118 32738 14170
rect 32738 14118 32752 14170
rect 32776 14118 32790 14170
rect 32790 14118 32802 14170
rect 32802 14118 32832 14170
rect 32856 14118 32866 14170
rect 32866 14118 32912 14170
rect 32616 14116 32672 14118
rect 32696 14116 32752 14118
rect 32776 14116 32832 14118
rect 32856 14116 32912 14118
rect 37616 14170 37672 14172
rect 37696 14170 37752 14172
rect 37776 14170 37832 14172
rect 37856 14170 37912 14172
rect 37616 14118 37662 14170
rect 37662 14118 37672 14170
rect 37696 14118 37726 14170
rect 37726 14118 37738 14170
rect 37738 14118 37752 14170
rect 37776 14118 37790 14170
rect 37790 14118 37802 14170
rect 37802 14118 37832 14170
rect 37856 14118 37866 14170
rect 37866 14118 37912 14170
rect 37616 14116 37672 14118
rect 37696 14116 37752 14118
rect 37776 14116 37832 14118
rect 37856 14116 37912 14118
rect 42616 14170 42672 14172
rect 42696 14170 42752 14172
rect 42776 14170 42832 14172
rect 42856 14170 42912 14172
rect 42616 14118 42662 14170
rect 42662 14118 42672 14170
rect 42696 14118 42726 14170
rect 42726 14118 42738 14170
rect 42738 14118 42752 14170
rect 42776 14118 42790 14170
rect 42790 14118 42802 14170
rect 42802 14118 42832 14170
rect 42856 14118 42866 14170
rect 42866 14118 42912 14170
rect 42616 14116 42672 14118
rect 42696 14116 42752 14118
rect 42776 14116 42832 14118
rect 42856 14116 42912 14118
rect 47616 14170 47672 14172
rect 47696 14170 47752 14172
rect 47776 14170 47832 14172
rect 47856 14170 47912 14172
rect 47616 14118 47662 14170
rect 47662 14118 47672 14170
rect 47696 14118 47726 14170
rect 47726 14118 47738 14170
rect 47738 14118 47752 14170
rect 47776 14118 47790 14170
rect 47790 14118 47802 14170
rect 47802 14118 47832 14170
rect 47856 14118 47866 14170
rect 47866 14118 47912 14170
rect 47616 14116 47672 14118
rect 47696 14116 47752 14118
rect 47776 14116 47832 14118
rect 47856 14116 47912 14118
rect 52616 14170 52672 14172
rect 52696 14170 52752 14172
rect 52776 14170 52832 14172
rect 52856 14170 52912 14172
rect 52616 14118 52662 14170
rect 52662 14118 52672 14170
rect 52696 14118 52726 14170
rect 52726 14118 52738 14170
rect 52738 14118 52752 14170
rect 52776 14118 52790 14170
rect 52790 14118 52802 14170
rect 52802 14118 52832 14170
rect 52856 14118 52866 14170
rect 52866 14118 52912 14170
rect 52616 14116 52672 14118
rect 52696 14116 52752 14118
rect 52776 14116 52832 14118
rect 52856 14116 52912 14118
rect 57616 14170 57672 14172
rect 57696 14170 57752 14172
rect 57776 14170 57832 14172
rect 57856 14170 57912 14172
rect 57616 14118 57662 14170
rect 57662 14118 57672 14170
rect 57696 14118 57726 14170
rect 57726 14118 57738 14170
rect 57738 14118 57752 14170
rect 57776 14118 57790 14170
rect 57790 14118 57802 14170
rect 57802 14118 57832 14170
rect 57856 14118 57866 14170
rect 57866 14118 57912 14170
rect 57616 14116 57672 14118
rect 57696 14116 57752 14118
rect 57776 14116 57832 14118
rect 57856 14116 57912 14118
rect 58530 13912 58586 13968
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 21956 13626 22012 13628
rect 22036 13626 22092 13628
rect 22116 13626 22172 13628
rect 22196 13626 22252 13628
rect 21956 13574 22002 13626
rect 22002 13574 22012 13626
rect 22036 13574 22066 13626
rect 22066 13574 22078 13626
rect 22078 13574 22092 13626
rect 22116 13574 22130 13626
rect 22130 13574 22142 13626
rect 22142 13574 22172 13626
rect 22196 13574 22206 13626
rect 22206 13574 22252 13626
rect 21956 13572 22012 13574
rect 22036 13572 22092 13574
rect 22116 13572 22172 13574
rect 22196 13572 22252 13574
rect 26956 13626 27012 13628
rect 27036 13626 27092 13628
rect 27116 13626 27172 13628
rect 27196 13626 27252 13628
rect 26956 13574 27002 13626
rect 27002 13574 27012 13626
rect 27036 13574 27066 13626
rect 27066 13574 27078 13626
rect 27078 13574 27092 13626
rect 27116 13574 27130 13626
rect 27130 13574 27142 13626
rect 27142 13574 27172 13626
rect 27196 13574 27206 13626
rect 27206 13574 27252 13626
rect 26956 13572 27012 13574
rect 27036 13572 27092 13574
rect 27116 13572 27172 13574
rect 27196 13572 27252 13574
rect 31956 13626 32012 13628
rect 32036 13626 32092 13628
rect 32116 13626 32172 13628
rect 32196 13626 32252 13628
rect 31956 13574 32002 13626
rect 32002 13574 32012 13626
rect 32036 13574 32066 13626
rect 32066 13574 32078 13626
rect 32078 13574 32092 13626
rect 32116 13574 32130 13626
rect 32130 13574 32142 13626
rect 32142 13574 32172 13626
rect 32196 13574 32206 13626
rect 32206 13574 32252 13626
rect 31956 13572 32012 13574
rect 32036 13572 32092 13574
rect 32116 13572 32172 13574
rect 32196 13572 32252 13574
rect 36956 13626 37012 13628
rect 37036 13626 37092 13628
rect 37116 13626 37172 13628
rect 37196 13626 37252 13628
rect 36956 13574 37002 13626
rect 37002 13574 37012 13626
rect 37036 13574 37066 13626
rect 37066 13574 37078 13626
rect 37078 13574 37092 13626
rect 37116 13574 37130 13626
rect 37130 13574 37142 13626
rect 37142 13574 37172 13626
rect 37196 13574 37206 13626
rect 37206 13574 37252 13626
rect 36956 13572 37012 13574
rect 37036 13572 37092 13574
rect 37116 13572 37172 13574
rect 37196 13572 37252 13574
rect 41956 13626 42012 13628
rect 42036 13626 42092 13628
rect 42116 13626 42172 13628
rect 42196 13626 42252 13628
rect 41956 13574 42002 13626
rect 42002 13574 42012 13626
rect 42036 13574 42066 13626
rect 42066 13574 42078 13626
rect 42078 13574 42092 13626
rect 42116 13574 42130 13626
rect 42130 13574 42142 13626
rect 42142 13574 42172 13626
rect 42196 13574 42206 13626
rect 42206 13574 42252 13626
rect 41956 13572 42012 13574
rect 42036 13572 42092 13574
rect 42116 13572 42172 13574
rect 42196 13572 42252 13574
rect 46956 13626 47012 13628
rect 47036 13626 47092 13628
rect 47116 13626 47172 13628
rect 47196 13626 47252 13628
rect 46956 13574 47002 13626
rect 47002 13574 47012 13626
rect 47036 13574 47066 13626
rect 47066 13574 47078 13626
rect 47078 13574 47092 13626
rect 47116 13574 47130 13626
rect 47130 13574 47142 13626
rect 47142 13574 47172 13626
rect 47196 13574 47206 13626
rect 47206 13574 47252 13626
rect 46956 13572 47012 13574
rect 47036 13572 47092 13574
rect 47116 13572 47172 13574
rect 47196 13572 47252 13574
rect 51956 13626 52012 13628
rect 52036 13626 52092 13628
rect 52116 13626 52172 13628
rect 52196 13626 52252 13628
rect 51956 13574 52002 13626
rect 52002 13574 52012 13626
rect 52036 13574 52066 13626
rect 52066 13574 52078 13626
rect 52078 13574 52092 13626
rect 52116 13574 52130 13626
rect 52130 13574 52142 13626
rect 52142 13574 52172 13626
rect 52196 13574 52206 13626
rect 52206 13574 52252 13626
rect 51956 13572 52012 13574
rect 52036 13572 52092 13574
rect 52116 13572 52172 13574
rect 52196 13572 52252 13574
rect 56956 13626 57012 13628
rect 57036 13626 57092 13628
rect 57116 13626 57172 13628
rect 57196 13626 57252 13628
rect 56956 13574 57002 13626
rect 57002 13574 57012 13626
rect 57036 13574 57066 13626
rect 57066 13574 57078 13626
rect 57078 13574 57092 13626
rect 57116 13574 57130 13626
rect 57130 13574 57142 13626
rect 57142 13574 57172 13626
rect 57196 13574 57206 13626
rect 57206 13574 57252 13626
rect 56956 13572 57012 13574
rect 57036 13572 57092 13574
rect 57116 13572 57172 13574
rect 57196 13572 57252 13574
rect 58530 13096 58586 13152
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 22616 13082 22672 13084
rect 22696 13082 22752 13084
rect 22776 13082 22832 13084
rect 22856 13082 22912 13084
rect 22616 13030 22662 13082
rect 22662 13030 22672 13082
rect 22696 13030 22726 13082
rect 22726 13030 22738 13082
rect 22738 13030 22752 13082
rect 22776 13030 22790 13082
rect 22790 13030 22802 13082
rect 22802 13030 22832 13082
rect 22856 13030 22866 13082
rect 22866 13030 22912 13082
rect 22616 13028 22672 13030
rect 22696 13028 22752 13030
rect 22776 13028 22832 13030
rect 22856 13028 22912 13030
rect 27616 13082 27672 13084
rect 27696 13082 27752 13084
rect 27776 13082 27832 13084
rect 27856 13082 27912 13084
rect 27616 13030 27662 13082
rect 27662 13030 27672 13082
rect 27696 13030 27726 13082
rect 27726 13030 27738 13082
rect 27738 13030 27752 13082
rect 27776 13030 27790 13082
rect 27790 13030 27802 13082
rect 27802 13030 27832 13082
rect 27856 13030 27866 13082
rect 27866 13030 27912 13082
rect 27616 13028 27672 13030
rect 27696 13028 27752 13030
rect 27776 13028 27832 13030
rect 27856 13028 27912 13030
rect 32616 13082 32672 13084
rect 32696 13082 32752 13084
rect 32776 13082 32832 13084
rect 32856 13082 32912 13084
rect 32616 13030 32662 13082
rect 32662 13030 32672 13082
rect 32696 13030 32726 13082
rect 32726 13030 32738 13082
rect 32738 13030 32752 13082
rect 32776 13030 32790 13082
rect 32790 13030 32802 13082
rect 32802 13030 32832 13082
rect 32856 13030 32866 13082
rect 32866 13030 32912 13082
rect 32616 13028 32672 13030
rect 32696 13028 32752 13030
rect 32776 13028 32832 13030
rect 32856 13028 32912 13030
rect 37616 13082 37672 13084
rect 37696 13082 37752 13084
rect 37776 13082 37832 13084
rect 37856 13082 37912 13084
rect 37616 13030 37662 13082
rect 37662 13030 37672 13082
rect 37696 13030 37726 13082
rect 37726 13030 37738 13082
rect 37738 13030 37752 13082
rect 37776 13030 37790 13082
rect 37790 13030 37802 13082
rect 37802 13030 37832 13082
rect 37856 13030 37866 13082
rect 37866 13030 37912 13082
rect 37616 13028 37672 13030
rect 37696 13028 37752 13030
rect 37776 13028 37832 13030
rect 37856 13028 37912 13030
rect 42616 13082 42672 13084
rect 42696 13082 42752 13084
rect 42776 13082 42832 13084
rect 42856 13082 42912 13084
rect 42616 13030 42662 13082
rect 42662 13030 42672 13082
rect 42696 13030 42726 13082
rect 42726 13030 42738 13082
rect 42738 13030 42752 13082
rect 42776 13030 42790 13082
rect 42790 13030 42802 13082
rect 42802 13030 42832 13082
rect 42856 13030 42866 13082
rect 42866 13030 42912 13082
rect 42616 13028 42672 13030
rect 42696 13028 42752 13030
rect 42776 13028 42832 13030
rect 42856 13028 42912 13030
rect 47616 13082 47672 13084
rect 47696 13082 47752 13084
rect 47776 13082 47832 13084
rect 47856 13082 47912 13084
rect 47616 13030 47662 13082
rect 47662 13030 47672 13082
rect 47696 13030 47726 13082
rect 47726 13030 47738 13082
rect 47738 13030 47752 13082
rect 47776 13030 47790 13082
rect 47790 13030 47802 13082
rect 47802 13030 47832 13082
rect 47856 13030 47866 13082
rect 47866 13030 47912 13082
rect 47616 13028 47672 13030
rect 47696 13028 47752 13030
rect 47776 13028 47832 13030
rect 47856 13028 47912 13030
rect 52616 13082 52672 13084
rect 52696 13082 52752 13084
rect 52776 13082 52832 13084
rect 52856 13082 52912 13084
rect 52616 13030 52662 13082
rect 52662 13030 52672 13082
rect 52696 13030 52726 13082
rect 52726 13030 52738 13082
rect 52738 13030 52752 13082
rect 52776 13030 52790 13082
rect 52790 13030 52802 13082
rect 52802 13030 52832 13082
rect 52856 13030 52866 13082
rect 52866 13030 52912 13082
rect 52616 13028 52672 13030
rect 52696 13028 52752 13030
rect 52776 13028 52832 13030
rect 52856 13028 52912 13030
rect 57616 13082 57672 13084
rect 57696 13082 57752 13084
rect 57776 13082 57832 13084
rect 57856 13082 57912 13084
rect 57616 13030 57662 13082
rect 57662 13030 57672 13082
rect 57696 13030 57726 13082
rect 57726 13030 57738 13082
rect 57738 13030 57752 13082
rect 57776 13030 57790 13082
rect 57790 13030 57802 13082
rect 57802 13030 57832 13082
rect 57856 13030 57866 13082
rect 57866 13030 57912 13082
rect 57616 13028 57672 13030
rect 57696 13028 57752 13030
rect 57776 13028 57832 13030
rect 57856 13028 57912 13030
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 21956 12538 22012 12540
rect 22036 12538 22092 12540
rect 22116 12538 22172 12540
rect 22196 12538 22252 12540
rect 21956 12486 22002 12538
rect 22002 12486 22012 12538
rect 22036 12486 22066 12538
rect 22066 12486 22078 12538
rect 22078 12486 22092 12538
rect 22116 12486 22130 12538
rect 22130 12486 22142 12538
rect 22142 12486 22172 12538
rect 22196 12486 22206 12538
rect 22206 12486 22252 12538
rect 21956 12484 22012 12486
rect 22036 12484 22092 12486
rect 22116 12484 22172 12486
rect 22196 12484 22252 12486
rect 26956 12538 27012 12540
rect 27036 12538 27092 12540
rect 27116 12538 27172 12540
rect 27196 12538 27252 12540
rect 26956 12486 27002 12538
rect 27002 12486 27012 12538
rect 27036 12486 27066 12538
rect 27066 12486 27078 12538
rect 27078 12486 27092 12538
rect 27116 12486 27130 12538
rect 27130 12486 27142 12538
rect 27142 12486 27172 12538
rect 27196 12486 27206 12538
rect 27206 12486 27252 12538
rect 26956 12484 27012 12486
rect 27036 12484 27092 12486
rect 27116 12484 27172 12486
rect 27196 12484 27252 12486
rect 31956 12538 32012 12540
rect 32036 12538 32092 12540
rect 32116 12538 32172 12540
rect 32196 12538 32252 12540
rect 31956 12486 32002 12538
rect 32002 12486 32012 12538
rect 32036 12486 32066 12538
rect 32066 12486 32078 12538
rect 32078 12486 32092 12538
rect 32116 12486 32130 12538
rect 32130 12486 32142 12538
rect 32142 12486 32172 12538
rect 32196 12486 32206 12538
rect 32206 12486 32252 12538
rect 31956 12484 32012 12486
rect 32036 12484 32092 12486
rect 32116 12484 32172 12486
rect 32196 12484 32252 12486
rect 36956 12538 37012 12540
rect 37036 12538 37092 12540
rect 37116 12538 37172 12540
rect 37196 12538 37252 12540
rect 36956 12486 37002 12538
rect 37002 12486 37012 12538
rect 37036 12486 37066 12538
rect 37066 12486 37078 12538
rect 37078 12486 37092 12538
rect 37116 12486 37130 12538
rect 37130 12486 37142 12538
rect 37142 12486 37172 12538
rect 37196 12486 37206 12538
rect 37206 12486 37252 12538
rect 36956 12484 37012 12486
rect 37036 12484 37092 12486
rect 37116 12484 37172 12486
rect 37196 12484 37252 12486
rect 41956 12538 42012 12540
rect 42036 12538 42092 12540
rect 42116 12538 42172 12540
rect 42196 12538 42252 12540
rect 41956 12486 42002 12538
rect 42002 12486 42012 12538
rect 42036 12486 42066 12538
rect 42066 12486 42078 12538
rect 42078 12486 42092 12538
rect 42116 12486 42130 12538
rect 42130 12486 42142 12538
rect 42142 12486 42172 12538
rect 42196 12486 42206 12538
rect 42206 12486 42252 12538
rect 41956 12484 42012 12486
rect 42036 12484 42092 12486
rect 42116 12484 42172 12486
rect 42196 12484 42252 12486
rect 46956 12538 47012 12540
rect 47036 12538 47092 12540
rect 47116 12538 47172 12540
rect 47196 12538 47252 12540
rect 46956 12486 47002 12538
rect 47002 12486 47012 12538
rect 47036 12486 47066 12538
rect 47066 12486 47078 12538
rect 47078 12486 47092 12538
rect 47116 12486 47130 12538
rect 47130 12486 47142 12538
rect 47142 12486 47172 12538
rect 47196 12486 47206 12538
rect 47206 12486 47252 12538
rect 46956 12484 47012 12486
rect 47036 12484 47092 12486
rect 47116 12484 47172 12486
rect 47196 12484 47252 12486
rect 51956 12538 52012 12540
rect 52036 12538 52092 12540
rect 52116 12538 52172 12540
rect 52196 12538 52252 12540
rect 51956 12486 52002 12538
rect 52002 12486 52012 12538
rect 52036 12486 52066 12538
rect 52066 12486 52078 12538
rect 52078 12486 52092 12538
rect 52116 12486 52130 12538
rect 52130 12486 52142 12538
rect 52142 12486 52172 12538
rect 52196 12486 52206 12538
rect 52206 12486 52252 12538
rect 51956 12484 52012 12486
rect 52036 12484 52092 12486
rect 52116 12484 52172 12486
rect 52196 12484 52252 12486
rect 56956 12538 57012 12540
rect 57036 12538 57092 12540
rect 57116 12538 57172 12540
rect 57196 12538 57252 12540
rect 56956 12486 57002 12538
rect 57002 12486 57012 12538
rect 57036 12486 57066 12538
rect 57066 12486 57078 12538
rect 57078 12486 57092 12538
rect 57116 12486 57130 12538
rect 57130 12486 57142 12538
rect 57142 12486 57172 12538
rect 57196 12486 57206 12538
rect 57206 12486 57252 12538
rect 56956 12484 57012 12486
rect 57036 12484 57092 12486
rect 57116 12484 57172 12486
rect 57196 12484 57252 12486
rect 58530 12280 58586 12336
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 22616 11994 22672 11996
rect 22696 11994 22752 11996
rect 22776 11994 22832 11996
rect 22856 11994 22912 11996
rect 22616 11942 22662 11994
rect 22662 11942 22672 11994
rect 22696 11942 22726 11994
rect 22726 11942 22738 11994
rect 22738 11942 22752 11994
rect 22776 11942 22790 11994
rect 22790 11942 22802 11994
rect 22802 11942 22832 11994
rect 22856 11942 22866 11994
rect 22866 11942 22912 11994
rect 22616 11940 22672 11942
rect 22696 11940 22752 11942
rect 22776 11940 22832 11942
rect 22856 11940 22912 11942
rect 27616 11994 27672 11996
rect 27696 11994 27752 11996
rect 27776 11994 27832 11996
rect 27856 11994 27912 11996
rect 27616 11942 27662 11994
rect 27662 11942 27672 11994
rect 27696 11942 27726 11994
rect 27726 11942 27738 11994
rect 27738 11942 27752 11994
rect 27776 11942 27790 11994
rect 27790 11942 27802 11994
rect 27802 11942 27832 11994
rect 27856 11942 27866 11994
rect 27866 11942 27912 11994
rect 27616 11940 27672 11942
rect 27696 11940 27752 11942
rect 27776 11940 27832 11942
rect 27856 11940 27912 11942
rect 32616 11994 32672 11996
rect 32696 11994 32752 11996
rect 32776 11994 32832 11996
rect 32856 11994 32912 11996
rect 32616 11942 32662 11994
rect 32662 11942 32672 11994
rect 32696 11942 32726 11994
rect 32726 11942 32738 11994
rect 32738 11942 32752 11994
rect 32776 11942 32790 11994
rect 32790 11942 32802 11994
rect 32802 11942 32832 11994
rect 32856 11942 32866 11994
rect 32866 11942 32912 11994
rect 32616 11940 32672 11942
rect 32696 11940 32752 11942
rect 32776 11940 32832 11942
rect 32856 11940 32912 11942
rect 37616 11994 37672 11996
rect 37696 11994 37752 11996
rect 37776 11994 37832 11996
rect 37856 11994 37912 11996
rect 37616 11942 37662 11994
rect 37662 11942 37672 11994
rect 37696 11942 37726 11994
rect 37726 11942 37738 11994
rect 37738 11942 37752 11994
rect 37776 11942 37790 11994
rect 37790 11942 37802 11994
rect 37802 11942 37832 11994
rect 37856 11942 37866 11994
rect 37866 11942 37912 11994
rect 37616 11940 37672 11942
rect 37696 11940 37752 11942
rect 37776 11940 37832 11942
rect 37856 11940 37912 11942
rect 42616 11994 42672 11996
rect 42696 11994 42752 11996
rect 42776 11994 42832 11996
rect 42856 11994 42912 11996
rect 42616 11942 42662 11994
rect 42662 11942 42672 11994
rect 42696 11942 42726 11994
rect 42726 11942 42738 11994
rect 42738 11942 42752 11994
rect 42776 11942 42790 11994
rect 42790 11942 42802 11994
rect 42802 11942 42832 11994
rect 42856 11942 42866 11994
rect 42866 11942 42912 11994
rect 42616 11940 42672 11942
rect 42696 11940 42752 11942
rect 42776 11940 42832 11942
rect 42856 11940 42912 11942
rect 47616 11994 47672 11996
rect 47696 11994 47752 11996
rect 47776 11994 47832 11996
rect 47856 11994 47912 11996
rect 47616 11942 47662 11994
rect 47662 11942 47672 11994
rect 47696 11942 47726 11994
rect 47726 11942 47738 11994
rect 47738 11942 47752 11994
rect 47776 11942 47790 11994
rect 47790 11942 47802 11994
rect 47802 11942 47832 11994
rect 47856 11942 47866 11994
rect 47866 11942 47912 11994
rect 47616 11940 47672 11942
rect 47696 11940 47752 11942
rect 47776 11940 47832 11942
rect 47856 11940 47912 11942
rect 52616 11994 52672 11996
rect 52696 11994 52752 11996
rect 52776 11994 52832 11996
rect 52856 11994 52912 11996
rect 52616 11942 52662 11994
rect 52662 11942 52672 11994
rect 52696 11942 52726 11994
rect 52726 11942 52738 11994
rect 52738 11942 52752 11994
rect 52776 11942 52790 11994
rect 52790 11942 52802 11994
rect 52802 11942 52832 11994
rect 52856 11942 52866 11994
rect 52866 11942 52912 11994
rect 52616 11940 52672 11942
rect 52696 11940 52752 11942
rect 52776 11940 52832 11942
rect 52856 11940 52912 11942
rect 57616 11994 57672 11996
rect 57696 11994 57752 11996
rect 57776 11994 57832 11996
rect 57856 11994 57912 11996
rect 57616 11942 57662 11994
rect 57662 11942 57672 11994
rect 57696 11942 57726 11994
rect 57726 11942 57738 11994
rect 57738 11942 57752 11994
rect 57776 11942 57790 11994
rect 57790 11942 57802 11994
rect 57802 11942 57832 11994
rect 57856 11942 57866 11994
rect 57866 11942 57912 11994
rect 57616 11940 57672 11942
rect 57696 11940 57752 11942
rect 57776 11940 57832 11942
rect 57856 11940 57912 11942
rect 58530 11500 58532 11520
rect 58532 11500 58584 11520
rect 58584 11500 58586 11520
rect 58530 11464 58586 11500
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 21956 11450 22012 11452
rect 22036 11450 22092 11452
rect 22116 11450 22172 11452
rect 22196 11450 22252 11452
rect 21956 11398 22002 11450
rect 22002 11398 22012 11450
rect 22036 11398 22066 11450
rect 22066 11398 22078 11450
rect 22078 11398 22092 11450
rect 22116 11398 22130 11450
rect 22130 11398 22142 11450
rect 22142 11398 22172 11450
rect 22196 11398 22206 11450
rect 22206 11398 22252 11450
rect 21956 11396 22012 11398
rect 22036 11396 22092 11398
rect 22116 11396 22172 11398
rect 22196 11396 22252 11398
rect 26956 11450 27012 11452
rect 27036 11450 27092 11452
rect 27116 11450 27172 11452
rect 27196 11450 27252 11452
rect 26956 11398 27002 11450
rect 27002 11398 27012 11450
rect 27036 11398 27066 11450
rect 27066 11398 27078 11450
rect 27078 11398 27092 11450
rect 27116 11398 27130 11450
rect 27130 11398 27142 11450
rect 27142 11398 27172 11450
rect 27196 11398 27206 11450
rect 27206 11398 27252 11450
rect 26956 11396 27012 11398
rect 27036 11396 27092 11398
rect 27116 11396 27172 11398
rect 27196 11396 27252 11398
rect 31956 11450 32012 11452
rect 32036 11450 32092 11452
rect 32116 11450 32172 11452
rect 32196 11450 32252 11452
rect 31956 11398 32002 11450
rect 32002 11398 32012 11450
rect 32036 11398 32066 11450
rect 32066 11398 32078 11450
rect 32078 11398 32092 11450
rect 32116 11398 32130 11450
rect 32130 11398 32142 11450
rect 32142 11398 32172 11450
rect 32196 11398 32206 11450
rect 32206 11398 32252 11450
rect 31956 11396 32012 11398
rect 32036 11396 32092 11398
rect 32116 11396 32172 11398
rect 32196 11396 32252 11398
rect 36956 11450 37012 11452
rect 37036 11450 37092 11452
rect 37116 11450 37172 11452
rect 37196 11450 37252 11452
rect 36956 11398 37002 11450
rect 37002 11398 37012 11450
rect 37036 11398 37066 11450
rect 37066 11398 37078 11450
rect 37078 11398 37092 11450
rect 37116 11398 37130 11450
rect 37130 11398 37142 11450
rect 37142 11398 37172 11450
rect 37196 11398 37206 11450
rect 37206 11398 37252 11450
rect 36956 11396 37012 11398
rect 37036 11396 37092 11398
rect 37116 11396 37172 11398
rect 37196 11396 37252 11398
rect 41956 11450 42012 11452
rect 42036 11450 42092 11452
rect 42116 11450 42172 11452
rect 42196 11450 42252 11452
rect 41956 11398 42002 11450
rect 42002 11398 42012 11450
rect 42036 11398 42066 11450
rect 42066 11398 42078 11450
rect 42078 11398 42092 11450
rect 42116 11398 42130 11450
rect 42130 11398 42142 11450
rect 42142 11398 42172 11450
rect 42196 11398 42206 11450
rect 42206 11398 42252 11450
rect 41956 11396 42012 11398
rect 42036 11396 42092 11398
rect 42116 11396 42172 11398
rect 42196 11396 42252 11398
rect 46956 11450 47012 11452
rect 47036 11450 47092 11452
rect 47116 11450 47172 11452
rect 47196 11450 47252 11452
rect 46956 11398 47002 11450
rect 47002 11398 47012 11450
rect 47036 11398 47066 11450
rect 47066 11398 47078 11450
rect 47078 11398 47092 11450
rect 47116 11398 47130 11450
rect 47130 11398 47142 11450
rect 47142 11398 47172 11450
rect 47196 11398 47206 11450
rect 47206 11398 47252 11450
rect 46956 11396 47012 11398
rect 47036 11396 47092 11398
rect 47116 11396 47172 11398
rect 47196 11396 47252 11398
rect 51956 11450 52012 11452
rect 52036 11450 52092 11452
rect 52116 11450 52172 11452
rect 52196 11450 52252 11452
rect 51956 11398 52002 11450
rect 52002 11398 52012 11450
rect 52036 11398 52066 11450
rect 52066 11398 52078 11450
rect 52078 11398 52092 11450
rect 52116 11398 52130 11450
rect 52130 11398 52142 11450
rect 52142 11398 52172 11450
rect 52196 11398 52206 11450
rect 52206 11398 52252 11450
rect 51956 11396 52012 11398
rect 52036 11396 52092 11398
rect 52116 11396 52172 11398
rect 52196 11396 52252 11398
rect 56956 11450 57012 11452
rect 57036 11450 57092 11452
rect 57116 11450 57172 11452
rect 57196 11450 57252 11452
rect 56956 11398 57002 11450
rect 57002 11398 57012 11450
rect 57036 11398 57066 11450
rect 57066 11398 57078 11450
rect 57078 11398 57092 11450
rect 57116 11398 57130 11450
rect 57130 11398 57142 11450
rect 57142 11398 57172 11450
rect 57196 11398 57206 11450
rect 57206 11398 57252 11450
rect 56956 11396 57012 11398
rect 57036 11396 57092 11398
rect 57116 11396 57172 11398
rect 57196 11396 57252 11398
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 22616 10906 22672 10908
rect 22696 10906 22752 10908
rect 22776 10906 22832 10908
rect 22856 10906 22912 10908
rect 22616 10854 22662 10906
rect 22662 10854 22672 10906
rect 22696 10854 22726 10906
rect 22726 10854 22738 10906
rect 22738 10854 22752 10906
rect 22776 10854 22790 10906
rect 22790 10854 22802 10906
rect 22802 10854 22832 10906
rect 22856 10854 22866 10906
rect 22866 10854 22912 10906
rect 22616 10852 22672 10854
rect 22696 10852 22752 10854
rect 22776 10852 22832 10854
rect 22856 10852 22912 10854
rect 27616 10906 27672 10908
rect 27696 10906 27752 10908
rect 27776 10906 27832 10908
rect 27856 10906 27912 10908
rect 27616 10854 27662 10906
rect 27662 10854 27672 10906
rect 27696 10854 27726 10906
rect 27726 10854 27738 10906
rect 27738 10854 27752 10906
rect 27776 10854 27790 10906
rect 27790 10854 27802 10906
rect 27802 10854 27832 10906
rect 27856 10854 27866 10906
rect 27866 10854 27912 10906
rect 27616 10852 27672 10854
rect 27696 10852 27752 10854
rect 27776 10852 27832 10854
rect 27856 10852 27912 10854
rect 32616 10906 32672 10908
rect 32696 10906 32752 10908
rect 32776 10906 32832 10908
rect 32856 10906 32912 10908
rect 32616 10854 32662 10906
rect 32662 10854 32672 10906
rect 32696 10854 32726 10906
rect 32726 10854 32738 10906
rect 32738 10854 32752 10906
rect 32776 10854 32790 10906
rect 32790 10854 32802 10906
rect 32802 10854 32832 10906
rect 32856 10854 32866 10906
rect 32866 10854 32912 10906
rect 32616 10852 32672 10854
rect 32696 10852 32752 10854
rect 32776 10852 32832 10854
rect 32856 10852 32912 10854
rect 37616 10906 37672 10908
rect 37696 10906 37752 10908
rect 37776 10906 37832 10908
rect 37856 10906 37912 10908
rect 37616 10854 37662 10906
rect 37662 10854 37672 10906
rect 37696 10854 37726 10906
rect 37726 10854 37738 10906
rect 37738 10854 37752 10906
rect 37776 10854 37790 10906
rect 37790 10854 37802 10906
rect 37802 10854 37832 10906
rect 37856 10854 37866 10906
rect 37866 10854 37912 10906
rect 37616 10852 37672 10854
rect 37696 10852 37752 10854
rect 37776 10852 37832 10854
rect 37856 10852 37912 10854
rect 42616 10906 42672 10908
rect 42696 10906 42752 10908
rect 42776 10906 42832 10908
rect 42856 10906 42912 10908
rect 42616 10854 42662 10906
rect 42662 10854 42672 10906
rect 42696 10854 42726 10906
rect 42726 10854 42738 10906
rect 42738 10854 42752 10906
rect 42776 10854 42790 10906
rect 42790 10854 42802 10906
rect 42802 10854 42832 10906
rect 42856 10854 42866 10906
rect 42866 10854 42912 10906
rect 42616 10852 42672 10854
rect 42696 10852 42752 10854
rect 42776 10852 42832 10854
rect 42856 10852 42912 10854
rect 47616 10906 47672 10908
rect 47696 10906 47752 10908
rect 47776 10906 47832 10908
rect 47856 10906 47912 10908
rect 47616 10854 47662 10906
rect 47662 10854 47672 10906
rect 47696 10854 47726 10906
rect 47726 10854 47738 10906
rect 47738 10854 47752 10906
rect 47776 10854 47790 10906
rect 47790 10854 47802 10906
rect 47802 10854 47832 10906
rect 47856 10854 47866 10906
rect 47866 10854 47912 10906
rect 47616 10852 47672 10854
rect 47696 10852 47752 10854
rect 47776 10852 47832 10854
rect 47856 10852 47912 10854
rect 52616 10906 52672 10908
rect 52696 10906 52752 10908
rect 52776 10906 52832 10908
rect 52856 10906 52912 10908
rect 52616 10854 52662 10906
rect 52662 10854 52672 10906
rect 52696 10854 52726 10906
rect 52726 10854 52738 10906
rect 52738 10854 52752 10906
rect 52776 10854 52790 10906
rect 52790 10854 52802 10906
rect 52802 10854 52832 10906
rect 52856 10854 52866 10906
rect 52866 10854 52912 10906
rect 52616 10852 52672 10854
rect 52696 10852 52752 10854
rect 52776 10852 52832 10854
rect 52856 10852 52912 10854
rect 57616 10906 57672 10908
rect 57696 10906 57752 10908
rect 57776 10906 57832 10908
rect 57856 10906 57912 10908
rect 57616 10854 57662 10906
rect 57662 10854 57672 10906
rect 57696 10854 57726 10906
rect 57726 10854 57738 10906
rect 57738 10854 57752 10906
rect 57776 10854 57790 10906
rect 57790 10854 57802 10906
rect 57802 10854 57832 10906
rect 57856 10854 57866 10906
rect 57866 10854 57912 10906
rect 57616 10852 57672 10854
rect 57696 10852 57752 10854
rect 57776 10852 57832 10854
rect 57856 10852 57912 10854
rect 58530 10648 58586 10704
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 21956 10362 22012 10364
rect 22036 10362 22092 10364
rect 22116 10362 22172 10364
rect 22196 10362 22252 10364
rect 21956 10310 22002 10362
rect 22002 10310 22012 10362
rect 22036 10310 22066 10362
rect 22066 10310 22078 10362
rect 22078 10310 22092 10362
rect 22116 10310 22130 10362
rect 22130 10310 22142 10362
rect 22142 10310 22172 10362
rect 22196 10310 22206 10362
rect 22206 10310 22252 10362
rect 21956 10308 22012 10310
rect 22036 10308 22092 10310
rect 22116 10308 22172 10310
rect 22196 10308 22252 10310
rect 26956 10362 27012 10364
rect 27036 10362 27092 10364
rect 27116 10362 27172 10364
rect 27196 10362 27252 10364
rect 26956 10310 27002 10362
rect 27002 10310 27012 10362
rect 27036 10310 27066 10362
rect 27066 10310 27078 10362
rect 27078 10310 27092 10362
rect 27116 10310 27130 10362
rect 27130 10310 27142 10362
rect 27142 10310 27172 10362
rect 27196 10310 27206 10362
rect 27206 10310 27252 10362
rect 26956 10308 27012 10310
rect 27036 10308 27092 10310
rect 27116 10308 27172 10310
rect 27196 10308 27252 10310
rect 31956 10362 32012 10364
rect 32036 10362 32092 10364
rect 32116 10362 32172 10364
rect 32196 10362 32252 10364
rect 31956 10310 32002 10362
rect 32002 10310 32012 10362
rect 32036 10310 32066 10362
rect 32066 10310 32078 10362
rect 32078 10310 32092 10362
rect 32116 10310 32130 10362
rect 32130 10310 32142 10362
rect 32142 10310 32172 10362
rect 32196 10310 32206 10362
rect 32206 10310 32252 10362
rect 31956 10308 32012 10310
rect 32036 10308 32092 10310
rect 32116 10308 32172 10310
rect 32196 10308 32252 10310
rect 36956 10362 37012 10364
rect 37036 10362 37092 10364
rect 37116 10362 37172 10364
rect 37196 10362 37252 10364
rect 36956 10310 37002 10362
rect 37002 10310 37012 10362
rect 37036 10310 37066 10362
rect 37066 10310 37078 10362
rect 37078 10310 37092 10362
rect 37116 10310 37130 10362
rect 37130 10310 37142 10362
rect 37142 10310 37172 10362
rect 37196 10310 37206 10362
rect 37206 10310 37252 10362
rect 36956 10308 37012 10310
rect 37036 10308 37092 10310
rect 37116 10308 37172 10310
rect 37196 10308 37252 10310
rect 41956 10362 42012 10364
rect 42036 10362 42092 10364
rect 42116 10362 42172 10364
rect 42196 10362 42252 10364
rect 41956 10310 42002 10362
rect 42002 10310 42012 10362
rect 42036 10310 42066 10362
rect 42066 10310 42078 10362
rect 42078 10310 42092 10362
rect 42116 10310 42130 10362
rect 42130 10310 42142 10362
rect 42142 10310 42172 10362
rect 42196 10310 42206 10362
rect 42206 10310 42252 10362
rect 41956 10308 42012 10310
rect 42036 10308 42092 10310
rect 42116 10308 42172 10310
rect 42196 10308 42252 10310
rect 46956 10362 47012 10364
rect 47036 10362 47092 10364
rect 47116 10362 47172 10364
rect 47196 10362 47252 10364
rect 46956 10310 47002 10362
rect 47002 10310 47012 10362
rect 47036 10310 47066 10362
rect 47066 10310 47078 10362
rect 47078 10310 47092 10362
rect 47116 10310 47130 10362
rect 47130 10310 47142 10362
rect 47142 10310 47172 10362
rect 47196 10310 47206 10362
rect 47206 10310 47252 10362
rect 46956 10308 47012 10310
rect 47036 10308 47092 10310
rect 47116 10308 47172 10310
rect 47196 10308 47252 10310
rect 51956 10362 52012 10364
rect 52036 10362 52092 10364
rect 52116 10362 52172 10364
rect 52196 10362 52252 10364
rect 51956 10310 52002 10362
rect 52002 10310 52012 10362
rect 52036 10310 52066 10362
rect 52066 10310 52078 10362
rect 52078 10310 52092 10362
rect 52116 10310 52130 10362
rect 52130 10310 52142 10362
rect 52142 10310 52172 10362
rect 52196 10310 52206 10362
rect 52206 10310 52252 10362
rect 51956 10308 52012 10310
rect 52036 10308 52092 10310
rect 52116 10308 52172 10310
rect 52196 10308 52252 10310
rect 56956 10362 57012 10364
rect 57036 10362 57092 10364
rect 57116 10362 57172 10364
rect 57196 10362 57252 10364
rect 56956 10310 57002 10362
rect 57002 10310 57012 10362
rect 57036 10310 57066 10362
rect 57066 10310 57078 10362
rect 57078 10310 57092 10362
rect 57116 10310 57130 10362
rect 57130 10310 57142 10362
rect 57142 10310 57172 10362
rect 57196 10310 57206 10362
rect 57206 10310 57252 10362
rect 56956 10308 57012 10310
rect 57036 10308 57092 10310
rect 57116 10308 57172 10310
rect 57196 10308 57252 10310
rect 58530 9832 58586 9888
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 22616 9818 22672 9820
rect 22696 9818 22752 9820
rect 22776 9818 22832 9820
rect 22856 9818 22912 9820
rect 22616 9766 22662 9818
rect 22662 9766 22672 9818
rect 22696 9766 22726 9818
rect 22726 9766 22738 9818
rect 22738 9766 22752 9818
rect 22776 9766 22790 9818
rect 22790 9766 22802 9818
rect 22802 9766 22832 9818
rect 22856 9766 22866 9818
rect 22866 9766 22912 9818
rect 22616 9764 22672 9766
rect 22696 9764 22752 9766
rect 22776 9764 22832 9766
rect 22856 9764 22912 9766
rect 27616 9818 27672 9820
rect 27696 9818 27752 9820
rect 27776 9818 27832 9820
rect 27856 9818 27912 9820
rect 27616 9766 27662 9818
rect 27662 9766 27672 9818
rect 27696 9766 27726 9818
rect 27726 9766 27738 9818
rect 27738 9766 27752 9818
rect 27776 9766 27790 9818
rect 27790 9766 27802 9818
rect 27802 9766 27832 9818
rect 27856 9766 27866 9818
rect 27866 9766 27912 9818
rect 27616 9764 27672 9766
rect 27696 9764 27752 9766
rect 27776 9764 27832 9766
rect 27856 9764 27912 9766
rect 32616 9818 32672 9820
rect 32696 9818 32752 9820
rect 32776 9818 32832 9820
rect 32856 9818 32912 9820
rect 32616 9766 32662 9818
rect 32662 9766 32672 9818
rect 32696 9766 32726 9818
rect 32726 9766 32738 9818
rect 32738 9766 32752 9818
rect 32776 9766 32790 9818
rect 32790 9766 32802 9818
rect 32802 9766 32832 9818
rect 32856 9766 32866 9818
rect 32866 9766 32912 9818
rect 32616 9764 32672 9766
rect 32696 9764 32752 9766
rect 32776 9764 32832 9766
rect 32856 9764 32912 9766
rect 37616 9818 37672 9820
rect 37696 9818 37752 9820
rect 37776 9818 37832 9820
rect 37856 9818 37912 9820
rect 37616 9766 37662 9818
rect 37662 9766 37672 9818
rect 37696 9766 37726 9818
rect 37726 9766 37738 9818
rect 37738 9766 37752 9818
rect 37776 9766 37790 9818
rect 37790 9766 37802 9818
rect 37802 9766 37832 9818
rect 37856 9766 37866 9818
rect 37866 9766 37912 9818
rect 37616 9764 37672 9766
rect 37696 9764 37752 9766
rect 37776 9764 37832 9766
rect 37856 9764 37912 9766
rect 42616 9818 42672 9820
rect 42696 9818 42752 9820
rect 42776 9818 42832 9820
rect 42856 9818 42912 9820
rect 42616 9766 42662 9818
rect 42662 9766 42672 9818
rect 42696 9766 42726 9818
rect 42726 9766 42738 9818
rect 42738 9766 42752 9818
rect 42776 9766 42790 9818
rect 42790 9766 42802 9818
rect 42802 9766 42832 9818
rect 42856 9766 42866 9818
rect 42866 9766 42912 9818
rect 42616 9764 42672 9766
rect 42696 9764 42752 9766
rect 42776 9764 42832 9766
rect 42856 9764 42912 9766
rect 47616 9818 47672 9820
rect 47696 9818 47752 9820
rect 47776 9818 47832 9820
rect 47856 9818 47912 9820
rect 47616 9766 47662 9818
rect 47662 9766 47672 9818
rect 47696 9766 47726 9818
rect 47726 9766 47738 9818
rect 47738 9766 47752 9818
rect 47776 9766 47790 9818
rect 47790 9766 47802 9818
rect 47802 9766 47832 9818
rect 47856 9766 47866 9818
rect 47866 9766 47912 9818
rect 47616 9764 47672 9766
rect 47696 9764 47752 9766
rect 47776 9764 47832 9766
rect 47856 9764 47912 9766
rect 52616 9818 52672 9820
rect 52696 9818 52752 9820
rect 52776 9818 52832 9820
rect 52856 9818 52912 9820
rect 52616 9766 52662 9818
rect 52662 9766 52672 9818
rect 52696 9766 52726 9818
rect 52726 9766 52738 9818
rect 52738 9766 52752 9818
rect 52776 9766 52790 9818
rect 52790 9766 52802 9818
rect 52802 9766 52832 9818
rect 52856 9766 52866 9818
rect 52866 9766 52912 9818
rect 52616 9764 52672 9766
rect 52696 9764 52752 9766
rect 52776 9764 52832 9766
rect 52856 9764 52912 9766
rect 57616 9818 57672 9820
rect 57696 9818 57752 9820
rect 57776 9818 57832 9820
rect 57856 9818 57912 9820
rect 57616 9766 57662 9818
rect 57662 9766 57672 9818
rect 57696 9766 57726 9818
rect 57726 9766 57738 9818
rect 57738 9766 57752 9818
rect 57776 9766 57790 9818
rect 57790 9766 57802 9818
rect 57802 9766 57832 9818
rect 57856 9766 57866 9818
rect 57866 9766 57912 9818
rect 57616 9764 57672 9766
rect 57696 9764 57752 9766
rect 57776 9764 57832 9766
rect 57856 9764 57912 9766
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 21956 9274 22012 9276
rect 22036 9274 22092 9276
rect 22116 9274 22172 9276
rect 22196 9274 22252 9276
rect 21956 9222 22002 9274
rect 22002 9222 22012 9274
rect 22036 9222 22066 9274
rect 22066 9222 22078 9274
rect 22078 9222 22092 9274
rect 22116 9222 22130 9274
rect 22130 9222 22142 9274
rect 22142 9222 22172 9274
rect 22196 9222 22206 9274
rect 22206 9222 22252 9274
rect 21956 9220 22012 9222
rect 22036 9220 22092 9222
rect 22116 9220 22172 9222
rect 22196 9220 22252 9222
rect 26956 9274 27012 9276
rect 27036 9274 27092 9276
rect 27116 9274 27172 9276
rect 27196 9274 27252 9276
rect 26956 9222 27002 9274
rect 27002 9222 27012 9274
rect 27036 9222 27066 9274
rect 27066 9222 27078 9274
rect 27078 9222 27092 9274
rect 27116 9222 27130 9274
rect 27130 9222 27142 9274
rect 27142 9222 27172 9274
rect 27196 9222 27206 9274
rect 27206 9222 27252 9274
rect 26956 9220 27012 9222
rect 27036 9220 27092 9222
rect 27116 9220 27172 9222
rect 27196 9220 27252 9222
rect 31956 9274 32012 9276
rect 32036 9274 32092 9276
rect 32116 9274 32172 9276
rect 32196 9274 32252 9276
rect 31956 9222 32002 9274
rect 32002 9222 32012 9274
rect 32036 9222 32066 9274
rect 32066 9222 32078 9274
rect 32078 9222 32092 9274
rect 32116 9222 32130 9274
rect 32130 9222 32142 9274
rect 32142 9222 32172 9274
rect 32196 9222 32206 9274
rect 32206 9222 32252 9274
rect 31956 9220 32012 9222
rect 32036 9220 32092 9222
rect 32116 9220 32172 9222
rect 32196 9220 32252 9222
rect 36956 9274 37012 9276
rect 37036 9274 37092 9276
rect 37116 9274 37172 9276
rect 37196 9274 37252 9276
rect 36956 9222 37002 9274
rect 37002 9222 37012 9274
rect 37036 9222 37066 9274
rect 37066 9222 37078 9274
rect 37078 9222 37092 9274
rect 37116 9222 37130 9274
rect 37130 9222 37142 9274
rect 37142 9222 37172 9274
rect 37196 9222 37206 9274
rect 37206 9222 37252 9274
rect 36956 9220 37012 9222
rect 37036 9220 37092 9222
rect 37116 9220 37172 9222
rect 37196 9220 37252 9222
rect 41956 9274 42012 9276
rect 42036 9274 42092 9276
rect 42116 9274 42172 9276
rect 42196 9274 42252 9276
rect 41956 9222 42002 9274
rect 42002 9222 42012 9274
rect 42036 9222 42066 9274
rect 42066 9222 42078 9274
rect 42078 9222 42092 9274
rect 42116 9222 42130 9274
rect 42130 9222 42142 9274
rect 42142 9222 42172 9274
rect 42196 9222 42206 9274
rect 42206 9222 42252 9274
rect 41956 9220 42012 9222
rect 42036 9220 42092 9222
rect 42116 9220 42172 9222
rect 42196 9220 42252 9222
rect 46956 9274 47012 9276
rect 47036 9274 47092 9276
rect 47116 9274 47172 9276
rect 47196 9274 47252 9276
rect 46956 9222 47002 9274
rect 47002 9222 47012 9274
rect 47036 9222 47066 9274
rect 47066 9222 47078 9274
rect 47078 9222 47092 9274
rect 47116 9222 47130 9274
rect 47130 9222 47142 9274
rect 47142 9222 47172 9274
rect 47196 9222 47206 9274
rect 47206 9222 47252 9274
rect 46956 9220 47012 9222
rect 47036 9220 47092 9222
rect 47116 9220 47172 9222
rect 47196 9220 47252 9222
rect 51956 9274 52012 9276
rect 52036 9274 52092 9276
rect 52116 9274 52172 9276
rect 52196 9274 52252 9276
rect 51956 9222 52002 9274
rect 52002 9222 52012 9274
rect 52036 9222 52066 9274
rect 52066 9222 52078 9274
rect 52078 9222 52092 9274
rect 52116 9222 52130 9274
rect 52130 9222 52142 9274
rect 52142 9222 52172 9274
rect 52196 9222 52206 9274
rect 52206 9222 52252 9274
rect 51956 9220 52012 9222
rect 52036 9220 52092 9222
rect 52116 9220 52172 9222
rect 52196 9220 52252 9222
rect 56956 9274 57012 9276
rect 57036 9274 57092 9276
rect 57116 9274 57172 9276
rect 57196 9274 57252 9276
rect 56956 9222 57002 9274
rect 57002 9222 57012 9274
rect 57036 9222 57066 9274
rect 57066 9222 57078 9274
rect 57078 9222 57092 9274
rect 57116 9222 57130 9274
rect 57130 9222 57142 9274
rect 57142 9222 57172 9274
rect 57196 9222 57206 9274
rect 57206 9222 57252 9274
rect 56956 9220 57012 9222
rect 57036 9220 57092 9222
rect 57116 9220 57172 9222
rect 57196 9220 57252 9222
rect 58530 9016 58586 9072
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 22616 8730 22672 8732
rect 22696 8730 22752 8732
rect 22776 8730 22832 8732
rect 22856 8730 22912 8732
rect 22616 8678 22662 8730
rect 22662 8678 22672 8730
rect 22696 8678 22726 8730
rect 22726 8678 22738 8730
rect 22738 8678 22752 8730
rect 22776 8678 22790 8730
rect 22790 8678 22802 8730
rect 22802 8678 22832 8730
rect 22856 8678 22866 8730
rect 22866 8678 22912 8730
rect 22616 8676 22672 8678
rect 22696 8676 22752 8678
rect 22776 8676 22832 8678
rect 22856 8676 22912 8678
rect 27616 8730 27672 8732
rect 27696 8730 27752 8732
rect 27776 8730 27832 8732
rect 27856 8730 27912 8732
rect 27616 8678 27662 8730
rect 27662 8678 27672 8730
rect 27696 8678 27726 8730
rect 27726 8678 27738 8730
rect 27738 8678 27752 8730
rect 27776 8678 27790 8730
rect 27790 8678 27802 8730
rect 27802 8678 27832 8730
rect 27856 8678 27866 8730
rect 27866 8678 27912 8730
rect 27616 8676 27672 8678
rect 27696 8676 27752 8678
rect 27776 8676 27832 8678
rect 27856 8676 27912 8678
rect 32616 8730 32672 8732
rect 32696 8730 32752 8732
rect 32776 8730 32832 8732
rect 32856 8730 32912 8732
rect 32616 8678 32662 8730
rect 32662 8678 32672 8730
rect 32696 8678 32726 8730
rect 32726 8678 32738 8730
rect 32738 8678 32752 8730
rect 32776 8678 32790 8730
rect 32790 8678 32802 8730
rect 32802 8678 32832 8730
rect 32856 8678 32866 8730
rect 32866 8678 32912 8730
rect 32616 8676 32672 8678
rect 32696 8676 32752 8678
rect 32776 8676 32832 8678
rect 32856 8676 32912 8678
rect 37616 8730 37672 8732
rect 37696 8730 37752 8732
rect 37776 8730 37832 8732
rect 37856 8730 37912 8732
rect 37616 8678 37662 8730
rect 37662 8678 37672 8730
rect 37696 8678 37726 8730
rect 37726 8678 37738 8730
rect 37738 8678 37752 8730
rect 37776 8678 37790 8730
rect 37790 8678 37802 8730
rect 37802 8678 37832 8730
rect 37856 8678 37866 8730
rect 37866 8678 37912 8730
rect 37616 8676 37672 8678
rect 37696 8676 37752 8678
rect 37776 8676 37832 8678
rect 37856 8676 37912 8678
rect 42616 8730 42672 8732
rect 42696 8730 42752 8732
rect 42776 8730 42832 8732
rect 42856 8730 42912 8732
rect 42616 8678 42662 8730
rect 42662 8678 42672 8730
rect 42696 8678 42726 8730
rect 42726 8678 42738 8730
rect 42738 8678 42752 8730
rect 42776 8678 42790 8730
rect 42790 8678 42802 8730
rect 42802 8678 42832 8730
rect 42856 8678 42866 8730
rect 42866 8678 42912 8730
rect 42616 8676 42672 8678
rect 42696 8676 42752 8678
rect 42776 8676 42832 8678
rect 42856 8676 42912 8678
rect 47616 8730 47672 8732
rect 47696 8730 47752 8732
rect 47776 8730 47832 8732
rect 47856 8730 47912 8732
rect 47616 8678 47662 8730
rect 47662 8678 47672 8730
rect 47696 8678 47726 8730
rect 47726 8678 47738 8730
rect 47738 8678 47752 8730
rect 47776 8678 47790 8730
rect 47790 8678 47802 8730
rect 47802 8678 47832 8730
rect 47856 8678 47866 8730
rect 47866 8678 47912 8730
rect 47616 8676 47672 8678
rect 47696 8676 47752 8678
rect 47776 8676 47832 8678
rect 47856 8676 47912 8678
rect 52616 8730 52672 8732
rect 52696 8730 52752 8732
rect 52776 8730 52832 8732
rect 52856 8730 52912 8732
rect 52616 8678 52662 8730
rect 52662 8678 52672 8730
rect 52696 8678 52726 8730
rect 52726 8678 52738 8730
rect 52738 8678 52752 8730
rect 52776 8678 52790 8730
rect 52790 8678 52802 8730
rect 52802 8678 52832 8730
rect 52856 8678 52866 8730
rect 52866 8678 52912 8730
rect 52616 8676 52672 8678
rect 52696 8676 52752 8678
rect 52776 8676 52832 8678
rect 52856 8676 52912 8678
rect 57616 8730 57672 8732
rect 57696 8730 57752 8732
rect 57776 8730 57832 8732
rect 57856 8730 57912 8732
rect 57616 8678 57662 8730
rect 57662 8678 57672 8730
rect 57696 8678 57726 8730
rect 57726 8678 57738 8730
rect 57738 8678 57752 8730
rect 57776 8678 57790 8730
rect 57790 8678 57802 8730
rect 57802 8678 57832 8730
rect 57856 8678 57866 8730
rect 57866 8678 57912 8730
rect 57616 8676 57672 8678
rect 57696 8676 57752 8678
rect 57776 8676 57832 8678
rect 57856 8676 57912 8678
rect 58530 8200 58586 8256
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 21956 8186 22012 8188
rect 22036 8186 22092 8188
rect 22116 8186 22172 8188
rect 22196 8186 22252 8188
rect 21956 8134 22002 8186
rect 22002 8134 22012 8186
rect 22036 8134 22066 8186
rect 22066 8134 22078 8186
rect 22078 8134 22092 8186
rect 22116 8134 22130 8186
rect 22130 8134 22142 8186
rect 22142 8134 22172 8186
rect 22196 8134 22206 8186
rect 22206 8134 22252 8186
rect 21956 8132 22012 8134
rect 22036 8132 22092 8134
rect 22116 8132 22172 8134
rect 22196 8132 22252 8134
rect 26956 8186 27012 8188
rect 27036 8186 27092 8188
rect 27116 8186 27172 8188
rect 27196 8186 27252 8188
rect 26956 8134 27002 8186
rect 27002 8134 27012 8186
rect 27036 8134 27066 8186
rect 27066 8134 27078 8186
rect 27078 8134 27092 8186
rect 27116 8134 27130 8186
rect 27130 8134 27142 8186
rect 27142 8134 27172 8186
rect 27196 8134 27206 8186
rect 27206 8134 27252 8186
rect 26956 8132 27012 8134
rect 27036 8132 27092 8134
rect 27116 8132 27172 8134
rect 27196 8132 27252 8134
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 36956 8186 37012 8188
rect 37036 8186 37092 8188
rect 37116 8186 37172 8188
rect 37196 8186 37252 8188
rect 36956 8134 37002 8186
rect 37002 8134 37012 8186
rect 37036 8134 37066 8186
rect 37066 8134 37078 8186
rect 37078 8134 37092 8186
rect 37116 8134 37130 8186
rect 37130 8134 37142 8186
rect 37142 8134 37172 8186
rect 37196 8134 37206 8186
rect 37206 8134 37252 8186
rect 36956 8132 37012 8134
rect 37036 8132 37092 8134
rect 37116 8132 37172 8134
rect 37196 8132 37252 8134
rect 41956 8186 42012 8188
rect 42036 8186 42092 8188
rect 42116 8186 42172 8188
rect 42196 8186 42252 8188
rect 41956 8134 42002 8186
rect 42002 8134 42012 8186
rect 42036 8134 42066 8186
rect 42066 8134 42078 8186
rect 42078 8134 42092 8186
rect 42116 8134 42130 8186
rect 42130 8134 42142 8186
rect 42142 8134 42172 8186
rect 42196 8134 42206 8186
rect 42206 8134 42252 8186
rect 41956 8132 42012 8134
rect 42036 8132 42092 8134
rect 42116 8132 42172 8134
rect 42196 8132 42252 8134
rect 46956 8186 47012 8188
rect 47036 8186 47092 8188
rect 47116 8186 47172 8188
rect 47196 8186 47252 8188
rect 46956 8134 47002 8186
rect 47002 8134 47012 8186
rect 47036 8134 47066 8186
rect 47066 8134 47078 8186
rect 47078 8134 47092 8186
rect 47116 8134 47130 8186
rect 47130 8134 47142 8186
rect 47142 8134 47172 8186
rect 47196 8134 47206 8186
rect 47206 8134 47252 8186
rect 46956 8132 47012 8134
rect 47036 8132 47092 8134
rect 47116 8132 47172 8134
rect 47196 8132 47252 8134
rect 51956 8186 52012 8188
rect 52036 8186 52092 8188
rect 52116 8186 52172 8188
rect 52196 8186 52252 8188
rect 51956 8134 52002 8186
rect 52002 8134 52012 8186
rect 52036 8134 52066 8186
rect 52066 8134 52078 8186
rect 52078 8134 52092 8186
rect 52116 8134 52130 8186
rect 52130 8134 52142 8186
rect 52142 8134 52172 8186
rect 52196 8134 52206 8186
rect 52206 8134 52252 8186
rect 51956 8132 52012 8134
rect 52036 8132 52092 8134
rect 52116 8132 52172 8134
rect 52196 8132 52252 8134
rect 56956 8186 57012 8188
rect 57036 8186 57092 8188
rect 57116 8186 57172 8188
rect 57196 8186 57252 8188
rect 56956 8134 57002 8186
rect 57002 8134 57012 8186
rect 57036 8134 57066 8186
rect 57066 8134 57078 8186
rect 57078 8134 57092 8186
rect 57116 8134 57130 8186
rect 57130 8134 57142 8186
rect 57142 8134 57172 8186
rect 57196 8134 57206 8186
rect 57206 8134 57252 8186
rect 56956 8132 57012 8134
rect 57036 8132 57092 8134
rect 57116 8132 57172 8134
rect 57196 8132 57252 8134
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 22616 7642 22672 7644
rect 22696 7642 22752 7644
rect 22776 7642 22832 7644
rect 22856 7642 22912 7644
rect 22616 7590 22662 7642
rect 22662 7590 22672 7642
rect 22696 7590 22726 7642
rect 22726 7590 22738 7642
rect 22738 7590 22752 7642
rect 22776 7590 22790 7642
rect 22790 7590 22802 7642
rect 22802 7590 22832 7642
rect 22856 7590 22866 7642
rect 22866 7590 22912 7642
rect 22616 7588 22672 7590
rect 22696 7588 22752 7590
rect 22776 7588 22832 7590
rect 22856 7588 22912 7590
rect 27616 7642 27672 7644
rect 27696 7642 27752 7644
rect 27776 7642 27832 7644
rect 27856 7642 27912 7644
rect 27616 7590 27662 7642
rect 27662 7590 27672 7642
rect 27696 7590 27726 7642
rect 27726 7590 27738 7642
rect 27738 7590 27752 7642
rect 27776 7590 27790 7642
rect 27790 7590 27802 7642
rect 27802 7590 27832 7642
rect 27856 7590 27866 7642
rect 27866 7590 27912 7642
rect 27616 7588 27672 7590
rect 27696 7588 27752 7590
rect 27776 7588 27832 7590
rect 27856 7588 27912 7590
rect 32616 7642 32672 7644
rect 32696 7642 32752 7644
rect 32776 7642 32832 7644
rect 32856 7642 32912 7644
rect 32616 7590 32662 7642
rect 32662 7590 32672 7642
rect 32696 7590 32726 7642
rect 32726 7590 32738 7642
rect 32738 7590 32752 7642
rect 32776 7590 32790 7642
rect 32790 7590 32802 7642
rect 32802 7590 32832 7642
rect 32856 7590 32866 7642
rect 32866 7590 32912 7642
rect 32616 7588 32672 7590
rect 32696 7588 32752 7590
rect 32776 7588 32832 7590
rect 32856 7588 32912 7590
rect 37616 7642 37672 7644
rect 37696 7642 37752 7644
rect 37776 7642 37832 7644
rect 37856 7642 37912 7644
rect 37616 7590 37662 7642
rect 37662 7590 37672 7642
rect 37696 7590 37726 7642
rect 37726 7590 37738 7642
rect 37738 7590 37752 7642
rect 37776 7590 37790 7642
rect 37790 7590 37802 7642
rect 37802 7590 37832 7642
rect 37856 7590 37866 7642
rect 37866 7590 37912 7642
rect 37616 7588 37672 7590
rect 37696 7588 37752 7590
rect 37776 7588 37832 7590
rect 37856 7588 37912 7590
rect 42616 7642 42672 7644
rect 42696 7642 42752 7644
rect 42776 7642 42832 7644
rect 42856 7642 42912 7644
rect 42616 7590 42662 7642
rect 42662 7590 42672 7642
rect 42696 7590 42726 7642
rect 42726 7590 42738 7642
rect 42738 7590 42752 7642
rect 42776 7590 42790 7642
rect 42790 7590 42802 7642
rect 42802 7590 42832 7642
rect 42856 7590 42866 7642
rect 42866 7590 42912 7642
rect 42616 7588 42672 7590
rect 42696 7588 42752 7590
rect 42776 7588 42832 7590
rect 42856 7588 42912 7590
rect 47616 7642 47672 7644
rect 47696 7642 47752 7644
rect 47776 7642 47832 7644
rect 47856 7642 47912 7644
rect 47616 7590 47662 7642
rect 47662 7590 47672 7642
rect 47696 7590 47726 7642
rect 47726 7590 47738 7642
rect 47738 7590 47752 7642
rect 47776 7590 47790 7642
rect 47790 7590 47802 7642
rect 47802 7590 47832 7642
rect 47856 7590 47866 7642
rect 47866 7590 47912 7642
rect 47616 7588 47672 7590
rect 47696 7588 47752 7590
rect 47776 7588 47832 7590
rect 47856 7588 47912 7590
rect 52616 7642 52672 7644
rect 52696 7642 52752 7644
rect 52776 7642 52832 7644
rect 52856 7642 52912 7644
rect 52616 7590 52662 7642
rect 52662 7590 52672 7642
rect 52696 7590 52726 7642
rect 52726 7590 52738 7642
rect 52738 7590 52752 7642
rect 52776 7590 52790 7642
rect 52790 7590 52802 7642
rect 52802 7590 52832 7642
rect 52856 7590 52866 7642
rect 52866 7590 52912 7642
rect 52616 7588 52672 7590
rect 52696 7588 52752 7590
rect 52776 7588 52832 7590
rect 52856 7588 52912 7590
rect 57616 7642 57672 7644
rect 57696 7642 57752 7644
rect 57776 7642 57832 7644
rect 57856 7642 57912 7644
rect 57616 7590 57662 7642
rect 57662 7590 57672 7642
rect 57696 7590 57726 7642
rect 57726 7590 57738 7642
rect 57738 7590 57752 7642
rect 57776 7590 57790 7642
rect 57790 7590 57802 7642
rect 57802 7590 57832 7642
rect 57856 7590 57866 7642
rect 57866 7590 57912 7642
rect 57616 7588 57672 7590
rect 57696 7588 57752 7590
rect 57776 7588 57832 7590
rect 57856 7588 57912 7590
rect 58530 7384 58586 7440
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 21956 7098 22012 7100
rect 22036 7098 22092 7100
rect 22116 7098 22172 7100
rect 22196 7098 22252 7100
rect 21956 7046 22002 7098
rect 22002 7046 22012 7098
rect 22036 7046 22066 7098
rect 22066 7046 22078 7098
rect 22078 7046 22092 7098
rect 22116 7046 22130 7098
rect 22130 7046 22142 7098
rect 22142 7046 22172 7098
rect 22196 7046 22206 7098
rect 22206 7046 22252 7098
rect 21956 7044 22012 7046
rect 22036 7044 22092 7046
rect 22116 7044 22172 7046
rect 22196 7044 22252 7046
rect 26956 7098 27012 7100
rect 27036 7098 27092 7100
rect 27116 7098 27172 7100
rect 27196 7098 27252 7100
rect 26956 7046 27002 7098
rect 27002 7046 27012 7098
rect 27036 7046 27066 7098
rect 27066 7046 27078 7098
rect 27078 7046 27092 7098
rect 27116 7046 27130 7098
rect 27130 7046 27142 7098
rect 27142 7046 27172 7098
rect 27196 7046 27206 7098
rect 27206 7046 27252 7098
rect 26956 7044 27012 7046
rect 27036 7044 27092 7046
rect 27116 7044 27172 7046
rect 27196 7044 27252 7046
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 36956 7098 37012 7100
rect 37036 7098 37092 7100
rect 37116 7098 37172 7100
rect 37196 7098 37252 7100
rect 36956 7046 37002 7098
rect 37002 7046 37012 7098
rect 37036 7046 37066 7098
rect 37066 7046 37078 7098
rect 37078 7046 37092 7098
rect 37116 7046 37130 7098
rect 37130 7046 37142 7098
rect 37142 7046 37172 7098
rect 37196 7046 37206 7098
rect 37206 7046 37252 7098
rect 36956 7044 37012 7046
rect 37036 7044 37092 7046
rect 37116 7044 37172 7046
rect 37196 7044 37252 7046
rect 41956 7098 42012 7100
rect 42036 7098 42092 7100
rect 42116 7098 42172 7100
rect 42196 7098 42252 7100
rect 41956 7046 42002 7098
rect 42002 7046 42012 7098
rect 42036 7046 42066 7098
rect 42066 7046 42078 7098
rect 42078 7046 42092 7098
rect 42116 7046 42130 7098
rect 42130 7046 42142 7098
rect 42142 7046 42172 7098
rect 42196 7046 42206 7098
rect 42206 7046 42252 7098
rect 41956 7044 42012 7046
rect 42036 7044 42092 7046
rect 42116 7044 42172 7046
rect 42196 7044 42252 7046
rect 46956 7098 47012 7100
rect 47036 7098 47092 7100
rect 47116 7098 47172 7100
rect 47196 7098 47252 7100
rect 46956 7046 47002 7098
rect 47002 7046 47012 7098
rect 47036 7046 47066 7098
rect 47066 7046 47078 7098
rect 47078 7046 47092 7098
rect 47116 7046 47130 7098
rect 47130 7046 47142 7098
rect 47142 7046 47172 7098
rect 47196 7046 47206 7098
rect 47206 7046 47252 7098
rect 46956 7044 47012 7046
rect 47036 7044 47092 7046
rect 47116 7044 47172 7046
rect 47196 7044 47252 7046
rect 51956 7098 52012 7100
rect 52036 7098 52092 7100
rect 52116 7098 52172 7100
rect 52196 7098 52252 7100
rect 51956 7046 52002 7098
rect 52002 7046 52012 7098
rect 52036 7046 52066 7098
rect 52066 7046 52078 7098
rect 52078 7046 52092 7098
rect 52116 7046 52130 7098
rect 52130 7046 52142 7098
rect 52142 7046 52172 7098
rect 52196 7046 52206 7098
rect 52206 7046 52252 7098
rect 51956 7044 52012 7046
rect 52036 7044 52092 7046
rect 52116 7044 52172 7046
rect 52196 7044 52252 7046
rect 56956 7098 57012 7100
rect 57036 7098 57092 7100
rect 57116 7098 57172 7100
rect 57196 7098 57252 7100
rect 56956 7046 57002 7098
rect 57002 7046 57012 7098
rect 57036 7046 57066 7098
rect 57066 7046 57078 7098
rect 57078 7046 57092 7098
rect 57116 7046 57130 7098
rect 57130 7046 57142 7098
rect 57142 7046 57172 7098
rect 57196 7046 57206 7098
rect 57206 7046 57252 7098
rect 56956 7044 57012 7046
rect 57036 7044 57092 7046
rect 57116 7044 57172 7046
rect 57196 7044 57252 7046
rect 58530 6568 58586 6624
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 22616 6554 22672 6556
rect 22696 6554 22752 6556
rect 22776 6554 22832 6556
rect 22856 6554 22912 6556
rect 22616 6502 22662 6554
rect 22662 6502 22672 6554
rect 22696 6502 22726 6554
rect 22726 6502 22738 6554
rect 22738 6502 22752 6554
rect 22776 6502 22790 6554
rect 22790 6502 22802 6554
rect 22802 6502 22832 6554
rect 22856 6502 22866 6554
rect 22866 6502 22912 6554
rect 22616 6500 22672 6502
rect 22696 6500 22752 6502
rect 22776 6500 22832 6502
rect 22856 6500 22912 6502
rect 27616 6554 27672 6556
rect 27696 6554 27752 6556
rect 27776 6554 27832 6556
rect 27856 6554 27912 6556
rect 27616 6502 27662 6554
rect 27662 6502 27672 6554
rect 27696 6502 27726 6554
rect 27726 6502 27738 6554
rect 27738 6502 27752 6554
rect 27776 6502 27790 6554
rect 27790 6502 27802 6554
rect 27802 6502 27832 6554
rect 27856 6502 27866 6554
rect 27866 6502 27912 6554
rect 27616 6500 27672 6502
rect 27696 6500 27752 6502
rect 27776 6500 27832 6502
rect 27856 6500 27912 6502
rect 32616 6554 32672 6556
rect 32696 6554 32752 6556
rect 32776 6554 32832 6556
rect 32856 6554 32912 6556
rect 32616 6502 32662 6554
rect 32662 6502 32672 6554
rect 32696 6502 32726 6554
rect 32726 6502 32738 6554
rect 32738 6502 32752 6554
rect 32776 6502 32790 6554
rect 32790 6502 32802 6554
rect 32802 6502 32832 6554
rect 32856 6502 32866 6554
rect 32866 6502 32912 6554
rect 32616 6500 32672 6502
rect 32696 6500 32752 6502
rect 32776 6500 32832 6502
rect 32856 6500 32912 6502
rect 37616 6554 37672 6556
rect 37696 6554 37752 6556
rect 37776 6554 37832 6556
rect 37856 6554 37912 6556
rect 37616 6502 37662 6554
rect 37662 6502 37672 6554
rect 37696 6502 37726 6554
rect 37726 6502 37738 6554
rect 37738 6502 37752 6554
rect 37776 6502 37790 6554
rect 37790 6502 37802 6554
rect 37802 6502 37832 6554
rect 37856 6502 37866 6554
rect 37866 6502 37912 6554
rect 37616 6500 37672 6502
rect 37696 6500 37752 6502
rect 37776 6500 37832 6502
rect 37856 6500 37912 6502
rect 42616 6554 42672 6556
rect 42696 6554 42752 6556
rect 42776 6554 42832 6556
rect 42856 6554 42912 6556
rect 42616 6502 42662 6554
rect 42662 6502 42672 6554
rect 42696 6502 42726 6554
rect 42726 6502 42738 6554
rect 42738 6502 42752 6554
rect 42776 6502 42790 6554
rect 42790 6502 42802 6554
rect 42802 6502 42832 6554
rect 42856 6502 42866 6554
rect 42866 6502 42912 6554
rect 42616 6500 42672 6502
rect 42696 6500 42752 6502
rect 42776 6500 42832 6502
rect 42856 6500 42912 6502
rect 47616 6554 47672 6556
rect 47696 6554 47752 6556
rect 47776 6554 47832 6556
rect 47856 6554 47912 6556
rect 47616 6502 47662 6554
rect 47662 6502 47672 6554
rect 47696 6502 47726 6554
rect 47726 6502 47738 6554
rect 47738 6502 47752 6554
rect 47776 6502 47790 6554
rect 47790 6502 47802 6554
rect 47802 6502 47832 6554
rect 47856 6502 47866 6554
rect 47866 6502 47912 6554
rect 47616 6500 47672 6502
rect 47696 6500 47752 6502
rect 47776 6500 47832 6502
rect 47856 6500 47912 6502
rect 52616 6554 52672 6556
rect 52696 6554 52752 6556
rect 52776 6554 52832 6556
rect 52856 6554 52912 6556
rect 52616 6502 52662 6554
rect 52662 6502 52672 6554
rect 52696 6502 52726 6554
rect 52726 6502 52738 6554
rect 52738 6502 52752 6554
rect 52776 6502 52790 6554
rect 52790 6502 52802 6554
rect 52802 6502 52832 6554
rect 52856 6502 52866 6554
rect 52866 6502 52912 6554
rect 52616 6500 52672 6502
rect 52696 6500 52752 6502
rect 52776 6500 52832 6502
rect 52856 6500 52912 6502
rect 57616 6554 57672 6556
rect 57696 6554 57752 6556
rect 57776 6554 57832 6556
rect 57856 6554 57912 6556
rect 57616 6502 57662 6554
rect 57662 6502 57672 6554
rect 57696 6502 57726 6554
rect 57726 6502 57738 6554
rect 57738 6502 57752 6554
rect 57776 6502 57790 6554
rect 57790 6502 57802 6554
rect 57802 6502 57832 6554
rect 57856 6502 57866 6554
rect 57866 6502 57912 6554
rect 57616 6500 57672 6502
rect 57696 6500 57752 6502
rect 57776 6500 57832 6502
rect 57856 6500 57912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 21956 6010 22012 6012
rect 22036 6010 22092 6012
rect 22116 6010 22172 6012
rect 22196 6010 22252 6012
rect 21956 5958 22002 6010
rect 22002 5958 22012 6010
rect 22036 5958 22066 6010
rect 22066 5958 22078 6010
rect 22078 5958 22092 6010
rect 22116 5958 22130 6010
rect 22130 5958 22142 6010
rect 22142 5958 22172 6010
rect 22196 5958 22206 6010
rect 22206 5958 22252 6010
rect 21956 5956 22012 5958
rect 22036 5956 22092 5958
rect 22116 5956 22172 5958
rect 22196 5956 22252 5958
rect 26956 6010 27012 6012
rect 27036 6010 27092 6012
rect 27116 6010 27172 6012
rect 27196 6010 27252 6012
rect 26956 5958 27002 6010
rect 27002 5958 27012 6010
rect 27036 5958 27066 6010
rect 27066 5958 27078 6010
rect 27078 5958 27092 6010
rect 27116 5958 27130 6010
rect 27130 5958 27142 6010
rect 27142 5958 27172 6010
rect 27196 5958 27206 6010
rect 27206 5958 27252 6010
rect 26956 5956 27012 5958
rect 27036 5956 27092 5958
rect 27116 5956 27172 5958
rect 27196 5956 27252 5958
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 36956 6010 37012 6012
rect 37036 6010 37092 6012
rect 37116 6010 37172 6012
rect 37196 6010 37252 6012
rect 36956 5958 37002 6010
rect 37002 5958 37012 6010
rect 37036 5958 37066 6010
rect 37066 5958 37078 6010
rect 37078 5958 37092 6010
rect 37116 5958 37130 6010
rect 37130 5958 37142 6010
rect 37142 5958 37172 6010
rect 37196 5958 37206 6010
rect 37206 5958 37252 6010
rect 36956 5956 37012 5958
rect 37036 5956 37092 5958
rect 37116 5956 37172 5958
rect 37196 5956 37252 5958
rect 41956 6010 42012 6012
rect 42036 6010 42092 6012
rect 42116 6010 42172 6012
rect 42196 6010 42252 6012
rect 41956 5958 42002 6010
rect 42002 5958 42012 6010
rect 42036 5958 42066 6010
rect 42066 5958 42078 6010
rect 42078 5958 42092 6010
rect 42116 5958 42130 6010
rect 42130 5958 42142 6010
rect 42142 5958 42172 6010
rect 42196 5958 42206 6010
rect 42206 5958 42252 6010
rect 41956 5956 42012 5958
rect 42036 5956 42092 5958
rect 42116 5956 42172 5958
rect 42196 5956 42252 5958
rect 46956 6010 47012 6012
rect 47036 6010 47092 6012
rect 47116 6010 47172 6012
rect 47196 6010 47252 6012
rect 46956 5958 47002 6010
rect 47002 5958 47012 6010
rect 47036 5958 47066 6010
rect 47066 5958 47078 6010
rect 47078 5958 47092 6010
rect 47116 5958 47130 6010
rect 47130 5958 47142 6010
rect 47142 5958 47172 6010
rect 47196 5958 47206 6010
rect 47206 5958 47252 6010
rect 46956 5956 47012 5958
rect 47036 5956 47092 5958
rect 47116 5956 47172 5958
rect 47196 5956 47252 5958
rect 51956 6010 52012 6012
rect 52036 6010 52092 6012
rect 52116 6010 52172 6012
rect 52196 6010 52252 6012
rect 51956 5958 52002 6010
rect 52002 5958 52012 6010
rect 52036 5958 52066 6010
rect 52066 5958 52078 6010
rect 52078 5958 52092 6010
rect 52116 5958 52130 6010
rect 52130 5958 52142 6010
rect 52142 5958 52172 6010
rect 52196 5958 52206 6010
rect 52206 5958 52252 6010
rect 51956 5956 52012 5958
rect 52036 5956 52092 5958
rect 52116 5956 52172 5958
rect 52196 5956 52252 5958
rect 56956 6010 57012 6012
rect 57036 6010 57092 6012
rect 57116 6010 57172 6012
rect 57196 6010 57252 6012
rect 56956 5958 57002 6010
rect 57002 5958 57012 6010
rect 57036 5958 57066 6010
rect 57066 5958 57078 6010
rect 57078 5958 57092 6010
rect 57116 5958 57130 6010
rect 57130 5958 57142 6010
rect 57142 5958 57172 6010
rect 57196 5958 57206 6010
rect 57206 5958 57252 6010
rect 56956 5956 57012 5958
rect 57036 5956 57092 5958
rect 57116 5956 57172 5958
rect 57196 5956 57252 5958
rect 58530 5752 58586 5808
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 22616 5466 22672 5468
rect 22696 5466 22752 5468
rect 22776 5466 22832 5468
rect 22856 5466 22912 5468
rect 22616 5414 22662 5466
rect 22662 5414 22672 5466
rect 22696 5414 22726 5466
rect 22726 5414 22738 5466
rect 22738 5414 22752 5466
rect 22776 5414 22790 5466
rect 22790 5414 22802 5466
rect 22802 5414 22832 5466
rect 22856 5414 22866 5466
rect 22866 5414 22912 5466
rect 22616 5412 22672 5414
rect 22696 5412 22752 5414
rect 22776 5412 22832 5414
rect 22856 5412 22912 5414
rect 27616 5466 27672 5468
rect 27696 5466 27752 5468
rect 27776 5466 27832 5468
rect 27856 5466 27912 5468
rect 27616 5414 27662 5466
rect 27662 5414 27672 5466
rect 27696 5414 27726 5466
rect 27726 5414 27738 5466
rect 27738 5414 27752 5466
rect 27776 5414 27790 5466
rect 27790 5414 27802 5466
rect 27802 5414 27832 5466
rect 27856 5414 27866 5466
rect 27866 5414 27912 5466
rect 27616 5412 27672 5414
rect 27696 5412 27752 5414
rect 27776 5412 27832 5414
rect 27856 5412 27912 5414
rect 32616 5466 32672 5468
rect 32696 5466 32752 5468
rect 32776 5466 32832 5468
rect 32856 5466 32912 5468
rect 32616 5414 32662 5466
rect 32662 5414 32672 5466
rect 32696 5414 32726 5466
rect 32726 5414 32738 5466
rect 32738 5414 32752 5466
rect 32776 5414 32790 5466
rect 32790 5414 32802 5466
rect 32802 5414 32832 5466
rect 32856 5414 32866 5466
rect 32866 5414 32912 5466
rect 32616 5412 32672 5414
rect 32696 5412 32752 5414
rect 32776 5412 32832 5414
rect 32856 5412 32912 5414
rect 37616 5466 37672 5468
rect 37696 5466 37752 5468
rect 37776 5466 37832 5468
rect 37856 5466 37912 5468
rect 37616 5414 37662 5466
rect 37662 5414 37672 5466
rect 37696 5414 37726 5466
rect 37726 5414 37738 5466
rect 37738 5414 37752 5466
rect 37776 5414 37790 5466
rect 37790 5414 37802 5466
rect 37802 5414 37832 5466
rect 37856 5414 37866 5466
rect 37866 5414 37912 5466
rect 37616 5412 37672 5414
rect 37696 5412 37752 5414
rect 37776 5412 37832 5414
rect 37856 5412 37912 5414
rect 42616 5466 42672 5468
rect 42696 5466 42752 5468
rect 42776 5466 42832 5468
rect 42856 5466 42912 5468
rect 42616 5414 42662 5466
rect 42662 5414 42672 5466
rect 42696 5414 42726 5466
rect 42726 5414 42738 5466
rect 42738 5414 42752 5466
rect 42776 5414 42790 5466
rect 42790 5414 42802 5466
rect 42802 5414 42832 5466
rect 42856 5414 42866 5466
rect 42866 5414 42912 5466
rect 42616 5412 42672 5414
rect 42696 5412 42752 5414
rect 42776 5412 42832 5414
rect 42856 5412 42912 5414
rect 47616 5466 47672 5468
rect 47696 5466 47752 5468
rect 47776 5466 47832 5468
rect 47856 5466 47912 5468
rect 47616 5414 47662 5466
rect 47662 5414 47672 5466
rect 47696 5414 47726 5466
rect 47726 5414 47738 5466
rect 47738 5414 47752 5466
rect 47776 5414 47790 5466
rect 47790 5414 47802 5466
rect 47802 5414 47832 5466
rect 47856 5414 47866 5466
rect 47866 5414 47912 5466
rect 47616 5412 47672 5414
rect 47696 5412 47752 5414
rect 47776 5412 47832 5414
rect 47856 5412 47912 5414
rect 52616 5466 52672 5468
rect 52696 5466 52752 5468
rect 52776 5466 52832 5468
rect 52856 5466 52912 5468
rect 52616 5414 52662 5466
rect 52662 5414 52672 5466
rect 52696 5414 52726 5466
rect 52726 5414 52738 5466
rect 52738 5414 52752 5466
rect 52776 5414 52790 5466
rect 52790 5414 52802 5466
rect 52802 5414 52832 5466
rect 52856 5414 52866 5466
rect 52866 5414 52912 5466
rect 52616 5412 52672 5414
rect 52696 5412 52752 5414
rect 52776 5412 52832 5414
rect 52856 5412 52912 5414
rect 57616 5466 57672 5468
rect 57696 5466 57752 5468
rect 57776 5466 57832 5468
rect 57856 5466 57912 5468
rect 57616 5414 57662 5466
rect 57662 5414 57672 5466
rect 57696 5414 57726 5466
rect 57726 5414 57738 5466
rect 57738 5414 57752 5466
rect 57776 5414 57790 5466
rect 57790 5414 57802 5466
rect 57802 5414 57832 5466
rect 57856 5414 57866 5466
rect 57866 5414 57912 5466
rect 57616 5412 57672 5414
rect 57696 5412 57752 5414
rect 57776 5412 57832 5414
rect 57856 5412 57912 5414
rect 58530 4972 58532 4992
rect 58532 4972 58584 4992
rect 58584 4972 58586 4992
rect 58530 4936 58586 4972
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 21956 4922 22012 4924
rect 22036 4922 22092 4924
rect 22116 4922 22172 4924
rect 22196 4922 22252 4924
rect 21956 4870 22002 4922
rect 22002 4870 22012 4922
rect 22036 4870 22066 4922
rect 22066 4870 22078 4922
rect 22078 4870 22092 4922
rect 22116 4870 22130 4922
rect 22130 4870 22142 4922
rect 22142 4870 22172 4922
rect 22196 4870 22206 4922
rect 22206 4870 22252 4922
rect 21956 4868 22012 4870
rect 22036 4868 22092 4870
rect 22116 4868 22172 4870
rect 22196 4868 22252 4870
rect 26956 4922 27012 4924
rect 27036 4922 27092 4924
rect 27116 4922 27172 4924
rect 27196 4922 27252 4924
rect 26956 4870 27002 4922
rect 27002 4870 27012 4922
rect 27036 4870 27066 4922
rect 27066 4870 27078 4922
rect 27078 4870 27092 4922
rect 27116 4870 27130 4922
rect 27130 4870 27142 4922
rect 27142 4870 27172 4922
rect 27196 4870 27206 4922
rect 27206 4870 27252 4922
rect 26956 4868 27012 4870
rect 27036 4868 27092 4870
rect 27116 4868 27172 4870
rect 27196 4868 27252 4870
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 36956 4922 37012 4924
rect 37036 4922 37092 4924
rect 37116 4922 37172 4924
rect 37196 4922 37252 4924
rect 36956 4870 37002 4922
rect 37002 4870 37012 4922
rect 37036 4870 37066 4922
rect 37066 4870 37078 4922
rect 37078 4870 37092 4922
rect 37116 4870 37130 4922
rect 37130 4870 37142 4922
rect 37142 4870 37172 4922
rect 37196 4870 37206 4922
rect 37206 4870 37252 4922
rect 36956 4868 37012 4870
rect 37036 4868 37092 4870
rect 37116 4868 37172 4870
rect 37196 4868 37252 4870
rect 41956 4922 42012 4924
rect 42036 4922 42092 4924
rect 42116 4922 42172 4924
rect 42196 4922 42252 4924
rect 41956 4870 42002 4922
rect 42002 4870 42012 4922
rect 42036 4870 42066 4922
rect 42066 4870 42078 4922
rect 42078 4870 42092 4922
rect 42116 4870 42130 4922
rect 42130 4870 42142 4922
rect 42142 4870 42172 4922
rect 42196 4870 42206 4922
rect 42206 4870 42252 4922
rect 41956 4868 42012 4870
rect 42036 4868 42092 4870
rect 42116 4868 42172 4870
rect 42196 4868 42252 4870
rect 46956 4922 47012 4924
rect 47036 4922 47092 4924
rect 47116 4922 47172 4924
rect 47196 4922 47252 4924
rect 46956 4870 47002 4922
rect 47002 4870 47012 4922
rect 47036 4870 47066 4922
rect 47066 4870 47078 4922
rect 47078 4870 47092 4922
rect 47116 4870 47130 4922
rect 47130 4870 47142 4922
rect 47142 4870 47172 4922
rect 47196 4870 47206 4922
rect 47206 4870 47252 4922
rect 46956 4868 47012 4870
rect 47036 4868 47092 4870
rect 47116 4868 47172 4870
rect 47196 4868 47252 4870
rect 51956 4922 52012 4924
rect 52036 4922 52092 4924
rect 52116 4922 52172 4924
rect 52196 4922 52252 4924
rect 51956 4870 52002 4922
rect 52002 4870 52012 4922
rect 52036 4870 52066 4922
rect 52066 4870 52078 4922
rect 52078 4870 52092 4922
rect 52116 4870 52130 4922
rect 52130 4870 52142 4922
rect 52142 4870 52172 4922
rect 52196 4870 52206 4922
rect 52206 4870 52252 4922
rect 51956 4868 52012 4870
rect 52036 4868 52092 4870
rect 52116 4868 52172 4870
rect 52196 4868 52252 4870
rect 56956 4922 57012 4924
rect 57036 4922 57092 4924
rect 57116 4922 57172 4924
rect 57196 4922 57252 4924
rect 56956 4870 57002 4922
rect 57002 4870 57012 4922
rect 57036 4870 57066 4922
rect 57066 4870 57078 4922
rect 57078 4870 57092 4922
rect 57116 4870 57130 4922
rect 57130 4870 57142 4922
rect 57142 4870 57172 4922
rect 57196 4870 57206 4922
rect 57206 4870 57252 4922
rect 56956 4868 57012 4870
rect 57036 4868 57092 4870
rect 57116 4868 57172 4870
rect 57196 4868 57252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 22616 4378 22672 4380
rect 22696 4378 22752 4380
rect 22776 4378 22832 4380
rect 22856 4378 22912 4380
rect 22616 4326 22662 4378
rect 22662 4326 22672 4378
rect 22696 4326 22726 4378
rect 22726 4326 22738 4378
rect 22738 4326 22752 4378
rect 22776 4326 22790 4378
rect 22790 4326 22802 4378
rect 22802 4326 22832 4378
rect 22856 4326 22866 4378
rect 22866 4326 22912 4378
rect 22616 4324 22672 4326
rect 22696 4324 22752 4326
rect 22776 4324 22832 4326
rect 22856 4324 22912 4326
rect 27616 4378 27672 4380
rect 27696 4378 27752 4380
rect 27776 4378 27832 4380
rect 27856 4378 27912 4380
rect 27616 4326 27662 4378
rect 27662 4326 27672 4378
rect 27696 4326 27726 4378
rect 27726 4326 27738 4378
rect 27738 4326 27752 4378
rect 27776 4326 27790 4378
rect 27790 4326 27802 4378
rect 27802 4326 27832 4378
rect 27856 4326 27866 4378
rect 27866 4326 27912 4378
rect 27616 4324 27672 4326
rect 27696 4324 27752 4326
rect 27776 4324 27832 4326
rect 27856 4324 27912 4326
rect 32616 4378 32672 4380
rect 32696 4378 32752 4380
rect 32776 4378 32832 4380
rect 32856 4378 32912 4380
rect 32616 4326 32662 4378
rect 32662 4326 32672 4378
rect 32696 4326 32726 4378
rect 32726 4326 32738 4378
rect 32738 4326 32752 4378
rect 32776 4326 32790 4378
rect 32790 4326 32802 4378
rect 32802 4326 32832 4378
rect 32856 4326 32866 4378
rect 32866 4326 32912 4378
rect 32616 4324 32672 4326
rect 32696 4324 32752 4326
rect 32776 4324 32832 4326
rect 32856 4324 32912 4326
rect 37616 4378 37672 4380
rect 37696 4378 37752 4380
rect 37776 4378 37832 4380
rect 37856 4378 37912 4380
rect 37616 4326 37662 4378
rect 37662 4326 37672 4378
rect 37696 4326 37726 4378
rect 37726 4326 37738 4378
rect 37738 4326 37752 4378
rect 37776 4326 37790 4378
rect 37790 4326 37802 4378
rect 37802 4326 37832 4378
rect 37856 4326 37866 4378
rect 37866 4326 37912 4378
rect 37616 4324 37672 4326
rect 37696 4324 37752 4326
rect 37776 4324 37832 4326
rect 37856 4324 37912 4326
rect 42616 4378 42672 4380
rect 42696 4378 42752 4380
rect 42776 4378 42832 4380
rect 42856 4378 42912 4380
rect 42616 4326 42662 4378
rect 42662 4326 42672 4378
rect 42696 4326 42726 4378
rect 42726 4326 42738 4378
rect 42738 4326 42752 4378
rect 42776 4326 42790 4378
rect 42790 4326 42802 4378
rect 42802 4326 42832 4378
rect 42856 4326 42866 4378
rect 42866 4326 42912 4378
rect 42616 4324 42672 4326
rect 42696 4324 42752 4326
rect 42776 4324 42832 4326
rect 42856 4324 42912 4326
rect 47616 4378 47672 4380
rect 47696 4378 47752 4380
rect 47776 4378 47832 4380
rect 47856 4378 47912 4380
rect 47616 4326 47662 4378
rect 47662 4326 47672 4378
rect 47696 4326 47726 4378
rect 47726 4326 47738 4378
rect 47738 4326 47752 4378
rect 47776 4326 47790 4378
rect 47790 4326 47802 4378
rect 47802 4326 47832 4378
rect 47856 4326 47866 4378
rect 47866 4326 47912 4378
rect 47616 4324 47672 4326
rect 47696 4324 47752 4326
rect 47776 4324 47832 4326
rect 47856 4324 47912 4326
rect 52616 4378 52672 4380
rect 52696 4378 52752 4380
rect 52776 4378 52832 4380
rect 52856 4378 52912 4380
rect 52616 4326 52662 4378
rect 52662 4326 52672 4378
rect 52696 4326 52726 4378
rect 52726 4326 52738 4378
rect 52738 4326 52752 4378
rect 52776 4326 52790 4378
rect 52790 4326 52802 4378
rect 52802 4326 52832 4378
rect 52856 4326 52866 4378
rect 52866 4326 52912 4378
rect 52616 4324 52672 4326
rect 52696 4324 52752 4326
rect 52776 4324 52832 4326
rect 52856 4324 52912 4326
rect 57616 4378 57672 4380
rect 57696 4378 57752 4380
rect 57776 4378 57832 4380
rect 57856 4378 57912 4380
rect 57616 4326 57662 4378
rect 57662 4326 57672 4378
rect 57696 4326 57726 4378
rect 57726 4326 57738 4378
rect 57738 4326 57752 4378
rect 57776 4326 57790 4378
rect 57790 4326 57802 4378
rect 57802 4326 57832 4378
rect 57856 4326 57866 4378
rect 57866 4326 57912 4378
rect 57616 4324 57672 4326
rect 57696 4324 57752 4326
rect 57776 4324 57832 4326
rect 57856 4324 57912 4326
rect 58530 4120 58586 4176
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 21956 3834 22012 3836
rect 22036 3834 22092 3836
rect 22116 3834 22172 3836
rect 22196 3834 22252 3836
rect 21956 3782 22002 3834
rect 22002 3782 22012 3834
rect 22036 3782 22066 3834
rect 22066 3782 22078 3834
rect 22078 3782 22092 3834
rect 22116 3782 22130 3834
rect 22130 3782 22142 3834
rect 22142 3782 22172 3834
rect 22196 3782 22206 3834
rect 22206 3782 22252 3834
rect 21956 3780 22012 3782
rect 22036 3780 22092 3782
rect 22116 3780 22172 3782
rect 22196 3780 22252 3782
rect 26956 3834 27012 3836
rect 27036 3834 27092 3836
rect 27116 3834 27172 3836
rect 27196 3834 27252 3836
rect 26956 3782 27002 3834
rect 27002 3782 27012 3834
rect 27036 3782 27066 3834
rect 27066 3782 27078 3834
rect 27078 3782 27092 3834
rect 27116 3782 27130 3834
rect 27130 3782 27142 3834
rect 27142 3782 27172 3834
rect 27196 3782 27206 3834
rect 27206 3782 27252 3834
rect 26956 3780 27012 3782
rect 27036 3780 27092 3782
rect 27116 3780 27172 3782
rect 27196 3780 27252 3782
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 36956 3834 37012 3836
rect 37036 3834 37092 3836
rect 37116 3834 37172 3836
rect 37196 3834 37252 3836
rect 36956 3782 37002 3834
rect 37002 3782 37012 3834
rect 37036 3782 37066 3834
rect 37066 3782 37078 3834
rect 37078 3782 37092 3834
rect 37116 3782 37130 3834
rect 37130 3782 37142 3834
rect 37142 3782 37172 3834
rect 37196 3782 37206 3834
rect 37206 3782 37252 3834
rect 36956 3780 37012 3782
rect 37036 3780 37092 3782
rect 37116 3780 37172 3782
rect 37196 3780 37252 3782
rect 41956 3834 42012 3836
rect 42036 3834 42092 3836
rect 42116 3834 42172 3836
rect 42196 3834 42252 3836
rect 41956 3782 42002 3834
rect 42002 3782 42012 3834
rect 42036 3782 42066 3834
rect 42066 3782 42078 3834
rect 42078 3782 42092 3834
rect 42116 3782 42130 3834
rect 42130 3782 42142 3834
rect 42142 3782 42172 3834
rect 42196 3782 42206 3834
rect 42206 3782 42252 3834
rect 41956 3780 42012 3782
rect 42036 3780 42092 3782
rect 42116 3780 42172 3782
rect 42196 3780 42252 3782
rect 46956 3834 47012 3836
rect 47036 3834 47092 3836
rect 47116 3834 47172 3836
rect 47196 3834 47252 3836
rect 46956 3782 47002 3834
rect 47002 3782 47012 3834
rect 47036 3782 47066 3834
rect 47066 3782 47078 3834
rect 47078 3782 47092 3834
rect 47116 3782 47130 3834
rect 47130 3782 47142 3834
rect 47142 3782 47172 3834
rect 47196 3782 47206 3834
rect 47206 3782 47252 3834
rect 46956 3780 47012 3782
rect 47036 3780 47092 3782
rect 47116 3780 47172 3782
rect 47196 3780 47252 3782
rect 51956 3834 52012 3836
rect 52036 3834 52092 3836
rect 52116 3834 52172 3836
rect 52196 3834 52252 3836
rect 51956 3782 52002 3834
rect 52002 3782 52012 3834
rect 52036 3782 52066 3834
rect 52066 3782 52078 3834
rect 52078 3782 52092 3834
rect 52116 3782 52130 3834
rect 52130 3782 52142 3834
rect 52142 3782 52172 3834
rect 52196 3782 52206 3834
rect 52206 3782 52252 3834
rect 51956 3780 52012 3782
rect 52036 3780 52092 3782
rect 52116 3780 52172 3782
rect 52196 3780 52252 3782
rect 56956 3834 57012 3836
rect 57036 3834 57092 3836
rect 57116 3834 57172 3836
rect 57196 3834 57252 3836
rect 56956 3782 57002 3834
rect 57002 3782 57012 3834
rect 57036 3782 57066 3834
rect 57066 3782 57078 3834
rect 57078 3782 57092 3834
rect 57116 3782 57130 3834
rect 57130 3782 57142 3834
rect 57142 3782 57172 3834
rect 57196 3782 57206 3834
rect 57206 3782 57252 3834
rect 56956 3780 57012 3782
rect 57036 3780 57092 3782
rect 57116 3780 57172 3782
rect 57196 3780 57252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 22616 3290 22672 3292
rect 22696 3290 22752 3292
rect 22776 3290 22832 3292
rect 22856 3290 22912 3292
rect 22616 3238 22662 3290
rect 22662 3238 22672 3290
rect 22696 3238 22726 3290
rect 22726 3238 22738 3290
rect 22738 3238 22752 3290
rect 22776 3238 22790 3290
rect 22790 3238 22802 3290
rect 22802 3238 22832 3290
rect 22856 3238 22866 3290
rect 22866 3238 22912 3290
rect 22616 3236 22672 3238
rect 22696 3236 22752 3238
rect 22776 3236 22832 3238
rect 22856 3236 22912 3238
rect 27616 3290 27672 3292
rect 27696 3290 27752 3292
rect 27776 3290 27832 3292
rect 27856 3290 27912 3292
rect 27616 3238 27662 3290
rect 27662 3238 27672 3290
rect 27696 3238 27726 3290
rect 27726 3238 27738 3290
rect 27738 3238 27752 3290
rect 27776 3238 27790 3290
rect 27790 3238 27802 3290
rect 27802 3238 27832 3290
rect 27856 3238 27866 3290
rect 27866 3238 27912 3290
rect 27616 3236 27672 3238
rect 27696 3236 27752 3238
rect 27776 3236 27832 3238
rect 27856 3236 27912 3238
rect 32616 3290 32672 3292
rect 32696 3290 32752 3292
rect 32776 3290 32832 3292
rect 32856 3290 32912 3292
rect 32616 3238 32662 3290
rect 32662 3238 32672 3290
rect 32696 3238 32726 3290
rect 32726 3238 32738 3290
rect 32738 3238 32752 3290
rect 32776 3238 32790 3290
rect 32790 3238 32802 3290
rect 32802 3238 32832 3290
rect 32856 3238 32866 3290
rect 32866 3238 32912 3290
rect 32616 3236 32672 3238
rect 32696 3236 32752 3238
rect 32776 3236 32832 3238
rect 32856 3236 32912 3238
rect 37616 3290 37672 3292
rect 37696 3290 37752 3292
rect 37776 3290 37832 3292
rect 37856 3290 37912 3292
rect 37616 3238 37662 3290
rect 37662 3238 37672 3290
rect 37696 3238 37726 3290
rect 37726 3238 37738 3290
rect 37738 3238 37752 3290
rect 37776 3238 37790 3290
rect 37790 3238 37802 3290
rect 37802 3238 37832 3290
rect 37856 3238 37866 3290
rect 37866 3238 37912 3290
rect 37616 3236 37672 3238
rect 37696 3236 37752 3238
rect 37776 3236 37832 3238
rect 37856 3236 37912 3238
rect 42616 3290 42672 3292
rect 42696 3290 42752 3292
rect 42776 3290 42832 3292
rect 42856 3290 42912 3292
rect 42616 3238 42662 3290
rect 42662 3238 42672 3290
rect 42696 3238 42726 3290
rect 42726 3238 42738 3290
rect 42738 3238 42752 3290
rect 42776 3238 42790 3290
rect 42790 3238 42802 3290
rect 42802 3238 42832 3290
rect 42856 3238 42866 3290
rect 42866 3238 42912 3290
rect 42616 3236 42672 3238
rect 42696 3236 42752 3238
rect 42776 3236 42832 3238
rect 42856 3236 42912 3238
rect 47616 3290 47672 3292
rect 47696 3290 47752 3292
rect 47776 3290 47832 3292
rect 47856 3290 47912 3292
rect 47616 3238 47662 3290
rect 47662 3238 47672 3290
rect 47696 3238 47726 3290
rect 47726 3238 47738 3290
rect 47738 3238 47752 3290
rect 47776 3238 47790 3290
rect 47790 3238 47802 3290
rect 47802 3238 47832 3290
rect 47856 3238 47866 3290
rect 47866 3238 47912 3290
rect 47616 3236 47672 3238
rect 47696 3236 47752 3238
rect 47776 3236 47832 3238
rect 47856 3236 47912 3238
rect 52616 3290 52672 3292
rect 52696 3290 52752 3292
rect 52776 3290 52832 3292
rect 52856 3290 52912 3292
rect 52616 3238 52662 3290
rect 52662 3238 52672 3290
rect 52696 3238 52726 3290
rect 52726 3238 52738 3290
rect 52738 3238 52752 3290
rect 52776 3238 52790 3290
rect 52790 3238 52802 3290
rect 52802 3238 52832 3290
rect 52856 3238 52866 3290
rect 52866 3238 52912 3290
rect 52616 3236 52672 3238
rect 52696 3236 52752 3238
rect 52776 3236 52832 3238
rect 52856 3236 52912 3238
rect 57616 3290 57672 3292
rect 57696 3290 57752 3292
rect 57776 3290 57832 3292
rect 57856 3290 57912 3292
rect 57616 3238 57662 3290
rect 57662 3238 57672 3290
rect 57696 3238 57726 3290
rect 57726 3238 57738 3290
rect 57738 3238 57752 3290
rect 57776 3238 57790 3290
rect 57790 3238 57802 3290
rect 57802 3238 57832 3290
rect 57856 3238 57866 3290
rect 57866 3238 57912 3290
rect 57616 3236 57672 3238
rect 57696 3236 57752 3238
rect 57776 3236 57832 3238
rect 57856 3236 57912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 21956 2746 22012 2748
rect 22036 2746 22092 2748
rect 22116 2746 22172 2748
rect 22196 2746 22252 2748
rect 21956 2694 22002 2746
rect 22002 2694 22012 2746
rect 22036 2694 22066 2746
rect 22066 2694 22078 2746
rect 22078 2694 22092 2746
rect 22116 2694 22130 2746
rect 22130 2694 22142 2746
rect 22142 2694 22172 2746
rect 22196 2694 22206 2746
rect 22206 2694 22252 2746
rect 21956 2692 22012 2694
rect 22036 2692 22092 2694
rect 22116 2692 22172 2694
rect 22196 2692 22252 2694
rect 26956 2746 27012 2748
rect 27036 2746 27092 2748
rect 27116 2746 27172 2748
rect 27196 2746 27252 2748
rect 26956 2694 27002 2746
rect 27002 2694 27012 2746
rect 27036 2694 27066 2746
rect 27066 2694 27078 2746
rect 27078 2694 27092 2746
rect 27116 2694 27130 2746
rect 27130 2694 27142 2746
rect 27142 2694 27172 2746
rect 27196 2694 27206 2746
rect 27206 2694 27252 2746
rect 26956 2692 27012 2694
rect 27036 2692 27092 2694
rect 27116 2692 27172 2694
rect 27196 2692 27252 2694
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 36956 2746 37012 2748
rect 37036 2746 37092 2748
rect 37116 2746 37172 2748
rect 37196 2746 37252 2748
rect 36956 2694 37002 2746
rect 37002 2694 37012 2746
rect 37036 2694 37066 2746
rect 37066 2694 37078 2746
rect 37078 2694 37092 2746
rect 37116 2694 37130 2746
rect 37130 2694 37142 2746
rect 37142 2694 37172 2746
rect 37196 2694 37206 2746
rect 37206 2694 37252 2746
rect 36956 2692 37012 2694
rect 37036 2692 37092 2694
rect 37116 2692 37172 2694
rect 37196 2692 37252 2694
rect 41956 2746 42012 2748
rect 42036 2746 42092 2748
rect 42116 2746 42172 2748
rect 42196 2746 42252 2748
rect 41956 2694 42002 2746
rect 42002 2694 42012 2746
rect 42036 2694 42066 2746
rect 42066 2694 42078 2746
rect 42078 2694 42092 2746
rect 42116 2694 42130 2746
rect 42130 2694 42142 2746
rect 42142 2694 42172 2746
rect 42196 2694 42206 2746
rect 42206 2694 42252 2746
rect 41956 2692 42012 2694
rect 42036 2692 42092 2694
rect 42116 2692 42172 2694
rect 42196 2692 42252 2694
rect 46956 2746 47012 2748
rect 47036 2746 47092 2748
rect 47116 2746 47172 2748
rect 47196 2746 47252 2748
rect 46956 2694 47002 2746
rect 47002 2694 47012 2746
rect 47036 2694 47066 2746
rect 47066 2694 47078 2746
rect 47078 2694 47092 2746
rect 47116 2694 47130 2746
rect 47130 2694 47142 2746
rect 47142 2694 47172 2746
rect 47196 2694 47206 2746
rect 47206 2694 47252 2746
rect 46956 2692 47012 2694
rect 47036 2692 47092 2694
rect 47116 2692 47172 2694
rect 47196 2692 47252 2694
rect 51956 2746 52012 2748
rect 52036 2746 52092 2748
rect 52116 2746 52172 2748
rect 52196 2746 52252 2748
rect 51956 2694 52002 2746
rect 52002 2694 52012 2746
rect 52036 2694 52066 2746
rect 52066 2694 52078 2746
rect 52078 2694 52092 2746
rect 52116 2694 52130 2746
rect 52130 2694 52142 2746
rect 52142 2694 52172 2746
rect 52196 2694 52206 2746
rect 52206 2694 52252 2746
rect 51956 2692 52012 2694
rect 52036 2692 52092 2694
rect 52116 2692 52172 2694
rect 52196 2692 52252 2694
rect 56956 2746 57012 2748
rect 57036 2746 57092 2748
rect 57116 2746 57172 2748
rect 57196 2746 57252 2748
rect 56956 2694 57002 2746
rect 57002 2694 57012 2746
rect 57036 2694 57066 2746
rect 57066 2694 57078 2746
rect 57078 2694 57092 2746
rect 57116 2694 57130 2746
rect 57130 2694 57142 2746
rect 57142 2694 57172 2746
rect 57196 2694 57206 2746
rect 57206 2694 57252 2746
rect 56956 2692 57012 2694
rect 57036 2692 57092 2694
rect 57116 2692 57172 2694
rect 57196 2692 57252 2694
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
rect 22616 2202 22672 2204
rect 22696 2202 22752 2204
rect 22776 2202 22832 2204
rect 22856 2202 22912 2204
rect 22616 2150 22662 2202
rect 22662 2150 22672 2202
rect 22696 2150 22726 2202
rect 22726 2150 22738 2202
rect 22738 2150 22752 2202
rect 22776 2150 22790 2202
rect 22790 2150 22802 2202
rect 22802 2150 22832 2202
rect 22856 2150 22866 2202
rect 22866 2150 22912 2202
rect 22616 2148 22672 2150
rect 22696 2148 22752 2150
rect 22776 2148 22832 2150
rect 22856 2148 22912 2150
rect 27616 2202 27672 2204
rect 27696 2202 27752 2204
rect 27776 2202 27832 2204
rect 27856 2202 27912 2204
rect 27616 2150 27662 2202
rect 27662 2150 27672 2202
rect 27696 2150 27726 2202
rect 27726 2150 27738 2202
rect 27738 2150 27752 2202
rect 27776 2150 27790 2202
rect 27790 2150 27802 2202
rect 27802 2150 27832 2202
rect 27856 2150 27866 2202
rect 27866 2150 27912 2202
rect 27616 2148 27672 2150
rect 27696 2148 27752 2150
rect 27776 2148 27832 2150
rect 27856 2148 27912 2150
rect 32616 2202 32672 2204
rect 32696 2202 32752 2204
rect 32776 2202 32832 2204
rect 32856 2202 32912 2204
rect 32616 2150 32662 2202
rect 32662 2150 32672 2202
rect 32696 2150 32726 2202
rect 32726 2150 32738 2202
rect 32738 2150 32752 2202
rect 32776 2150 32790 2202
rect 32790 2150 32802 2202
rect 32802 2150 32832 2202
rect 32856 2150 32866 2202
rect 32866 2150 32912 2202
rect 32616 2148 32672 2150
rect 32696 2148 32752 2150
rect 32776 2148 32832 2150
rect 32856 2148 32912 2150
rect 37616 2202 37672 2204
rect 37696 2202 37752 2204
rect 37776 2202 37832 2204
rect 37856 2202 37912 2204
rect 37616 2150 37662 2202
rect 37662 2150 37672 2202
rect 37696 2150 37726 2202
rect 37726 2150 37738 2202
rect 37738 2150 37752 2202
rect 37776 2150 37790 2202
rect 37790 2150 37802 2202
rect 37802 2150 37832 2202
rect 37856 2150 37866 2202
rect 37866 2150 37912 2202
rect 37616 2148 37672 2150
rect 37696 2148 37752 2150
rect 37776 2148 37832 2150
rect 37856 2148 37912 2150
rect 42616 2202 42672 2204
rect 42696 2202 42752 2204
rect 42776 2202 42832 2204
rect 42856 2202 42912 2204
rect 42616 2150 42662 2202
rect 42662 2150 42672 2202
rect 42696 2150 42726 2202
rect 42726 2150 42738 2202
rect 42738 2150 42752 2202
rect 42776 2150 42790 2202
rect 42790 2150 42802 2202
rect 42802 2150 42832 2202
rect 42856 2150 42866 2202
rect 42866 2150 42912 2202
rect 42616 2148 42672 2150
rect 42696 2148 42752 2150
rect 42776 2148 42832 2150
rect 42856 2148 42912 2150
rect 47616 2202 47672 2204
rect 47696 2202 47752 2204
rect 47776 2202 47832 2204
rect 47856 2202 47912 2204
rect 47616 2150 47662 2202
rect 47662 2150 47672 2202
rect 47696 2150 47726 2202
rect 47726 2150 47738 2202
rect 47738 2150 47752 2202
rect 47776 2150 47790 2202
rect 47790 2150 47802 2202
rect 47802 2150 47832 2202
rect 47856 2150 47866 2202
rect 47866 2150 47912 2202
rect 47616 2148 47672 2150
rect 47696 2148 47752 2150
rect 47776 2148 47832 2150
rect 47856 2148 47912 2150
rect 52616 2202 52672 2204
rect 52696 2202 52752 2204
rect 52776 2202 52832 2204
rect 52856 2202 52912 2204
rect 52616 2150 52662 2202
rect 52662 2150 52672 2202
rect 52696 2150 52726 2202
rect 52726 2150 52738 2202
rect 52738 2150 52752 2202
rect 52776 2150 52790 2202
rect 52790 2150 52802 2202
rect 52802 2150 52832 2202
rect 52856 2150 52866 2202
rect 52866 2150 52912 2202
rect 52616 2148 52672 2150
rect 52696 2148 52752 2150
rect 52776 2148 52832 2150
rect 52856 2148 52912 2150
rect 57616 2202 57672 2204
rect 57696 2202 57752 2204
rect 57776 2202 57832 2204
rect 57856 2202 57912 2204
rect 57616 2150 57662 2202
rect 57662 2150 57672 2202
rect 57696 2150 57726 2202
rect 57726 2150 57738 2202
rect 57738 2150 57752 2202
rect 57776 2150 57790 2202
rect 57790 2150 57802 2202
rect 57802 2150 57832 2202
rect 57856 2150 57866 2202
rect 57866 2150 57912 2202
rect 57616 2148 57672 2150
rect 57696 2148 57752 2150
rect 57776 2148 57832 2150
rect 57856 2148 57912 2150
<< metal3 >>
rect 2606 57696 2922 57697
rect 2606 57632 2612 57696
rect 2676 57632 2692 57696
rect 2756 57632 2772 57696
rect 2836 57632 2852 57696
rect 2916 57632 2922 57696
rect 2606 57631 2922 57632
rect 7606 57696 7922 57697
rect 7606 57632 7612 57696
rect 7676 57632 7692 57696
rect 7756 57632 7772 57696
rect 7836 57632 7852 57696
rect 7916 57632 7922 57696
rect 7606 57631 7922 57632
rect 12606 57696 12922 57697
rect 12606 57632 12612 57696
rect 12676 57632 12692 57696
rect 12756 57632 12772 57696
rect 12836 57632 12852 57696
rect 12916 57632 12922 57696
rect 12606 57631 12922 57632
rect 17606 57696 17922 57697
rect 17606 57632 17612 57696
rect 17676 57632 17692 57696
rect 17756 57632 17772 57696
rect 17836 57632 17852 57696
rect 17916 57632 17922 57696
rect 17606 57631 17922 57632
rect 22606 57696 22922 57697
rect 22606 57632 22612 57696
rect 22676 57632 22692 57696
rect 22756 57632 22772 57696
rect 22836 57632 22852 57696
rect 22916 57632 22922 57696
rect 22606 57631 22922 57632
rect 27606 57696 27922 57697
rect 27606 57632 27612 57696
rect 27676 57632 27692 57696
rect 27756 57632 27772 57696
rect 27836 57632 27852 57696
rect 27916 57632 27922 57696
rect 27606 57631 27922 57632
rect 32606 57696 32922 57697
rect 32606 57632 32612 57696
rect 32676 57632 32692 57696
rect 32756 57632 32772 57696
rect 32836 57632 32852 57696
rect 32916 57632 32922 57696
rect 32606 57631 32922 57632
rect 37606 57696 37922 57697
rect 37606 57632 37612 57696
rect 37676 57632 37692 57696
rect 37756 57632 37772 57696
rect 37836 57632 37852 57696
rect 37916 57632 37922 57696
rect 37606 57631 37922 57632
rect 42606 57696 42922 57697
rect 42606 57632 42612 57696
rect 42676 57632 42692 57696
rect 42756 57632 42772 57696
rect 42836 57632 42852 57696
rect 42916 57632 42922 57696
rect 42606 57631 42922 57632
rect 47606 57696 47922 57697
rect 47606 57632 47612 57696
rect 47676 57632 47692 57696
rect 47756 57632 47772 57696
rect 47836 57632 47852 57696
rect 47916 57632 47922 57696
rect 47606 57631 47922 57632
rect 52606 57696 52922 57697
rect 52606 57632 52612 57696
rect 52676 57632 52692 57696
rect 52756 57632 52772 57696
rect 52836 57632 52852 57696
rect 52916 57632 52922 57696
rect 52606 57631 52922 57632
rect 57606 57696 57922 57697
rect 57606 57632 57612 57696
rect 57676 57632 57692 57696
rect 57756 57632 57772 57696
rect 57836 57632 57852 57696
rect 57916 57632 57922 57696
rect 57606 57631 57922 57632
rect 1946 57152 2262 57153
rect 1946 57088 1952 57152
rect 2016 57088 2032 57152
rect 2096 57088 2112 57152
rect 2176 57088 2192 57152
rect 2256 57088 2262 57152
rect 1946 57087 2262 57088
rect 6946 57152 7262 57153
rect 6946 57088 6952 57152
rect 7016 57088 7032 57152
rect 7096 57088 7112 57152
rect 7176 57088 7192 57152
rect 7256 57088 7262 57152
rect 6946 57087 7262 57088
rect 11946 57152 12262 57153
rect 11946 57088 11952 57152
rect 12016 57088 12032 57152
rect 12096 57088 12112 57152
rect 12176 57088 12192 57152
rect 12256 57088 12262 57152
rect 11946 57087 12262 57088
rect 16946 57152 17262 57153
rect 16946 57088 16952 57152
rect 17016 57088 17032 57152
rect 17096 57088 17112 57152
rect 17176 57088 17192 57152
rect 17256 57088 17262 57152
rect 16946 57087 17262 57088
rect 21946 57152 22262 57153
rect 21946 57088 21952 57152
rect 22016 57088 22032 57152
rect 22096 57088 22112 57152
rect 22176 57088 22192 57152
rect 22256 57088 22262 57152
rect 21946 57087 22262 57088
rect 26946 57152 27262 57153
rect 26946 57088 26952 57152
rect 27016 57088 27032 57152
rect 27096 57088 27112 57152
rect 27176 57088 27192 57152
rect 27256 57088 27262 57152
rect 26946 57087 27262 57088
rect 31946 57152 32262 57153
rect 31946 57088 31952 57152
rect 32016 57088 32032 57152
rect 32096 57088 32112 57152
rect 32176 57088 32192 57152
rect 32256 57088 32262 57152
rect 31946 57087 32262 57088
rect 36946 57152 37262 57153
rect 36946 57088 36952 57152
rect 37016 57088 37032 57152
rect 37096 57088 37112 57152
rect 37176 57088 37192 57152
rect 37256 57088 37262 57152
rect 36946 57087 37262 57088
rect 41946 57152 42262 57153
rect 41946 57088 41952 57152
rect 42016 57088 42032 57152
rect 42096 57088 42112 57152
rect 42176 57088 42192 57152
rect 42256 57088 42262 57152
rect 41946 57087 42262 57088
rect 46946 57152 47262 57153
rect 46946 57088 46952 57152
rect 47016 57088 47032 57152
rect 47096 57088 47112 57152
rect 47176 57088 47192 57152
rect 47256 57088 47262 57152
rect 46946 57087 47262 57088
rect 51946 57152 52262 57153
rect 51946 57088 51952 57152
rect 52016 57088 52032 57152
rect 52096 57088 52112 57152
rect 52176 57088 52192 57152
rect 52256 57088 52262 57152
rect 51946 57087 52262 57088
rect 56946 57152 57262 57153
rect 56946 57088 56952 57152
rect 57016 57088 57032 57152
rect 57096 57088 57112 57152
rect 57176 57088 57192 57152
rect 57256 57088 57262 57152
rect 56946 57087 57262 57088
rect 2606 56608 2922 56609
rect 2606 56544 2612 56608
rect 2676 56544 2692 56608
rect 2756 56544 2772 56608
rect 2836 56544 2852 56608
rect 2916 56544 2922 56608
rect 2606 56543 2922 56544
rect 7606 56608 7922 56609
rect 7606 56544 7612 56608
rect 7676 56544 7692 56608
rect 7756 56544 7772 56608
rect 7836 56544 7852 56608
rect 7916 56544 7922 56608
rect 7606 56543 7922 56544
rect 12606 56608 12922 56609
rect 12606 56544 12612 56608
rect 12676 56544 12692 56608
rect 12756 56544 12772 56608
rect 12836 56544 12852 56608
rect 12916 56544 12922 56608
rect 12606 56543 12922 56544
rect 17606 56608 17922 56609
rect 17606 56544 17612 56608
rect 17676 56544 17692 56608
rect 17756 56544 17772 56608
rect 17836 56544 17852 56608
rect 17916 56544 17922 56608
rect 17606 56543 17922 56544
rect 22606 56608 22922 56609
rect 22606 56544 22612 56608
rect 22676 56544 22692 56608
rect 22756 56544 22772 56608
rect 22836 56544 22852 56608
rect 22916 56544 22922 56608
rect 22606 56543 22922 56544
rect 27606 56608 27922 56609
rect 27606 56544 27612 56608
rect 27676 56544 27692 56608
rect 27756 56544 27772 56608
rect 27836 56544 27852 56608
rect 27916 56544 27922 56608
rect 27606 56543 27922 56544
rect 32606 56608 32922 56609
rect 32606 56544 32612 56608
rect 32676 56544 32692 56608
rect 32756 56544 32772 56608
rect 32836 56544 32852 56608
rect 32916 56544 32922 56608
rect 32606 56543 32922 56544
rect 37606 56608 37922 56609
rect 37606 56544 37612 56608
rect 37676 56544 37692 56608
rect 37756 56544 37772 56608
rect 37836 56544 37852 56608
rect 37916 56544 37922 56608
rect 37606 56543 37922 56544
rect 42606 56608 42922 56609
rect 42606 56544 42612 56608
rect 42676 56544 42692 56608
rect 42756 56544 42772 56608
rect 42836 56544 42852 56608
rect 42916 56544 42922 56608
rect 42606 56543 42922 56544
rect 47606 56608 47922 56609
rect 47606 56544 47612 56608
rect 47676 56544 47692 56608
rect 47756 56544 47772 56608
rect 47836 56544 47852 56608
rect 47916 56544 47922 56608
rect 47606 56543 47922 56544
rect 52606 56608 52922 56609
rect 52606 56544 52612 56608
rect 52676 56544 52692 56608
rect 52756 56544 52772 56608
rect 52836 56544 52852 56608
rect 52916 56544 52922 56608
rect 52606 56543 52922 56544
rect 57606 56608 57922 56609
rect 57606 56544 57612 56608
rect 57676 56544 57692 56608
rect 57756 56544 57772 56608
rect 57836 56544 57852 56608
rect 57916 56544 57922 56608
rect 57606 56543 57922 56544
rect 1946 56064 2262 56065
rect 1946 56000 1952 56064
rect 2016 56000 2032 56064
rect 2096 56000 2112 56064
rect 2176 56000 2192 56064
rect 2256 56000 2262 56064
rect 1946 55999 2262 56000
rect 6946 56064 7262 56065
rect 6946 56000 6952 56064
rect 7016 56000 7032 56064
rect 7096 56000 7112 56064
rect 7176 56000 7192 56064
rect 7256 56000 7262 56064
rect 6946 55999 7262 56000
rect 11946 56064 12262 56065
rect 11946 56000 11952 56064
rect 12016 56000 12032 56064
rect 12096 56000 12112 56064
rect 12176 56000 12192 56064
rect 12256 56000 12262 56064
rect 11946 55999 12262 56000
rect 16946 56064 17262 56065
rect 16946 56000 16952 56064
rect 17016 56000 17032 56064
rect 17096 56000 17112 56064
rect 17176 56000 17192 56064
rect 17256 56000 17262 56064
rect 16946 55999 17262 56000
rect 21946 56064 22262 56065
rect 21946 56000 21952 56064
rect 22016 56000 22032 56064
rect 22096 56000 22112 56064
rect 22176 56000 22192 56064
rect 22256 56000 22262 56064
rect 21946 55999 22262 56000
rect 26946 56064 27262 56065
rect 26946 56000 26952 56064
rect 27016 56000 27032 56064
rect 27096 56000 27112 56064
rect 27176 56000 27192 56064
rect 27256 56000 27262 56064
rect 26946 55999 27262 56000
rect 31946 56064 32262 56065
rect 31946 56000 31952 56064
rect 32016 56000 32032 56064
rect 32096 56000 32112 56064
rect 32176 56000 32192 56064
rect 32256 56000 32262 56064
rect 31946 55999 32262 56000
rect 36946 56064 37262 56065
rect 36946 56000 36952 56064
rect 37016 56000 37032 56064
rect 37096 56000 37112 56064
rect 37176 56000 37192 56064
rect 37256 56000 37262 56064
rect 36946 55999 37262 56000
rect 41946 56064 42262 56065
rect 41946 56000 41952 56064
rect 42016 56000 42032 56064
rect 42096 56000 42112 56064
rect 42176 56000 42192 56064
rect 42256 56000 42262 56064
rect 41946 55999 42262 56000
rect 46946 56064 47262 56065
rect 46946 56000 46952 56064
rect 47016 56000 47032 56064
rect 47096 56000 47112 56064
rect 47176 56000 47192 56064
rect 47256 56000 47262 56064
rect 46946 55999 47262 56000
rect 51946 56064 52262 56065
rect 51946 56000 51952 56064
rect 52016 56000 52032 56064
rect 52096 56000 52112 56064
rect 52176 56000 52192 56064
rect 52256 56000 52262 56064
rect 51946 55999 52262 56000
rect 56946 56064 57262 56065
rect 56946 56000 56952 56064
rect 57016 56000 57032 56064
rect 57096 56000 57112 56064
rect 57176 56000 57192 56064
rect 57256 56000 57262 56064
rect 56946 55999 57262 56000
rect 58525 55586 58591 55589
rect 59200 55586 60000 55616
rect 58525 55584 60000 55586
rect 58525 55528 58530 55584
rect 58586 55528 60000 55584
rect 58525 55526 60000 55528
rect 58525 55523 58591 55526
rect 2606 55520 2922 55521
rect 2606 55456 2612 55520
rect 2676 55456 2692 55520
rect 2756 55456 2772 55520
rect 2836 55456 2852 55520
rect 2916 55456 2922 55520
rect 2606 55455 2922 55456
rect 7606 55520 7922 55521
rect 7606 55456 7612 55520
rect 7676 55456 7692 55520
rect 7756 55456 7772 55520
rect 7836 55456 7852 55520
rect 7916 55456 7922 55520
rect 7606 55455 7922 55456
rect 12606 55520 12922 55521
rect 12606 55456 12612 55520
rect 12676 55456 12692 55520
rect 12756 55456 12772 55520
rect 12836 55456 12852 55520
rect 12916 55456 12922 55520
rect 12606 55455 12922 55456
rect 17606 55520 17922 55521
rect 17606 55456 17612 55520
rect 17676 55456 17692 55520
rect 17756 55456 17772 55520
rect 17836 55456 17852 55520
rect 17916 55456 17922 55520
rect 17606 55455 17922 55456
rect 22606 55520 22922 55521
rect 22606 55456 22612 55520
rect 22676 55456 22692 55520
rect 22756 55456 22772 55520
rect 22836 55456 22852 55520
rect 22916 55456 22922 55520
rect 22606 55455 22922 55456
rect 27606 55520 27922 55521
rect 27606 55456 27612 55520
rect 27676 55456 27692 55520
rect 27756 55456 27772 55520
rect 27836 55456 27852 55520
rect 27916 55456 27922 55520
rect 27606 55455 27922 55456
rect 32606 55520 32922 55521
rect 32606 55456 32612 55520
rect 32676 55456 32692 55520
rect 32756 55456 32772 55520
rect 32836 55456 32852 55520
rect 32916 55456 32922 55520
rect 32606 55455 32922 55456
rect 37606 55520 37922 55521
rect 37606 55456 37612 55520
rect 37676 55456 37692 55520
rect 37756 55456 37772 55520
rect 37836 55456 37852 55520
rect 37916 55456 37922 55520
rect 37606 55455 37922 55456
rect 42606 55520 42922 55521
rect 42606 55456 42612 55520
rect 42676 55456 42692 55520
rect 42756 55456 42772 55520
rect 42836 55456 42852 55520
rect 42916 55456 42922 55520
rect 42606 55455 42922 55456
rect 47606 55520 47922 55521
rect 47606 55456 47612 55520
rect 47676 55456 47692 55520
rect 47756 55456 47772 55520
rect 47836 55456 47852 55520
rect 47916 55456 47922 55520
rect 47606 55455 47922 55456
rect 52606 55520 52922 55521
rect 52606 55456 52612 55520
rect 52676 55456 52692 55520
rect 52756 55456 52772 55520
rect 52836 55456 52852 55520
rect 52916 55456 52922 55520
rect 52606 55455 52922 55456
rect 57606 55520 57922 55521
rect 57606 55456 57612 55520
rect 57676 55456 57692 55520
rect 57756 55456 57772 55520
rect 57836 55456 57852 55520
rect 57916 55456 57922 55520
rect 59200 55496 60000 55526
rect 57606 55455 57922 55456
rect 1946 54976 2262 54977
rect 1946 54912 1952 54976
rect 2016 54912 2032 54976
rect 2096 54912 2112 54976
rect 2176 54912 2192 54976
rect 2256 54912 2262 54976
rect 1946 54911 2262 54912
rect 6946 54976 7262 54977
rect 6946 54912 6952 54976
rect 7016 54912 7032 54976
rect 7096 54912 7112 54976
rect 7176 54912 7192 54976
rect 7256 54912 7262 54976
rect 6946 54911 7262 54912
rect 11946 54976 12262 54977
rect 11946 54912 11952 54976
rect 12016 54912 12032 54976
rect 12096 54912 12112 54976
rect 12176 54912 12192 54976
rect 12256 54912 12262 54976
rect 11946 54911 12262 54912
rect 16946 54976 17262 54977
rect 16946 54912 16952 54976
rect 17016 54912 17032 54976
rect 17096 54912 17112 54976
rect 17176 54912 17192 54976
rect 17256 54912 17262 54976
rect 16946 54911 17262 54912
rect 21946 54976 22262 54977
rect 21946 54912 21952 54976
rect 22016 54912 22032 54976
rect 22096 54912 22112 54976
rect 22176 54912 22192 54976
rect 22256 54912 22262 54976
rect 21946 54911 22262 54912
rect 26946 54976 27262 54977
rect 26946 54912 26952 54976
rect 27016 54912 27032 54976
rect 27096 54912 27112 54976
rect 27176 54912 27192 54976
rect 27256 54912 27262 54976
rect 26946 54911 27262 54912
rect 31946 54976 32262 54977
rect 31946 54912 31952 54976
rect 32016 54912 32032 54976
rect 32096 54912 32112 54976
rect 32176 54912 32192 54976
rect 32256 54912 32262 54976
rect 31946 54911 32262 54912
rect 36946 54976 37262 54977
rect 36946 54912 36952 54976
rect 37016 54912 37032 54976
rect 37096 54912 37112 54976
rect 37176 54912 37192 54976
rect 37256 54912 37262 54976
rect 36946 54911 37262 54912
rect 41946 54976 42262 54977
rect 41946 54912 41952 54976
rect 42016 54912 42032 54976
rect 42096 54912 42112 54976
rect 42176 54912 42192 54976
rect 42256 54912 42262 54976
rect 41946 54911 42262 54912
rect 46946 54976 47262 54977
rect 46946 54912 46952 54976
rect 47016 54912 47032 54976
rect 47096 54912 47112 54976
rect 47176 54912 47192 54976
rect 47256 54912 47262 54976
rect 46946 54911 47262 54912
rect 51946 54976 52262 54977
rect 51946 54912 51952 54976
rect 52016 54912 52032 54976
rect 52096 54912 52112 54976
rect 52176 54912 52192 54976
rect 52256 54912 52262 54976
rect 51946 54911 52262 54912
rect 56946 54976 57262 54977
rect 56946 54912 56952 54976
rect 57016 54912 57032 54976
rect 57096 54912 57112 54976
rect 57176 54912 57192 54976
rect 57256 54912 57262 54976
rect 56946 54911 57262 54912
rect 58525 54770 58591 54773
rect 59200 54770 60000 54800
rect 58525 54768 60000 54770
rect 58525 54712 58530 54768
rect 58586 54712 60000 54768
rect 58525 54710 60000 54712
rect 58525 54707 58591 54710
rect 59200 54680 60000 54710
rect 2606 54432 2922 54433
rect 2606 54368 2612 54432
rect 2676 54368 2692 54432
rect 2756 54368 2772 54432
rect 2836 54368 2852 54432
rect 2916 54368 2922 54432
rect 2606 54367 2922 54368
rect 7606 54432 7922 54433
rect 7606 54368 7612 54432
rect 7676 54368 7692 54432
rect 7756 54368 7772 54432
rect 7836 54368 7852 54432
rect 7916 54368 7922 54432
rect 7606 54367 7922 54368
rect 12606 54432 12922 54433
rect 12606 54368 12612 54432
rect 12676 54368 12692 54432
rect 12756 54368 12772 54432
rect 12836 54368 12852 54432
rect 12916 54368 12922 54432
rect 12606 54367 12922 54368
rect 17606 54432 17922 54433
rect 17606 54368 17612 54432
rect 17676 54368 17692 54432
rect 17756 54368 17772 54432
rect 17836 54368 17852 54432
rect 17916 54368 17922 54432
rect 17606 54367 17922 54368
rect 22606 54432 22922 54433
rect 22606 54368 22612 54432
rect 22676 54368 22692 54432
rect 22756 54368 22772 54432
rect 22836 54368 22852 54432
rect 22916 54368 22922 54432
rect 22606 54367 22922 54368
rect 27606 54432 27922 54433
rect 27606 54368 27612 54432
rect 27676 54368 27692 54432
rect 27756 54368 27772 54432
rect 27836 54368 27852 54432
rect 27916 54368 27922 54432
rect 27606 54367 27922 54368
rect 32606 54432 32922 54433
rect 32606 54368 32612 54432
rect 32676 54368 32692 54432
rect 32756 54368 32772 54432
rect 32836 54368 32852 54432
rect 32916 54368 32922 54432
rect 32606 54367 32922 54368
rect 37606 54432 37922 54433
rect 37606 54368 37612 54432
rect 37676 54368 37692 54432
rect 37756 54368 37772 54432
rect 37836 54368 37852 54432
rect 37916 54368 37922 54432
rect 37606 54367 37922 54368
rect 42606 54432 42922 54433
rect 42606 54368 42612 54432
rect 42676 54368 42692 54432
rect 42756 54368 42772 54432
rect 42836 54368 42852 54432
rect 42916 54368 42922 54432
rect 42606 54367 42922 54368
rect 47606 54432 47922 54433
rect 47606 54368 47612 54432
rect 47676 54368 47692 54432
rect 47756 54368 47772 54432
rect 47836 54368 47852 54432
rect 47916 54368 47922 54432
rect 47606 54367 47922 54368
rect 52606 54432 52922 54433
rect 52606 54368 52612 54432
rect 52676 54368 52692 54432
rect 52756 54368 52772 54432
rect 52836 54368 52852 54432
rect 52916 54368 52922 54432
rect 52606 54367 52922 54368
rect 57606 54432 57922 54433
rect 57606 54368 57612 54432
rect 57676 54368 57692 54432
rect 57756 54368 57772 54432
rect 57836 54368 57852 54432
rect 57916 54368 57922 54432
rect 57606 54367 57922 54368
rect 58525 53954 58591 53957
rect 59200 53954 60000 53984
rect 58525 53952 60000 53954
rect 58525 53896 58530 53952
rect 58586 53896 60000 53952
rect 58525 53894 60000 53896
rect 58525 53891 58591 53894
rect 1946 53888 2262 53889
rect 1946 53824 1952 53888
rect 2016 53824 2032 53888
rect 2096 53824 2112 53888
rect 2176 53824 2192 53888
rect 2256 53824 2262 53888
rect 1946 53823 2262 53824
rect 6946 53888 7262 53889
rect 6946 53824 6952 53888
rect 7016 53824 7032 53888
rect 7096 53824 7112 53888
rect 7176 53824 7192 53888
rect 7256 53824 7262 53888
rect 6946 53823 7262 53824
rect 11946 53888 12262 53889
rect 11946 53824 11952 53888
rect 12016 53824 12032 53888
rect 12096 53824 12112 53888
rect 12176 53824 12192 53888
rect 12256 53824 12262 53888
rect 11946 53823 12262 53824
rect 16946 53888 17262 53889
rect 16946 53824 16952 53888
rect 17016 53824 17032 53888
rect 17096 53824 17112 53888
rect 17176 53824 17192 53888
rect 17256 53824 17262 53888
rect 16946 53823 17262 53824
rect 21946 53888 22262 53889
rect 21946 53824 21952 53888
rect 22016 53824 22032 53888
rect 22096 53824 22112 53888
rect 22176 53824 22192 53888
rect 22256 53824 22262 53888
rect 21946 53823 22262 53824
rect 26946 53888 27262 53889
rect 26946 53824 26952 53888
rect 27016 53824 27032 53888
rect 27096 53824 27112 53888
rect 27176 53824 27192 53888
rect 27256 53824 27262 53888
rect 26946 53823 27262 53824
rect 31946 53888 32262 53889
rect 31946 53824 31952 53888
rect 32016 53824 32032 53888
rect 32096 53824 32112 53888
rect 32176 53824 32192 53888
rect 32256 53824 32262 53888
rect 31946 53823 32262 53824
rect 36946 53888 37262 53889
rect 36946 53824 36952 53888
rect 37016 53824 37032 53888
rect 37096 53824 37112 53888
rect 37176 53824 37192 53888
rect 37256 53824 37262 53888
rect 36946 53823 37262 53824
rect 41946 53888 42262 53889
rect 41946 53824 41952 53888
rect 42016 53824 42032 53888
rect 42096 53824 42112 53888
rect 42176 53824 42192 53888
rect 42256 53824 42262 53888
rect 41946 53823 42262 53824
rect 46946 53888 47262 53889
rect 46946 53824 46952 53888
rect 47016 53824 47032 53888
rect 47096 53824 47112 53888
rect 47176 53824 47192 53888
rect 47256 53824 47262 53888
rect 46946 53823 47262 53824
rect 51946 53888 52262 53889
rect 51946 53824 51952 53888
rect 52016 53824 52032 53888
rect 52096 53824 52112 53888
rect 52176 53824 52192 53888
rect 52256 53824 52262 53888
rect 51946 53823 52262 53824
rect 56946 53888 57262 53889
rect 56946 53824 56952 53888
rect 57016 53824 57032 53888
rect 57096 53824 57112 53888
rect 57176 53824 57192 53888
rect 57256 53824 57262 53888
rect 59200 53864 60000 53894
rect 56946 53823 57262 53824
rect 2606 53344 2922 53345
rect 2606 53280 2612 53344
rect 2676 53280 2692 53344
rect 2756 53280 2772 53344
rect 2836 53280 2852 53344
rect 2916 53280 2922 53344
rect 2606 53279 2922 53280
rect 7606 53344 7922 53345
rect 7606 53280 7612 53344
rect 7676 53280 7692 53344
rect 7756 53280 7772 53344
rect 7836 53280 7852 53344
rect 7916 53280 7922 53344
rect 7606 53279 7922 53280
rect 12606 53344 12922 53345
rect 12606 53280 12612 53344
rect 12676 53280 12692 53344
rect 12756 53280 12772 53344
rect 12836 53280 12852 53344
rect 12916 53280 12922 53344
rect 12606 53279 12922 53280
rect 17606 53344 17922 53345
rect 17606 53280 17612 53344
rect 17676 53280 17692 53344
rect 17756 53280 17772 53344
rect 17836 53280 17852 53344
rect 17916 53280 17922 53344
rect 17606 53279 17922 53280
rect 22606 53344 22922 53345
rect 22606 53280 22612 53344
rect 22676 53280 22692 53344
rect 22756 53280 22772 53344
rect 22836 53280 22852 53344
rect 22916 53280 22922 53344
rect 22606 53279 22922 53280
rect 27606 53344 27922 53345
rect 27606 53280 27612 53344
rect 27676 53280 27692 53344
rect 27756 53280 27772 53344
rect 27836 53280 27852 53344
rect 27916 53280 27922 53344
rect 27606 53279 27922 53280
rect 32606 53344 32922 53345
rect 32606 53280 32612 53344
rect 32676 53280 32692 53344
rect 32756 53280 32772 53344
rect 32836 53280 32852 53344
rect 32916 53280 32922 53344
rect 32606 53279 32922 53280
rect 37606 53344 37922 53345
rect 37606 53280 37612 53344
rect 37676 53280 37692 53344
rect 37756 53280 37772 53344
rect 37836 53280 37852 53344
rect 37916 53280 37922 53344
rect 37606 53279 37922 53280
rect 42606 53344 42922 53345
rect 42606 53280 42612 53344
rect 42676 53280 42692 53344
rect 42756 53280 42772 53344
rect 42836 53280 42852 53344
rect 42916 53280 42922 53344
rect 42606 53279 42922 53280
rect 47606 53344 47922 53345
rect 47606 53280 47612 53344
rect 47676 53280 47692 53344
rect 47756 53280 47772 53344
rect 47836 53280 47852 53344
rect 47916 53280 47922 53344
rect 47606 53279 47922 53280
rect 52606 53344 52922 53345
rect 52606 53280 52612 53344
rect 52676 53280 52692 53344
rect 52756 53280 52772 53344
rect 52836 53280 52852 53344
rect 52916 53280 52922 53344
rect 52606 53279 52922 53280
rect 57606 53344 57922 53345
rect 57606 53280 57612 53344
rect 57676 53280 57692 53344
rect 57756 53280 57772 53344
rect 57836 53280 57852 53344
rect 57916 53280 57922 53344
rect 57606 53279 57922 53280
rect 58525 53138 58591 53141
rect 59200 53138 60000 53168
rect 58525 53136 60000 53138
rect 58525 53080 58530 53136
rect 58586 53080 60000 53136
rect 58525 53078 60000 53080
rect 58525 53075 58591 53078
rect 59200 53048 60000 53078
rect 1946 52800 2262 52801
rect 1946 52736 1952 52800
rect 2016 52736 2032 52800
rect 2096 52736 2112 52800
rect 2176 52736 2192 52800
rect 2256 52736 2262 52800
rect 1946 52735 2262 52736
rect 6946 52800 7262 52801
rect 6946 52736 6952 52800
rect 7016 52736 7032 52800
rect 7096 52736 7112 52800
rect 7176 52736 7192 52800
rect 7256 52736 7262 52800
rect 6946 52735 7262 52736
rect 11946 52800 12262 52801
rect 11946 52736 11952 52800
rect 12016 52736 12032 52800
rect 12096 52736 12112 52800
rect 12176 52736 12192 52800
rect 12256 52736 12262 52800
rect 11946 52735 12262 52736
rect 16946 52800 17262 52801
rect 16946 52736 16952 52800
rect 17016 52736 17032 52800
rect 17096 52736 17112 52800
rect 17176 52736 17192 52800
rect 17256 52736 17262 52800
rect 16946 52735 17262 52736
rect 21946 52800 22262 52801
rect 21946 52736 21952 52800
rect 22016 52736 22032 52800
rect 22096 52736 22112 52800
rect 22176 52736 22192 52800
rect 22256 52736 22262 52800
rect 21946 52735 22262 52736
rect 26946 52800 27262 52801
rect 26946 52736 26952 52800
rect 27016 52736 27032 52800
rect 27096 52736 27112 52800
rect 27176 52736 27192 52800
rect 27256 52736 27262 52800
rect 26946 52735 27262 52736
rect 31946 52800 32262 52801
rect 31946 52736 31952 52800
rect 32016 52736 32032 52800
rect 32096 52736 32112 52800
rect 32176 52736 32192 52800
rect 32256 52736 32262 52800
rect 31946 52735 32262 52736
rect 36946 52800 37262 52801
rect 36946 52736 36952 52800
rect 37016 52736 37032 52800
rect 37096 52736 37112 52800
rect 37176 52736 37192 52800
rect 37256 52736 37262 52800
rect 36946 52735 37262 52736
rect 41946 52800 42262 52801
rect 41946 52736 41952 52800
rect 42016 52736 42032 52800
rect 42096 52736 42112 52800
rect 42176 52736 42192 52800
rect 42256 52736 42262 52800
rect 41946 52735 42262 52736
rect 46946 52800 47262 52801
rect 46946 52736 46952 52800
rect 47016 52736 47032 52800
rect 47096 52736 47112 52800
rect 47176 52736 47192 52800
rect 47256 52736 47262 52800
rect 46946 52735 47262 52736
rect 51946 52800 52262 52801
rect 51946 52736 51952 52800
rect 52016 52736 52032 52800
rect 52096 52736 52112 52800
rect 52176 52736 52192 52800
rect 52256 52736 52262 52800
rect 51946 52735 52262 52736
rect 56946 52800 57262 52801
rect 56946 52736 56952 52800
rect 57016 52736 57032 52800
rect 57096 52736 57112 52800
rect 57176 52736 57192 52800
rect 57256 52736 57262 52800
rect 56946 52735 57262 52736
rect 58525 52322 58591 52325
rect 59200 52322 60000 52352
rect 58525 52320 60000 52322
rect 58525 52264 58530 52320
rect 58586 52264 60000 52320
rect 58525 52262 60000 52264
rect 58525 52259 58591 52262
rect 2606 52256 2922 52257
rect 2606 52192 2612 52256
rect 2676 52192 2692 52256
rect 2756 52192 2772 52256
rect 2836 52192 2852 52256
rect 2916 52192 2922 52256
rect 2606 52191 2922 52192
rect 7606 52256 7922 52257
rect 7606 52192 7612 52256
rect 7676 52192 7692 52256
rect 7756 52192 7772 52256
rect 7836 52192 7852 52256
rect 7916 52192 7922 52256
rect 7606 52191 7922 52192
rect 12606 52256 12922 52257
rect 12606 52192 12612 52256
rect 12676 52192 12692 52256
rect 12756 52192 12772 52256
rect 12836 52192 12852 52256
rect 12916 52192 12922 52256
rect 12606 52191 12922 52192
rect 17606 52256 17922 52257
rect 17606 52192 17612 52256
rect 17676 52192 17692 52256
rect 17756 52192 17772 52256
rect 17836 52192 17852 52256
rect 17916 52192 17922 52256
rect 17606 52191 17922 52192
rect 22606 52256 22922 52257
rect 22606 52192 22612 52256
rect 22676 52192 22692 52256
rect 22756 52192 22772 52256
rect 22836 52192 22852 52256
rect 22916 52192 22922 52256
rect 22606 52191 22922 52192
rect 27606 52256 27922 52257
rect 27606 52192 27612 52256
rect 27676 52192 27692 52256
rect 27756 52192 27772 52256
rect 27836 52192 27852 52256
rect 27916 52192 27922 52256
rect 27606 52191 27922 52192
rect 32606 52256 32922 52257
rect 32606 52192 32612 52256
rect 32676 52192 32692 52256
rect 32756 52192 32772 52256
rect 32836 52192 32852 52256
rect 32916 52192 32922 52256
rect 32606 52191 32922 52192
rect 37606 52256 37922 52257
rect 37606 52192 37612 52256
rect 37676 52192 37692 52256
rect 37756 52192 37772 52256
rect 37836 52192 37852 52256
rect 37916 52192 37922 52256
rect 37606 52191 37922 52192
rect 42606 52256 42922 52257
rect 42606 52192 42612 52256
rect 42676 52192 42692 52256
rect 42756 52192 42772 52256
rect 42836 52192 42852 52256
rect 42916 52192 42922 52256
rect 42606 52191 42922 52192
rect 47606 52256 47922 52257
rect 47606 52192 47612 52256
rect 47676 52192 47692 52256
rect 47756 52192 47772 52256
rect 47836 52192 47852 52256
rect 47916 52192 47922 52256
rect 47606 52191 47922 52192
rect 52606 52256 52922 52257
rect 52606 52192 52612 52256
rect 52676 52192 52692 52256
rect 52756 52192 52772 52256
rect 52836 52192 52852 52256
rect 52916 52192 52922 52256
rect 52606 52191 52922 52192
rect 57606 52256 57922 52257
rect 57606 52192 57612 52256
rect 57676 52192 57692 52256
rect 57756 52192 57772 52256
rect 57836 52192 57852 52256
rect 57916 52192 57922 52256
rect 59200 52232 60000 52262
rect 57606 52191 57922 52192
rect 1946 51712 2262 51713
rect 1946 51648 1952 51712
rect 2016 51648 2032 51712
rect 2096 51648 2112 51712
rect 2176 51648 2192 51712
rect 2256 51648 2262 51712
rect 1946 51647 2262 51648
rect 6946 51712 7262 51713
rect 6946 51648 6952 51712
rect 7016 51648 7032 51712
rect 7096 51648 7112 51712
rect 7176 51648 7192 51712
rect 7256 51648 7262 51712
rect 6946 51647 7262 51648
rect 11946 51712 12262 51713
rect 11946 51648 11952 51712
rect 12016 51648 12032 51712
rect 12096 51648 12112 51712
rect 12176 51648 12192 51712
rect 12256 51648 12262 51712
rect 11946 51647 12262 51648
rect 16946 51712 17262 51713
rect 16946 51648 16952 51712
rect 17016 51648 17032 51712
rect 17096 51648 17112 51712
rect 17176 51648 17192 51712
rect 17256 51648 17262 51712
rect 16946 51647 17262 51648
rect 21946 51712 22262 51713
rect 21946 51648 21952 51712
rect 22016 51648 22032 51712
rect 22096 51648 22112 51712
rect 22176 51648 22192 51712
rect 22256 51648 22262 51712
rect 21946 51647 22262 51648
rect 26946 51712 27262 51713
rect 26946 51648 26952 51712
rect 27016 51648 27032 51712
rect 27096 51648 27112 51712
rect 27176 51648 27192 51712
rect 27256 51648 27262 51712
rect 26946 51647 27262 51648
rect 31946 51712 32262 51713
rect 31946 51648 31952 51712
rect 32016 51648 32032 51712
rect 32096 51648 32112 51712
rect 32176 51648 32192 51712
rect 32256 51648 32262 51712
rect 31946 51647 32262 51648
rect 36946 51712 37262 51713
rect 36946 51648 36952 51712
rect 37016 51648 37032 51712
rect 37096 51648 37112 51712
rect 37176 51648 37192 51712
rect 37256 51648 37262 51712
rect 36946 51647 37262 51648
rect 41946 51712 42262 51713
rect 41946 51648 41952 51712
rect 42016 51648 42032 51712
rect 42096 51648 42112 51712
rect 42176 51648 42192 51712
rect 42256 51648 42262 51712
rect 41946 51647 42262 51648
rect 46946 51712 47262 51713
rect 46946 51648 46952 51712
rect 47016 51648 47032 51712
rect 47096 51648 47112 51712
rect 47176 51648 47192 51712
rect 47256 51648 47262 51712
rect 46946 51647 47262 51648
rect 51946 51712 52262 51713
rect 51946 51648 51952 51712
rect 52016 51648 52032 51712
rect 52096 51648 52112 51712
rect 52176 51648 52192 51712
rect 52256 51648 52262 51712
rect 51946 51647 52262 51648
rect 56946 51712 57262 51713
rect 56946 51648 56952 51712
rect 57016 51648 57032 51712
rect 57096 51648 57112 51712
rect 57176 51648 57192 51712
rect 57256 51648 57262 51712
rect 56946 51647 57262 51648
rect 58525 51506 58591 51509
rect 59200 51506 60000 51536
rect 58525 51504 60000 51506
rect 58525 51448 58530 51504
rect 58586 51448 60000 51504
rect 58525 51446 60000 51448
rect 58525 51443 58591 51446
rect 59200 51416 60000 51446
rect 2606 51168 2922 51169
rect 2606 51104 2612 51168
rect 2676 51104 2692 51168
rect 2756 51104 2772 51168
rect 2836 51104 2852 51168
rect 2916 51104 2922 51168
rect 2606 51103 2922 51104
rect 7606 51168 7922 51169
rect 7606 51104 7612 51168
rect 7676 51104 7692 51168
rect 7756 51104 7772 51168
rect 7836 51104 7852 51168
rect 7916 51104 7922 51168
rect 7606 51103 7922 51104
rect 12606 51168 12922 51169
rect 12606 51104 12612 51168
rect 12676 51104 12692 51168
rect 12756 51104 12772 51168
rect 12836 51104 12852 51168
rect 12916 51104 12922 51168
rect 12606 51103 12922 51104
rect 17606 51168 17922 51169
rect 17606 51104 17612 51168
rect 17676 51104 17692 51168
rect 17756 51104 17772 51168
rect 17836 51104 17852 51168
rect 17916 51104 17922 51168
rect 17606 51103 17922 51104
rect 22606 51168 22922 51169
rect 22606 51104 22612 51168
rect 22676 51104 22692 51168
rect 22756 51104 22772 51168
rect 22836 51104 22852 51168
rect 22916 51104 22922 51168
rect 22606 51103 22922 51104
rect 27606 51168 27922 51169
rect 27606 51104 27612 51168
rect 27676 51104 27692 51168
rect 27756 51104 27772 51168
rect 27836 51104 27852 51168
rect 27916 51104 27922 51168
rect 27606 51103 27922 51104
rect 32606 51168 32922 51169
rect 32606 51104 32612 51168
rect 32676 51104 32692 51168
rect 32756 51104 32772 51168
rect 32836 51104 32852 51168
rect 32916 51104 32922 51168
rect 32606 51103 32922 51104
rect 37606 51168 37922 51169
rect 37606 51104 37612 51168
rect 37676 51104 37692 51168
rect 37756 51104 37772 51168
rect 37836 51104 37852 51168
rect 37916 51104 37922 51168
rect 37606 51103 37922 51104
rect 42606 51168 42922 51169
rect 42606 51104 42612 51168
rect 42676 51104 42692 51168
rect 42756 51104 42772 51168
rect 42836 51104 42852 51168
rect 42916 51104 42922 51168
rect 42606 51103 42922 51104
rect 47606 51168 47922 51169
rect 47606 51104 47612 51168
rect 47676 51104 47692 51168
rect 47756 51104 47772 51168
rect 47836 51104 47852 51168
rect 47916 51104 47922 51168
rect 47606 51103 47922 51104
rect 52606 51168 52922 51169
rect 52606 51104 52612 51168
rect 52676 51104 52692 51168
rect 52756 51104 52772 51168
rect 52836 51104 52852 51168
rect 52916 51104 52922 51168
rect 52606 51103 52922 51104
rect 57606 51168 57922 51169
rect 57606 51104 57612 51168
rect 57676 51104 57692 51168
rect 57756 51104 57772 51168
rect 57836 51104 57852 51168
rect 57916 51104 57922 51168
rect 57606 51103 57922 51104
rect 58525 50690 58591 50693
rect 59200 50690 60000 50720
rect 58525 50688 60000 50690
rect 58525 50632 58530 50688
rect 58586 50632 60000 50688
rect 58525 50630 60000 50632
rect 58525 50627 58591 50630
rect 1946 50624 2262 50625
rect 1946 50560 1952 50624
rect 2016 50560 2032 50624
rect 2096 50560 2112 50624
rect 2176 50560 2192 50624
rect 2256 50560 2262 50624
rect 1946 50559 2262 50560
rect 6946 50624 7262 50625
rect 6946 50560 6952 50624
rect 7016 50560 7032 50624
rect 7096 50560 7112 50624
rect 7176 50560 7192 50624
rect 7256 50560 7262 50624
rect 6946 50559 7262 50560
rect 11946 50624 12262 50625
rect 11946 50560 11952 50624
rect 12016 50560 12032 50624
rect 12096 50560 12112 50624
rect 12176 50560 12192 50624
rect 12256 50560 12262 50624
rect 11946 50559 12262 50560
rect 16946 50624 17262 50625
rect 16946 50560 16952 50624
rect 17016 50560 17032 50624
rect 17096 50560 17112 50624
rect 17176 50560 17192 50624
rect 17256 50560 17262 50624
rect 16946 50559 17262 50560
rect 21946 50624 22262 50625
rect 21946 50560 21952 50624
rect 22016 50560 22032 50624
rect 22096 50560 22112 50624
rect 22176 50560 22192 50624
rect 22256 50560 22262 50624
rect 21946 50559 22262 50560
rect 26946 50624 27262 50625
rect 26946 50560 26952 50624
rect 27016 50560 27032 50624
rect 27096 50560 27112 50624
rect 27176 50560 27192 50624
rect 27256 50560 27262 50624
rect 26946 50559 27262 50560
rect 31946 50624 32262 50625
rect 31946 50560 31952 50624
rect 32016 50560 32032 50624
rect 32096 50560 32112 50624
rect 32176 50560 32192 50624
rect 32256 50560 32262 50624
rect 31946 50559 32262 50560
rect 36946 50624 37262 50625
rect 36946 50560 36952 50624
rect 37016 50560 37032 50624
rect 37096 50560 37112 50624
rect 37176 50560 37192 50624
rect 37256 50560 37262 50624
rect 36946 50559 37262 50560
rect 41946 50624 42262 50625
rect 41946 50560 41952 50624
rect 42016 50560 42032 50624
rect 42096 50560 42112 50624
rect 42176 50560 42192 50624
rect 42256 50560 42262 50624
rect 41946 50559 42262 50560
rect 46946 50624 47262 50625
rect 46946 50560 46952 50624
rect 47016 50560 47032 50624
rect 47096 50560 47112 50624
rect 47176 50560 47192 50624
rect 47256 50560 47262 50624
rect 46946 50559 47262 50560
rect 51946 50624 52262 50625
rect 51946 50560 51952 50624
rect 52016 50560 52032 50624
rect 52096 50560 52112 50624
rect 52176 50560 52192 50624
rect 52256 50560 52262 50624
rect 51946 50559 52262 50560
rect 56946 50624 57262 50625
rect 56946 50560 56952 50624
rect 57016 50560 57032 50624
rect 57096 50560 57112 50624
rect 57176 50560 57192 50624
rect 57256 50560 57262 50624
rect 59200 50600 60000 50630
rect 56946 50559 57262 50560
rect 2606 50080 2922 50081
rect 2606 50016 2612 50080
rect 2676 50016 2692 50080
rect 2756 50016 2772 50080
rect 2836 50016 2852 50080
rect 2916 50016 2922 50080
rect 2606 50015 2922 50016
rect 7606 50080 7922 50081
rect 7606 50016 7612 50080
rect 7676 50016 7692 50080
rect 7756 50016 7772 50080
rect 7836 50016 7852 50080
rect 7916 50016 7922 50080
rect 7606 50015 7922 50016
rect 12606 50080 12922 50081
rect 12606 50016 12612 50080
rect 12676 50016 12692 50080
rect 12756 50016 12772 50080
rect 12836 50016 12852 50080
rect 12916 50016 12922 50080
rect 12606 50015 12922 50016
rect 17606 50080 17922 50081
rect 17606 50016 17612 50080
rect 17676 50016 17692 50080
rect 17756 50016 17772 50080
rect 17836 50016 17852 50080
rect 17916 50016 17922 50080
rect 17606 50015 17922 50016
rect 22606 50080 22922 50081
rect 22606 50016 22612 50080
rect 22676 50016 22692 50080
rect 22756 50016 22772 50080
rect 22836 50016 22852 50080
rect 22916 50016 22922 50080
rect 22606 50015 22922 50016
rect 27606 50080 27922 50081
rect 27606 50016 27612 50080
rect 27676 50016 27692 50080
rect 27756 50016 27772 50080
rect 27836 50016 27852 50080
rect 27916 50016 27922 50080
rect 27606 50015 27922 50016
rect 32606 50080 32922 50081
rect 32606 50016 32612 50080
rect 32676 50016 32692 50080
rect 32756 50016 32772 50080
rect 32836 50016 32852 50080
rect 32916 50016 32922 50080
rect 32606 50015 32922 50016
rect 37606 50080 37922 50081
rect 37606 50016 37612 50080
rect 37676 50016 37692 50080
rect 37756 50016 37772 50080
rect 37836 50016 37852 50080
rect 37916 50016 37922 50080
rect 37606 50015 37922 50016
rect 42606 50080 42922 50081
rect 42606 50016 42612 50080
rect 42676 50016 42692 50080
rect 42756 50016 42772 50080
rect 42836 50016 42852 50080
rect 42916 50016 42922 50080
rect 42606 50015 42922 50016
rect 47606 50080 47922 50081
rect 47606 50016 47612 50080
rect 47676 50016 47692 50080
rect 47756 50016 47772 50080
rect 47836 50016 47852 50080
rect 47916 50016 47922 50080
rect 47606 50015 47922 50016
rect 52606 50080 52922 50081
rect 52606 50016 52612 50080
rect 52676 50016 52692 50080
rect 52756 50016 52772 50080
rect 52836 50016 52852 50080
rect 52916 50016 52922 50080
rect 52606 50015 52922 50016
rect 57606 50080 57922 50081
rect 57606 50016 57612 50080
rect 57676 50016 57692 50080
rect 57756 50016 57772 50080
rect 57836 50016 57852 50080
rect 57916 50016 57922 50080
rect 57606 50015 57922 50016
rect 0 49784 800 49904
rect 58525 49874 58591 49877
rect 59200 49874 60000 49904
rect 58525 49872 60000 49874
rect 58525 49816 58530 49872
rect 58586 49816 60000 49872
rect 58525 49814 60000 49816
rect 58525 49811 58591 49814
rect 59200 49784 60000 49814
rect 1946 49536 2262 49537
rect 1946 49472 1952 49536
rect 2016 49472 2032 49536
rect 2096 49472 2112 49536
rect 2176 49472 2192 49536
rect 2256 49472 2262 49536
rect 1946 49471 2262 49472
rect 6946 49536 7262 49537
rect 6946 49472 6952 49536
rect 7016 49472 7032 49536
rect 7096 49472 7112 49536
rect 7176 49472 7192 49536
rect 7256 49472 7262 49536
rect 6946 49471 7262 49472
rect 11946 49536 12262 49537
rect 11946 49472 11952 49536
rect 12016 49472 12032 49536
rect 12096 49472 12112 49536
rect 12176 49472 12192 49536
rect 12256 49472 12262 49536
rect 11946 49471 12262 49472
rect 16946 49536 17262 49537
rect 16946 49472 16952 49536
rect 17016 49472 17032 49536
rect 17096 49472 17112 49536
rect 17176 49472 17192 49536
rect 17256 49472 17262 49536
rect 16946 49471 17262 49472
rect 21946 49536 22262 49537
rect 21946 49472 21952 49536
rect 22016 49472 22032 49536
rect 22096 49472 22112 49536
rect 22176 49472 22192 49536
rect 22256 49472 22262 49536
rect 21946 49471 22262 49472
rect 26946 49536 27262 49537
rect 26946 49472 26952 49536
rect 27016 49472 27032 49536
rect 27096 49472 27112 49536
rect 27176 49472 27192 49536
rect 27256 49472 27262 49536
rect 26946 49471 27262 49472
rect 31946 49536 32262 49537
rect 31946 49472 31952 49536
rect 32016 49472 32032 49536
rect 32096 49472 32112 49536
rect 32176 49472 32192 49536
rect 32256 49472 32262 49536
rect 31946 49471 32262 49472
rect 36946 49536 37262 49537
rect 36946 49472 36952 49536
rect 37016 49472 37032 49536
rect 37096 49472 37112 49536
rect 37176 49472 37192 49536
rect 37256 49472 37262 49536
rect 36946 49471 37262 49472
rect 41946 49536 42262 49537
rect 41946 49472 41952 49536
rect 42016 49472 42032 49536
rect 42096 49472 42112 49536
rect 42176 49472 42192 49536
rect 42256 49472 42262 49536
rect 41946 49471 42262 49472
rect 46946 49536 47262 49537
rect 46946 49472 46952 49536
rect 47016 49472 47032 49536
rect 47096 49472 47112 49536
rect 47176 49472 47192 49536
rect 47256 49472 47262 49536
rect 46946 49471 47262 49472
rect 51946 49536 52262 49537
rect 51946 49472 51952 49536
rect 52016 49472 52032 49536
rect 52096 49472 52112 49536
rect 52176 49472 52192 49536
rect 52256 49472 52262 49536
rect 51946 49471 52262 49472
rect 56946 49536 57262 49537
rect 56946 49472 56952 49536
rect 57016 49472 57032 49536
rect 57096 49472 57112 49536
rect 57176 49472 57192 49536
rect 57256 49472 57262 49536
rect 56946 49471 57262 49472
rect 58525 49058 58591 49061
rect 59200 49058 60000 49088
rect 58525 49056 60000 49058
rect 58525 49000 58530 49056
rect 58586 49000 60000 49056
rect 58525 48998 60000 49000
rect 58525 48995 58591 48998
rect 2606 48992 2922 48993
rect 2606 48928 2612 48992
rect 2676 48928 2692 48992
rect 2756 48928 2772 48992
rect 2836 48928 2852 48992
rect 2916 48928 2922 48992
rect 2606 48927 2922 48928
rect 7606 48992 7922 48993
rect 7606 48928 7612 48992
rect 7676 48928 7692 48992
rect 7756 48928 7772 48992
rect 7836 48928 7852 48992
rect 7916 48928 7922 48992
rect 7606 48927 7922 48928
rect 12606 48992 12922 48993
rect 12606 48928 12612 48992
rect 12676 48928 12692 48992
rect 12756 48928 12772 48992
rect 12836 48928 12852 48992
rect 12916 48928 12922 48992
rect 12606 48927 12922 48928
rect 17606 48992 17922 48993
rect 17606 48928 17612 48992
rect 17676 48928 17692 48992
rect 17756 48928 17772 48992
rect 17836 48928 17852 48992
rect 17916 48928 17922 48992
rect 17606 48927 17922 48928
rect 22606 48992 22922 48993
rect 22606 48928 22612 48992
rect 22676 48928 22692 48992
rect 22756 48928 22772 48992
rect 22836 48928 22852 48992
rect 22916 48928 22922 48992
rect 22606 48927 22922 48928
rect 27606 48992 27922 48993
rect 27606 48928 27612 48992
rect 27676 48928 27692 48992
rect 27756 48928 27772 48992
rect 27836 48928 27852 48992
rect 27916 48928 27922 48992
rect 27606 48927 27922 48928
rect 32606 48992 32922 48993
rect 32606 48928 32612 48992
rect 32676 48928 32692 48992
rect 32756 48928 32772 48992
rect 32836 48928 32852 48992
rect 32916 48928 32922 48992
rect 32606 48927 32922 48928
rect 37606 48992 37922 48993
rect 37606 48928 37612 48992
rect 37676 48928 37692 48992
rect 37756 48928 37772 48992
rect 37836 48928 37852 48992
rect 37916 48928 37922 48992
rect 37606 48927 37922 48928
rect 42606 48992 42922 48993
rect 42606 48928 42612 48992
rect 42676 48928 42692 48992
rect 42756 48928 42772 48992
rect 42836 48928 42852 48992
rect 42916 48928 42922 48992
rect 42606 48927 42922 48928
rect 47606 48992 47922 48993
rect 47606 48928 47612 48992
rect 47676 48928 47692 48992
rect 47756 48928 47772 48992
rect 47836 48928 47852 48992
rect 47916 48928 47922 48992
rect 47606 48927 47922 48928
rect 52606 48992 52922 48993
rect 52606 48928 52612 48992
rect 52676 48928 52692 48992
rect 52756 48928 52772 48992
rect 52836 48928 52852 48992
rect 52916 48928 52922 48992
rect 52606 48927 52922 48928
rect 57606 48992 57922 48993
rect 57606 48928 57612 48992
rect 57676 48928 57692 48992
rect 57756 48928 57772 48992
rect 57836 48928 57852 48992
rect 57916 48928 57922 48992
rect 59200 48968 60000 48998
rect 57606 48927 57922 48928
rect 1946 48448 2262 48449
rect 1946 48384 1952 48448
rect 2016 48384 2032 48448
rect 2096 48384 2112 48448
rect 2176 48384 2192 48448
rect 2256 48384 2262 48448
rect 1946 48383 2262 48384
rect 6946 48448 7262 48449
rect 6946 48384 6952 48448
rect 7016 48384 7032 48448
rect 7096 48384 7112 48448
rect 7176 48384 7192 48448
rect 7256 48384 7262 48448
rect 6946 48383 7262 48384
rect 11946 48448 12262 48449
rect 11946 48384 11952 48448
rect 12016 48384 12032 48448
rect 12096 48384 12112 48448
rect 12176 48384 12192 48448
rect 12256 48384 12262 48448
rect 11946 48383 12262 48384
rect 16946 48448 17262 48449
rect 16946 48384 16952 48448
rect 17016 48384 17032 48448
rect 17096 48384 17112 48448
rect 17176 48384 17192 48448
rect 17256 48384 17262 48448
rect 16946 48383 17262 48384
rect 21946 48448 22262 48449
rect 21946 48384 21952 48448
rect 22016 48384 22032 48448
rect 22096 48384 22112 48448
rect 22176 48384 22192 48448
rect 22256 48384 22262 48448
rect 21946 48383 22262 48384
rect 26946 48448 27262 48449
rect 26946 48384 26952 48448
rect 27016 48384 27032 48448
rect 27096 48384 27112 48448
rect 27176 48384 27192 48448
rect 27256 48384 27262 48448
rect 26946 48383 27262 48384
rect 31946 48448 32262 48449
rect 31946 48384 31952 48448
rect 32016 48384 32032 48448
rect 32096 48384 32112 48448
rect 32176 48384 32192 48448
rect 32256 48384 32262 48448
rect 31946 48383 32262 48384
rect 36946 48448 37262 48449
rect 36946 48384 36952 48448
rect 37016 48384 37032 48448
rect 37096 48384 37112 48448
rect 37176 48384 37192 48448
rect 37256 48384 37262 48448
rect 36946 48383 37262 48384
rect 41946 48448 42262 48449
rect 41946 48384 41952 48448
rect 42016 48384 42032 48448
rect 42096 48384 42112 48448
rect 42176 48384 42192 48448
rect 42256 48384 42262 48448
rect 41946 48383 42262 48384
rect 46946 48448 47262 48449
rect 46946 48384 46952 48448
rect 47016 48384 47032 48448
rect 47096 48384 47112 48448
rect 47176 48384 47192 48448
rect 47256 48384 47262 48448
rect 46946 48383 47262 48384
rect 51946 48448 52262 48449
rect 51946 48384 51952 48448
rect 52016 48384 52032 48448
rect 52096 48384 52112 48448
rect 52176 48384 52192 48448
rect 52256 48384 52262 48448
rect 51946 48383 52262 48384
rect 56946 48448 57262 48449
rect 56946 48384 56952 48448
rect 57016 48384 57032 48448
rect 57096 48384 57112 48448
rect 57176 48384 57192 48448
rect 57256 48384 57262 48448
rect 56946 48383 57262 48384
rect 58525 48242 58591 48245
rect 59200 48242 60000 48272
rect 58525 48240 60000 48242
rect 58525 48184 58530 48240
rect 58586 48184 60000 48240
rect 58525 48182 60000 48184
rect 58525 48179 58591 48182
rect 59200 48152 60000 48182
rect 2606 47904 2922 47905
rect 2606 47840 2612 47904
rect 2676 47840 2692 47904
rect 2756 47840 2772 47904
rect 2836 47840 2852 47904
rect 2916 47840 2922 47904
rect 2606 47839 2922 47840
rect 7606 47904 7922 47905
rect 7606 47840 7612 47904
rect 7676 47840 7692 47904
rect 7756 47840 7772 47904
rect 7836 47840 7852 47904
rect 7916 47840 7922 47904
rect 7606 47839 7922 47840
rect 12606 47904 12922 47905
rect 12606 47840 12612 47904
rect 12676 47840 12692 47904
rect 12756 47840 12772 47904
rect 12836 47840 12852 47904
rect 12916 47840 12922 47904
rect 12606 47839 12922 47840
rect 17606 47904 17922 47905
rect 17606 47840 17612 47904
rect 17676 47840 17692 47904
rect 17756 47840 17772 47904
rect 17836 47840 17852 47904
rect 17916 47840 17922 47904
rect 17606 47839 17922 47840
rect 22606 47904 22922 47905
rect 22606 47840 22612 47904
rect 22676 47840 22692 47904
rect 22756 47840 22772 47904
rect 22836 47840 22852 47904
rect 22916 47840 22922 47904
rect 22606 47839 22922 47840
rect 27606 47904 27922 47905
rect 27606 47840 27612 47904
rect 27676 47840 27692 47904
rect 27756 47840 27772 47904
rect 27836 47840 27852 47904
rect 27916 47840 27922 47904
rect 27606 47839 27922 47840
rect 32606 47904 32922 47905
rect 32606 47840 32612 47904
rect 32676 47840 32692 47904
rect 32756 47840 32772 47904
rect 32836 47840 32852 47904
rect 32916 47840 32922 47904
rect 32606 47839 32922 47840
rect 37606 47904 37922 47905
rect 37606 47840 37612 47904
rect 37676 47840 37692 47904
rect 37756 47840 37772 47904
rect 37836 47840 37852 47904
rect 37916 47840 37922 47904
rect 37606 47839 37922 47840
rect 42606 47904 42922 47905
rect 42606 47840 42612 47904
rect 42676 47840 42692 47904
rect 42756 47840 42772 47904
rect 42836 47840 42852 47904
rect 42916 47840 42922 47904
rect 42606 47839 42922 47840
rect 47606 47904 47922 47905
rect 47606 47840 47612 47904
rect 47676 47840 47692 47904
rect 47756 47840 47772 47904
rect 47836 47840 47852 47904
rect 47916 47840 47922 47904
rect 47606 47839 47922 47840
rect 52606 47904 52922 47905
rect 52606 47840 52612 47904
rect 52676 47840 52692 47904
rect 52756 47840 52772 47904
rect 52836 47840 52852 47904
rect 52916 47840 52922 47904
rect 52606 47839 52922 47840
rect 57606 47904 57922 47905
rect 57606 47840 57612 47904
rect 57676 47840 57692 47904
rect 57756 47840 57772 47904
rect 57836 47840 57852 47904
rect 57916 47840 57922 47904
rect 57606 47839 57922 47840
rect 58525 47426 58591 47429
rect 59200 47426 60000 47456
rect 58525 47424 60000 47426
rect 58525 47368 58530 47424
rect 58586 47368 60000 47424
rect 58525 47366 60000 47368
rect 58525 47363 58591 47366
rect 1946 47360 2262 47361
rect 1946 47296 1952 47360
rect 2016 47296 2032 47360
rect 2096 47296 2112 47360
rect 2176 47296 2192 47360
rect 2256 47296 2262 47360
rect 1946 47295 2262 47296
rect 6946 47360 7262 47361
rect 6946 47296 6952 47360
rect 7016 47296 7032 47360
rect 7096 47296 7112 47360
rect 7176 47296 7192 47360
rect 7256 47296 7262 47360
rect 6946 47295 7262 47296
rect 11946 47360 12262 47361
rect 11946 47296 11952 47360
rect 12016 47296 12032 47360
rect 12096 47296 12112 47360
rect 12176 47296 12192 47360
rect 12256 47296 12262 47360
rect 11946 47295 12262 47296
rect 16946 47360 17262 47361
rect 16946 47296 16952 47360
rect 17016 47296 17032 47360
rect 17096 47296 17112 47360
rect 17176 47296 17192 47360
rect 17256 47296 17262 47360
rect 16946 47295 17262 47296
rect 21946 47360 22262 47361
rect 21946 47296 21952 47360
rect 22016 47296 22032 47360
rect 22096 47296 22112 47360
rect 22176 47296 22192 47360
rect 22256 47296 22262 47360
rect 21946 47295 22262 47296
rect 26946 47360 27262 47361
rect 26946 47296 26952 47360
rect 27016 47296 27032 47360
rect 27096 47296 27112 47360
rect 27176 47296 27192 47360
rect 27256 47296 27262 47360
rect 26946 47295 27262 47296
rect 31946 47360 32262 47361
rect 31946 47296 31952 47360
rect 32016 47296 32032 47360
rect 32096 47296 32112 47360
rect 32176 47296 32192 47360
rect 32256 47296 32262 47360
rect 31946 47295 32262 47296
rect 36946 47360 37262 47361
rect 36946 47296 36952 47360
rect 37016 47296 37032 47360
rect 37096 47296 37112 47360
rect 37176 47296 37192 47360
rect 37256 47296 37262 47360
rect 36946 47295 37262 47296
rect 41946 47360 42262 47361
rect 41946 47296 41952 47360
rect 42016 47296 42032 47360
rect 42096 47296 42112 47360
rect 42176 47296 42192 47360
rect 42256 47296 42262 47360
rect 41946 47295 42262 47296
rect 46946 47360 47262 47361
rect 46946 47296 46952 47360
rect 47016 47296 47032 47360
rect 47096 47296 47112 47360
rect 47176 47296 47192 47360
rect 47256 47296 47262 47360
rect 46946 47295 47262 47296
rect 51946 47360 52262 47361
rect 51946 47296 51952 47360
rect 52016 47296 52032 47360
rect 52096 47296 52112 47360
rect 52176 47296 52192 47360
rect 52256 47296 52262 47360
rect 51946 47295 52262 47296
rect 56946 47360 57262 47361
rect 56946 47296 56952 47360
rect 57016 47296 57032 47360
rect 57096 47296 57112 47360
rect 57176 47296 57192 47360
rect 57256 47296 57262 47360
rect 59200 47336 60000 47366
rect 56946 47295 57262 47296
rect 2606 46816 2922 46817
rect 2606 46752 2612 46816
rect 2676 46752 2692 46816
rect 2756 46752 2772 46816
rect 2836 46752 2852 46816
rect 2916 46752 2922 46816
rect 2606 46751 2922 46752
rect 7606 46816 7922 46817
rect 7606 46752 7612 46816
rect 7676 46752 7692 46816
rect 7756 46752 7772 46816
rect 7836 46752 7852 46816
rect 7916 46752 7922 46816
rect 7606 46751 7922 46752
rect 12606 46816 12922 46817
rect 12606 46752 12612 46816
rect 12676 46752 12692 46816
rect 12756 46752 12772 46816
rect 12836 46752 12852 46816
rect 12916 46752 12922 46816
rect 12606 46751 12922 46752
rect 17606 46816 17922 46817
rect 17606 46752 17612 46816
rect 17676 46752 17692 46816
rect 17756 46752 17772 46816
rect 17836 46752 17852 46816
rect 17916 46752 17922 46816
rect 17606 46751 17922 46752
rect 22606 46816 22922 46817
rect 22606 46752 22612 46816
rect 22676 46752 22692 46816
rect 22756 46752 22772 46816
rect 22836 46752 22852 46816
rect 22916 46752 22922 46816
rect 22606 46751 22922 46752
rect 27606 46816 27922 46817
rect 27606 46752 27612 46816
rect 27676 46752 27692 46816
rect 27756 46752 27772 46816
rect 27836 46752 27852 46816
rect 27916 46752 27922 46816
rect 27606 46751 27922 46752
rect 32606 46816 32922 46817
rect 32606 46752 32612 46816
rect 32676 46752 32692 46816
rect 32756 46752 32772 46816
rect 32836 46752 32852 46816
rect 32916 46752 32922 46816
rect 32606 46751 32922 46752
rect 37606 46816 37922 46817
rect 37606 46752 37612 46816
rect 37676 46752 37692 46816
rect 37756 46752 37772 46816
rect 37836 46752 37852 46816
rect 37916 46752 37922 46816
rect 37606 46751 37922 46752
rect 42606 46816 42922 46817
rect 42606 46752 42612 46816
rect 42676 46752 42692 46816
rect 42756 46752 42772 46816
rect 42836 46752 42852 46816
rect 42916 46752 42922 46816
rect 42606 46751 42922 46752
rect 47606 46816 47922 46817
rect 47606 46752 47612 46816
rect 47676 46752 47692 46816
rect 47756 46752 47772 46816
rect 47836 46752 47852 46816
rect 47916 46752 47922 46816
rect 47606 46751 47922 46752
rect 52606 46816 52922 46817
rect 52606 46752 52612 46816
rect 52676 46752 52692 46816
rect 52756 46752 52772 46816
rect 52836 46752 52852 46816
rect 52916 46752 52922 46816
rect 52606 46751 52922 46752
rect 57606 46816 57922 46817
rect 57606 46752 57612 46816
rect 57676 46752 57692 46816
rect 57756 46752 57772 46816
rect 57836 46752 57852 46816
rect 57916 46752 57922 46816
rect 57606 46751 57922 46752
rect 58525 46610 58591 46613
rect 59200 46610 60000 46640
rect 58525 46608 60000 46610
rect 58525 46552 58530 46608
rect 58586 46552 60000 46608
rect 58525 46550 60000 46552
rect 58525 46547 58591 46550
rect 59200 46520 60000 46550
rect 1946 46272 2262 46273
rect 1946 46208 1952 46272
rect 2016 46208 2032 46272
rect 2096 46208 2112 46272
rect 2176 46208 2192 46272
rect 2256 46208 2262 46272
rect 1946 46207 2262 46208
rect 6946 46272 7262 46273
rect 6946 46208 6952 46272
rect 7016 46208 7032 46272
rect 7096 46208 7112 46272
rect 7176 46208 7192 46272
rect 7256 46208 7262 46272
rect 6946 46207 7262 46208
rect 11946 46272 12262 46273
rect 11946 46208 11952 46272
rect 12016 46208 12032 46272
rect 12096 46208 12112 46272
rect 12176 46208 12192 46272
rect 12256 46208 12262 46272
rect 11946 46207 12262 46208
rect 16946 46272 17262 46273
rect 16946 46208 16952 46272
rect 17016 46208 17032 46272
rect 17096 46208 17112 46272
rect 17176 46208 17192 46272
rect 17256 46208 17262 46272
rect 16946 46207 17262 46208
rect 21946 46272 22262 46273
rect 21946 46208 21952 46272
rect 22016 46208 22032 46272
rect 22096 46208 22112 46272
rect 22176 46208 22192 46272
rect 22256 46208 22262 46272
rect 21946 46207 22262 46208
rect 26946 46272 27262 46273
rect 26946 46208 26952 46272
rect 27016 46208 27032 46272
rect 27096 46208 27112 46272
rect 27176 46208 27192 46272
rect 27256 46208 27262 46272
rect 26946 46207 27262 46208
rect 31946 46272 32262 46273
rect 31946 46208 31952 46272
rect 32016 46208 32032 46272
rect 32096 46208 32112 46272
rect 32176 46208 32192 46272
rect 32256 46208 32262 46272
rect 31946 46207 32262 46208
rect 36946 46272 37262 46273
rect 36946 46208 36952 46272
rect 37016 46208 37032 46272
rect 37096 46208 37112 46272
rect 37176 46208 37192 46272
rect 37256 46208 37262 46272
rect 36946 46207 37262 46208
rect 41946 46272 42262 46273
rect 41946 46208 41952 46272
rect 42016 46208 42032 46272
rect 42096 46208 42112 46272
rect 42176 46208 42192 46272
rect 42256 46208 42262 46272
rect 41946 46207 42262 46208
rect 46946 46272 47262 46273
rect 46946 46208 46952 46272
rect 47016 46208 47032 46272
rect 47096 46208 47112 46272
rect 47176 46208 47192 46272
rect 47256 46208 47262 46272
rect 46946 46207 47262 46208
rect 51946 46272 52262 46273
rect 51946 46208 51952 46272
rect 52016 46208 52032 46272
rect 52096 46208 52112 46272
rect 52176 46208 52192 46272
rect 52256 46208 52262 46272
rect 51946 46207 52262 46208
rect 56946 46272 57262 46273
rect 56946 46208 56952 46272
rect 57016 46208 57032 46272
rect 57096 46208 57112 46272
rect 57176 46208 57192 46272
rect 57256 46208 57262 46272
rect 56946 46207 57262 46208
rect 58525 45794 58591 45797
rect 59200 45794 60000 45824
rect 58525 45792 60000 45794
rect 58525 45736 58530 45792
rect 58586 45736 60000 45792
rect 58525 45734 60000 45736
rect 58525 45731 58591 45734
rect 2606 45728 2922 45729
rect 2606 45664 2612 45728
rect 2676 45664 2692 45728
rect 2756 45664 2772 45728
rect 2836 45664 2852 45728
rect 2916 45664 2922 45728
rect 2606 45663 2922 45664
rect 7606 45728 7922 45729
rect 7606 45664 7612 45728
rect 7676 45664 7692 45728
rect 7756 45664 7772 45728
rect 7836 45664 7852 45728
rect 7916 45664 7922 45728
rect 7606 45663 7922 45664
rect 12606 45728 12922 45729
rect 12606 45664 12612 45728
rect 12676 45664 12692 45728
rect 12756 45664 12772 45728
rect 12836 45664 12852 45728
rect 12916 45664 12922 45728
rect 12606 45663 12922 45664
rect 17606 45728 17922 45729
rect 17606 45664 17612 45728
rect 17676 45664 17692 45728
rect 17756 45664 17772 45728
rect 17836 45664 17852 45728
rect 17916 45664 17922 45728
rect 17606 45663 17922 45664
rect 22606 45728 22922 45729
rect 22606 45664 22612 45728
rect 22676 45664 22692 45728
rect 22756 45664 22772 45728
rect 22836 45664 22852 45728
rect 22916 45664 22922 45728
rect 22606 45663 22922 45664
rect 27606 45728 27922 45729
rect 27606 45664 27612 45728
rect 27676 45664 27692 45728
rect 27756 45664 27772 45728
rect 27836 45664 27852 45728
rect 27916 45664 27922 45728
rect 27606 45663 27922 45664
rect 32606 45728 32922 45729
rect 32606 45664 32612 45728
rect 32676 45664 32692 45728
rect 32756 45664 32772 45728
rect 32836 45664 32852 45728
rect 32916 45664 32922 45728
rect 32606 45663 32922 45664
rect 37606 45728 37922 45729
rect 37606 45664 37612 45728
rect 37676 45664 37692 45728
rect 37756 45664 37772 45728
rect 37836 45664 37852 45728
rect 37916 45664 37922 45728
rect 37606 45663 37922 45664
rect 42606 45728 42922 45729
rect 42606 45664 42612 45728
rect 42676 45664 42692 45728
rect 42756 45664 42772 45728
rect 42836 45664 42852 45728
rect 42916 45664 42922 45728
rect 42606 45663 42922 45664
rect 47606 45728 47922 45729
rect 47606 45664 47612 45728
rect 47676 45664 47692 45728
rect 47756 45664 47772 45728
rect 47836 45664 47852 45728
rect 47916 45664 47922 45728
rect 47606 45663 47922 45664
rect 52606 45728 52922 45729
rect 52606 45664 52612 45728
rect 52676 45664 52692 45728
rect 52756 45664 52772 45728
rect 52836 45664 52852 45728
rect 52916 45664 52922 45728
rect 52606 45663 52922 45664
rect 57606 45728 57922 45729
rect 57606 45664 57612 45728
rect 57676 45664 57692 45728
rect 57756 45664 57772 45728
rect 57836 45664 57852 45728
rect 57916 45664 57922 45728
rect 59200 45704 60000 45734
rect 57606 45663 57922 45664
rect 1946 45184 2262 45185
rect 1946 45120 1952 45184
rect 2016 45120 2032 45184
rect 2096 45120 2112 45184
rect 2176 45120 2192 45184
rect 2256 45120 2262 45184
rect 1946 45119 2262 45120
rect 6946 45184 7262 45185
rect 6946 45120 6952 45184
rect 7016 45120 7032 45184
rect 7096 45120 7112 45184
rect 7176 45120 7192 45184
rect 7256 45120 7262 45184
rect 6946 45119 7262 45120
rect 11946 45184 12262 45185
rect 11946 45120 11952 45184
rect 12016 45120 12032 45184
rect 12096 45120 12112 45184
rect 12176 45120 12192 45184
rect 12256 45120 12262 45184
rect 11946 45119 12262 45120
rect 16946 45184 17262 45185
rect 16946 45120 16952 45184
rect 17016 45120 17032 45184
rect 17096 45120 17112 45184
rect 17176 45120 17192 45184
rect 17256 45120 17262 45184
rect 16946 45119 17262 45120
rect 21946 45184 22262 45185
rect 21946 45120 21952 45184
rect 22016 45120 22032 45184
rect 22096 45120 22112 45184
rect 22176 45120 22192 45184
rect 22256 45120 22262 45184
rect 21946 45119 22262 45120
rect 26946 45184 27262 45185
rect 26946 45120 26952 45184
rect 27016 45120 27032 45184
rect 27096 45120 27112 45184
rect 27176 45120 27192 45184
rect 27256 45120 27262 45184
rect 26946 45119 27262 45120
rect 31946 45184 32262 45185
rect 31946 45120 31952 45184
rect 32016 45120 32032 45184
rect 32096 45120 32112 45184
rect 32176 45120 32192 45184
rect 32256 45120 32262 45184
rect 31946 45119 32262 45120
rect 36946 45184 37262 45185
rect 36946 45120 36952 45184
rect 37016 45120 37032 45184
rect 37096 45120 37112 45184
rect 37176 45120 37192 45184
rect 37256 45120 37262 45184
rect 36946 45119 37262 45120
rect 41946 45184 42262 45185
rect 41946 45120 41952 45184
rect 42016 45120 42032 45184
rect 42096 45120 42112 45184
rect 42176 45120 42192 45184
rect 42256 45120 42262 45184
rect 41946 45119 42262 45120
rect 46946 45184 47262 45185
rect 46946 45120 46952 45184
rect 47016 45120 47032 45184
rect 47096 45120 47112 45184
rect 47176 45120 47192 45184
rect 47256 45120 47262 45184
rect 46946 45119 47262 45120
rect 51946 45184 52262 45185
rect 51946 45120 51952 45184
rect 52016 45120 52032 45184
rect 52096 45120 52112 45184
rect 52176 45120 52192 45184
rect 52256 45120 52262 45184
rect 51946 45119 52262 45120
rect 56946 45184 57262 45185
rect 56946 45120 56952 45184
rect 57016 45120 57032 45184
rect 57096 45120 57112 45184
rect 57176 45120 57192 45184
rect 57256 45120 57262 45184
rect 56946 45119 57262 45120
rect 58525 44978 58591 44981
rect 59200 44978 60000 45008
rect 58525 44976 60000 44978
rect 58525 44920 58530 44976
rect 58586 44920 60000 44976
rect 58525 44918 60000 44920
rect 58525 44915 58591 44918
rect 59200 44888 60000 44918
rect 2606 44640 2922 44641
rect 2606 44576 2612 44640
rect 2676 44576 2692 44640
rect 2756 44576 2772 44640
rect 2836 44576 2852 44640
rect 2916 44576 2922 44640
rect 2606 44575 2922 44576
rect 7606 44640 7922 44641
rect 7606 44576 7612 44640
rect 7676 44576 7692 44640
rect 7756 44576 7772 44640
rect 7836 44576 7852 44640
rect 7916 44576 7922 44640
rect 7606 44575 7922 44576
rect 12606 44640 12922 44641
rect 12606 44576 12612 44640
rect 12676 44576 12692 44640
rect 12756 44576 12772 44640
rect 12836 44576 12852 44640
rect 12916 44576 12922 44640
rect 12606 44575 12922 44576
rect 17606 44640 17922 44641
rect 17606 44576 17612 44640
rect 17676 44576 17692 44640
rect 17756 44576 17772 44640
rect 17836 44576 17852 44640
rect 17916 44576 17922 44640
rect 17606 44575 17922 44576
rect 22606 44640 22922 44641
rect 22606 44576 22612 44640
rect 22676 44576 22692 44640
rect 22756 44576 22772 44640
rect 22836 44576 22852 44640
rect 22916 44576 22922 44640
rect 22606 44575 22922 44576
rect 27606 44640 27922 44641
rect 27606 44576 27612 44640
rect 27676 44576 27692 44640
rect 27756 44576 27772 44640
rect 27836 44576 27852 44640
rect 27916 44576 27922 44640
rect 27606 44575 27922 44576
rect 32606 44640 32922 44641
rect 32606 44576 32612 44640
rect 32676 44576 32692 44640
rect 32756 44576 32772 44640
rect 32836 44576 32852 44640
rect 32916 44576 32922 44640
rect 32606 44575 32922 44576
rect 37606 44640 37922 44641
rect 37606 44576 37612 44640
rect 37676 44576 37692 44640
rect 37756 44576 37772 44640
rect 37836 44576 37852 44640
rect 37916 44576 37922 44640
rect 37606 44575 37922 44576
rect 42606 44640 42922 44641
rect 42606 44576 42612 44640
rect 42676 44576 42692 44640
rect 42756 44576 42772 44640
rect 42836 44576 42852 44640
rect 42916 44576 42922 44640
rect 42606 44575 42922 44576
rect 47606 44640 47922 44641
rect 47606 44576 47612 44640
rect 47676 44576 47692 44640
rect 47756 44576 47772 44640
rect 47836 44576 47852 44640
rect 47916 44576 47922 44640
rect 47606 44575 47922 44576
rect 52606 44640 52922 44641
rect 52606 44576 52612 44640
rect 52676 44576 52692 44640
rect 52756 44576 52772 44640
rect 52836 44576 52852 44640
rect 52916 44576 52922 44640
rect 52606 44575 52922 44576
rect 57606 44640 57922 44641
rect 57606 44576 57612 44640
rect 57676 44576 57692 44640
rect 57756 44576 57772 44640
rect 57836 44576 57852 44640
rect 57916 44576 57922 44640
rect 57606 44575 57922 44576
rect 58525 44162 58591 44165
rect 59200 44162 60000 44192
rect 58525 44160 60000 44162
rect 58525 44104 58530 44160
rect 58586 44104 60000 44160
rect 58525 44102 60000 44104
rect 58525 44099 58591 44102
rect 1946 44096 2262 44097
rect 1946 44032 1952 44096
rect 2016 44032 2032 44096
rect 2096 44032 2112 44096
rect 2176 44032 2192 44096
rect 2256 44032 2262 44096
rect 1946 44031 2262 44032
rect 6946 44096 7262 44097
rect 6946 44032 6952 44096
rect 7016 44032 7032 44096
rect 7096 44032 7112 44096
rect 7176 44032 7192 44096
rect 7256 44032 7262 44096
rect 6946 44031 7262 44032
rect 11946 44096 12262 44097
rect 11946 44032 11952 44096
rect 12016 44032 12032 44096
rect 12096 44032 12112 44096
rect 12176 44032 12192 44096
rect 12256 44032 12262 44096
rect 11946 44031 12262 44032
rect 16946 44096 17262 44097
rect 16946 44032 16952 44096
rect 17016 44032 17032 44096
rect 17096 44032 17112 44096
rect 17176 44032 17192 44096
rect 17256 44032 17262 44096
rect 16946 44031 17262 44032
rect 21946 44096 22262 44097
rect 21946 44032 21952 44096
rect 22016 44032 22032 44096
rect 22096 44032 22112 44096
rect 22176 44032 22192 44096
rect 22256 44032 22262 44096
rect 21946 44031 22262 44032
rect 26946 44096 27262 44097
rect 26946 44032 26952 44096
rect 27016 44032 27032 44096
rect 27096 44032 27112 44096
rect 27176 44032 27192 44096
rect 27256 44032 27262 44096
rect 26946 44031 27262 44032
rect 31946 44096 32262 44097
rect 31946 44032 31952 44096
rect 32016 44032 32032 44096
rect 32096 44032 32112 44096
rect 32176 44032 32192 44096
rect 32256 44032 32262 44096
rect 31946 44031 32262 44032
rect 36946 44096 37262 44097
rect 36946 44032 36952 44096
rect 37016 44032 37032 44096
rect 37096 44032 37112 44096
rect 37176 44032 37192 44096
rect 37256 44032 37262 44096
rect 36946 44031 37262 44032
rect 41946 44096 42262 44097
rect 41946 44032 41952 44096
rect 42016 44032 42032 44096
rect 42096 44032 42112 44096
rect 42176 44032 42192 44096
rect 42256 44032 42262 44096
rect 41946 44031 42262 44032
rect 46946 44096 47262 44097
rect 46946 44032 46952 44096
rect 47016 44032 47032 44096
rect 47096 44032 47112 44096
rect 47176 44032 47192 44096
rect 47256 44032 47262 44096
rect 46946 44031 47262 44032
rect 51946 44096 52262 44097
rect 51946 44032 51952 44096
rect 52016 44032 52032 44096
rect 52096 44032 52112 44096
rect 52176 44032 52192 44096
rect 52256 44032 52262 44096
rect 51946 44031 52262 44032
rect 56946 44096 57262 44097
rect 56946 44032 56952 44096
rect 57016 44032 57032 44096
rect 57096 44032 57112 44096
rect 57176 44032 57192 44096
rect 57256 44032 57262 44096
rect 59200 44072 60000 44102
rect 56946 44031 57262 44032
rect 2606 43552 2922 43553
rect 2606 43488 2612 43552
rect 2676 43488 2692 43552
rect 2756 43488 2772 43552
rect 2836 43488 2852 43552
rect 2916 43488 2922 43552
rect 2606 43487 2922 43488
rect 7606 43552 7922 43553
rect 7606 43488 7612 43552
rect 7676 43488 7692 43552
rect 7756 43488 7772 43552
rect 7836 43488 7852 43552
rect 7916 43488 7922 43552
rect 7606 43487 7922 43488
rect 12606 43552 12922 43553
rect 12606 43488 12612 43552
rect 12676 43488 12692 43552
rect 12756 43488 12772 43552
rect 12836 43488 12852 43552
rect 12916 43488 12922 43552
rect 12606 43487 12922 43488
rect 17606 43552 17922 43553
rect 17606 43488 17612 43552
rect 17676 43488 17692 43552
rect 17756 43488 17772 43552
rect 17836 43488 17852 43552
rect 17916 43488 17922 43552
rect 17606 43487 17922 43488
rect 22606 43552 22922 43553
rect 22606 43488 22612 43552
rect 22676 43488 22692 43552
rect 22756 43488 22772 43552
rect 22836 43488 22852 43552
rect 22916 43488 22922 43552
rect 22606 43487 22922 43488
rect 27606 43552 27922 43553
rect 27606 43488 27612 43552
rect 27676 43488 27692 43552
rect 27756 43488 27772 43552
rect 27836 43488 27852 43552
rect 27916 43488 27922 43552
rect 27606 43487 27922 43488
rect 32606 43552 32922 43553
rect 32606 43488 32612 43552
rect 32676 43488 32692 43552
rect 32756 43488 32772 43552
rect 32836 43488 32852 43552
rect 32916 43488 32922 43552
rect 32606 43487 32922 43488
rect 37606 43552 37922 43553
rect 37606 43488 37612 43552
rect 37676 43488 37692 43552
rect 37756 43488 37772 43552
rect 37836 43488 37852 43552
rect 37916 43488 37922 43552
rect 37606 43487 37922 43488
rect 42606 43552 42922 43553
rect 42606 43488 42612 43552
rect 42676 43488 42692 43552
rect 42756 43488 42772 43552
rect 42836 43488 42852 43552
rect 42916 43488 42922 43552
rect 42606 43487 42922 43488
rect 47606 43552 47922 43553
rect 47606 43488 47612 43552
rect 47676 43488 47692 43552
rect 47756 43488 47772 43552
rect 47836 43488 47852 43552
rect 47916 43488 47922 43552
rect 47606 43487 47922 43488
rect 52606 43552 52922 43553
rect 52606 43488 52612 43552
rect 52676 43488 52692 43552
rect 52756 43488 52772 43552
rect 52836 43488 52852 43552
rect 52916 43488 52922 43552
rect 52606 43487 52922 43488
rect 57606 43552 57922 43553
rect 57606 43488 57612 43552
rect 57676 43488 57692 43552
rect 57756 43488 57772 43552
rect 57836 43488 57852 43552
rect 57916 43488 57922 43552
rect 57606 43487 57922 43488
rect 58525 43346 58591 43349
rect 59200 43346 60000 43376
rect 58525 43344 60000 43346
rect 58525 43288 58530 43344
rect 58586 43288 60000 43344
rect 58525 43286 60000 43288
rect 58525 43283 58591 43286
rect 59200 43256 60000 43286
rect 1946 43008 2262 43009
rect 1946 42944 1952 43008
rect 2016 42944 2032 43008
rect 2096 42944 2112 43008
rect 2176 42944 2192 43008
rect 2256 42944 2262 43008
rect 1946 42943 2262 42944
rect 6946 43008 7262 43009
rect 6946 42944 6952 43008
rect 7016 42944 7032 43008
rect 7096 42944 7112 43008
rect 7176 42944 7192 43008
rect 7256 42944 7262 43008
rect 6946 42943 7262 42944
rect 11946 43008 12262 43009
rect 11946 42944 11952 43008
rect 12016 42944 12032 43008
rect 12096 42944 12112 43008
rect 12176 42944 12192 43008
rect 12256 42944 12262 43008
rect 11946 42943 12262 42944
rect 16946 43008 17262 43009
rect 16946 42944 16952 43008
rect 17016 42944 17032 43008
rect 17096 42944 17112 43008
rect 17176 42944 17192 43008
rect 17256 42944 17262 43008
rect 16946 42943 17262 42944
rect 21946 43008 22262 43009
rect 21946 42944 21952 43008
rect 22016 42944 22032 43008
rect 22096 42944 22112 43008
rect 22176 42944 22192 43008
rect 22256 42944 22262 43008
rect 21946 42943 22262 42944
rect 26946 43008 27262 43009
rect 26946 42944 26952 43008
rect 27016 42944 27032 43008
rect 27096 42944 27112 43008
rect 27176 42944 27192 43008
rect 27256 42944 27262 43008
rect 26946 42943 27262 42944
rect 31946 43008 32262 43009
rect 31946 42944 31952 43008
rect 32016 42944 32032 43008
rect 32096 42944 32112 43008
rect 32176 42944 32192 43008
rect 32256 42944 32262 43008
rect 31946 42943 32262 42944
rect 36946 43008 37262 43009
rect 36946 42944 36952 43008
rect 37016 42944 37032 43008
rect 37096 42944 37112 43008
rect 37176 42944 37192 43008
rect 37256 42944 37262 43008
rect 36946 42943 37262 42944
rect 41946 43008 42262 43009
rect 41946 42944 41952 43008
rect 42016 42944 42032 43008
rect 42096 42944 42112 43008
rect 42176 42944 42192 43008
rect 42256 42944 42262 43008
rect 41946 42943 42262 42944
rect 46946 43008 47262 43009
rect 46946 42944 46952 43008
rect 47016 42944 47032 43008
rect 47096 42944 47112 43008
rect 47176 42944 47192 43008
rect 47256 42944 47262 43008
rect 46946 42943 47262 42944
rect 51946 43008 52262 43009
rect 51946 42944 51952 43008
rect 52016 42944 52032 43008
rect 52096 42944 52112 43008
rect 52176 42944 52192 43008
rect 52256 42944 52262 43008
rect 51946 42943 52262 42944
rect 56946 43008 57262 43009
rect 56946 42944 56952 43008
rect 57016 42944 57032 43008
rect 57096 42944 57112 43008
rect 57176 42944 57192 43008
rect 57256 42944 57262 43008
rect 56946 42943 57262 42944
rect 58525 42530 58591 42533
rect 59200 42530 60000 42560
rect 58525 42528 60000 42530
rect 58525 42472 58530 42528
rect 58586 42472 60000 42528
rect 58525 42470 60000 42472
rect 58525 42467 58591 42470
rect 2606 42464 2922 42465
rect 2606 42400 2612 42464
rect 2676 42400 2692 42464
rect 2756 42400 2772 42464
rect 2836 42400 2852 42464
rect 2916 42400 2922 42464
rect 2606 42399 2922 42400
rect 7606 42464 7922 42465
rect 7606 42400 7612 42464
rect 7676 42400 7692 42464
rect 7756 42400 7772 42464
rect 7836 42400 7852 42464
rect 7916 42400 7922 42464
rect 7606 42399 7922 42400
rect 12606 42464 12922 42465
rect 12606 42400 12612 42464
rect 12676 42400 12692 42464
rect 12756 42400 12772 42464
rect 12836 42400 12852 42464
rect 12916 42400 12922 42464
rect 12606 42399 12922 42400
rect 17606 42464 17922 42465
rect 17606 42400 17612 42464
rect 17676 42400 17692 42464
rect 17756 42400 17772 42464
rect 17836 42400 17852 42464
rect 17916 42400 17922 42464
rect 17606 42399 17922 42400
rect 22606 42464 22922 42465
rect 22606 42400 22612 42464
rect 22676 42400 22692 42464
rect 22756 42400 22772 42464
rect 22836 42400 22852 42464
rect 22916 42400 22922 42464
rect 22606 42399 22922 42400
rect 27606 42464 27922 42465
rect 27606 42400 27612 42464
rect 27676 42400 27692 42464
rect 27756 42400 27772 42464
rect 27836 42400 27852 42464
rect 27916 42400 27922 42464
rect 27606 42399 27922 42400
rect 32606 42464 32922 42465
rect 32606 42400 32612 42464
rect 32676 42400 32692 42464
rect 32756 42400 32772 42464
rect 32836 42400 32852 42464
rect 32916 42400 32922 42464
rect 32606 42399 32922 42400
rect 37606 42464 37922 42465
rect 37606 42400 37612 42464
rect 37676 42400 37692 42464
rect 37756 42400 37772 42464
rect 37836 42400 37852 42464
rect 37916 42400 37922 42464
rect 37606 42399 37922 42400
rect 42606 42464 42922 42465
rect 42606 42400 42612 42464
rect 42676 42400 42692 42464
rect 42756 42400 42772 42464
rect 42836 42400 42852 42464
rect 42916 42400 42922 42464
rect 42606 42399 42922 42400
rect 47606 42464 47922 42465
rect 47606 42400 47612 42464
rect 47676 42400 47692 42464
rect 47756 42400 47772 42464
rect 47836 42400 47852 42464
rect 47916 42400 47922 42464
rect 47606 42399 47922 42400
rect 52606 42464 52922 42465
rect 52606 42400 52612 42464
rect 52676 42400 52692 42464
rect 52756 42400 52772 42464
rect 52836 42400 52852 42464
rect 52916 42400 52922 42464
rect 52606 42399 52922 42400
rect 57606 42464 57922 42465
rect 57606 42400 57612 42464
rect 57676 42400 57692 42464
rect 57756 42400 57772 42464
rect 57836 42400 57852 42464
rect 57916 42400 57922 42464
rect 59200 42440 60000 42470
rect 57606 42399 57922 42400
rect 1946 41920 2262 41921
rect 1946 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2262 41920
rect 1946 41855 2262 41856
rect 6946 41920 7262 41921
rect 6946 41856 6952 41920
rect 7016 41856 7032 41920
rect 7096 41856 7112 41920
rect 7176 41856 7192 41920
rect 7256 41856 7262 41920
rect 6946 41855 7262 41856
rect 11946 41920 12262 41921
rect 11946 41856 11952 41920
rect 12016 41856 12032 41920
rect 12096 41856 12112 41920
rect 12176 41856 12192 41920
rect 12256 41856 12262 41920
rect 11946 41855 12262 41856
rect 16946 41920 17262 41921
rect 16946 41856 16952 41920
rect 17016 41856 17032 41920
rect 17096 41856 17112 41920
rect 17176 41856 17192 41920
rect 17256 41856 17262 41920
rect 16946 41855 17262 41856
rect 21946 41920 22262 41921
rect 21946 41856 21952 41920
rect 22016 41856 22032 41920
rect 22096 41856 22112 41920
rect 22176 41856 22192 41920
rect 22256 41856 22262 41920
rect 21946 41855 22262 41856
rect 26946 41920 27262 41921
rect 26946 41856 26952 41920
rect 27016 41856 27032 41920
rect 27096 41856 27112 41920
rect 27176 41856 27192 41920
rect 27256 41856 27262 41920
rect 26946 41855 27262 41856
rect 31946 41920 32262 41921
rect 31946 41856 31952 41920
rect 32016 41856 32032 41920
rect 32096 41856 32112 41920
rect 32176 41856 32192 41920
rect 32256 41856 32262 41920
rect 31946 41855 32262 41856
rect 36946 41920 37262 41921
rect 36946 41856 36952 41920
rect 37016 41856 37032 41920
rect 37096 41856 37112 41920
rect 37176 41856 37192 41920
rect 37256 41856 37262 41920
rect 36946 41855 37262 41856
rect 41946 41920 42262 41921
rect 41946 41856 41952 41920
rect 42016 41856 42032 41920
rect 42096 41856 42112 41920
rect 42176 41856 42192 41920
rect 42256 41856 42262 41920
rect 41946 41855 42262 41856
rect 46946 41920 47262 41921
rect 46946 41856 46952 41920
rect 47016 41856 47032 41920
rect 47096 41856 47112 41920
rect 47176 41856 47192 41920
rect 47256 41856 47262 41920
rect 46946 41855 47262 41856
rect 51946 41920 52262 41921
rect 51946 41856 51952 41920
rect 52016 41856 52032 41920
rect 52096 41856 52112 41920
rect 52176 41856 52192 41920
rect 52256 41856 52262 41920
rect 51946 41855 52262 41856
rect 56946 41920 57262 41921
rect 56946 41856 56952 41920
rect 57016 41856 57032 41920
rect 57096 41856 57112 41920
rect 57176 41856 57192 41920
rect 57256 41856 57262 41920
rect 56946 41855 57262 41856
rect 58525 41714 58591 41717
rect 59200 41714 60000 41744
rect 58525 41712 60000 41714
rect 58525 41656 58530 41712
rect 58586 41656 60000 41712
rect 58525 41654 60000 41656
rect 58525 41651 58591 41654
rect 59200 41624 60000 41654
rect 2606 41376 2922 41377
rect 2606 41312 2612 41376
rect 2676 41312 2692 41376
rect 2756 41312 2772 41376
rect 2836 41312 2852 41376
rect 2916 41312 2922 41376
rect 2606 41311 2922 41312
rect 7606 41376 7922 41377
rect 7606 41312 7612 41376
rect 7676 41312 7692 41376
rect 7756 41312 7772 41376
rect 7836 41312 7852 41376
rect 7916 41312 7922 41376
rect 7606 41311 7922 41312
rect 12606 41376 12922 41377
rect 12606 41312 12612 41376
rect 12676 41312 12692 41376
rect 12756 41312 12772 41376
rect 12836 41312 12852 41376
rect 12916 41312 12922 41376
rect 12606 41311 12922 41312
rect 17606 41376 17922 41377
rect 17606 41312 17612 41376
rect 17676 41312 17692 41376
rect 17756 41312 17772 41376
rect 17836 41312 17852 41376
rect 17916 41312 17922 41376
rect 17606 41311 17922 41312
rect 22606 41376 22922 41377
rect 22606 41312 22612 41376
rect 22676 41312 22692 41376
rect 22756 41312 22772 41376
rect 22836 41312 22852 41376
rect 22916 41312 22922 41376
rect 22606 41311 22922 41312
rect 27606 41376 27922 41377
rect 27606 41312 27612 41376
rect 27676 41312 27692 41376
rect 27756 41312 27772 41376
rect 27836 41312 27852 41376
rect 27916 41312 27922 41376
rect 27606 41311 27922 41312
rect 32606 41376 32922 41377
rect 32606 41312 32612 41376
rect 32676 41312 32692 41376
rect 32756 41312 32772 41376
rect 32836 41312 32852 41376
rect 32916 41312 32922 41376
rect 32606 41311 32922 41312
rect 37606 41376 37922 41377
rect 37606 41312 37612 41376
rect 37676 41312 37692 41376
rect 37756 41312 37772 41376
rect 37836 41312 37852 41376
rect 37916 41312 37922 41376
rect 37606 41311 37922 41312
rect 42606 41376 42922 41377
rect 42606 41312 42612 41376
rect 42676 41312 42692 41376
rect 42756 41312 42772 41376
rect 42836 41312 42852 41376
rect 42916 41312 42922 41376
rect 42606 41311 42922 41312
rect 47606 41376 47922 41377
rect 47606 41312 47612 41376
rect 47676 41312 47692 41376
rect 47756 41312 47772 41376
rect 47836 41312 47852 41376
rect 47916 41312 47922 41376
rect 47606 41311 47922 41312
rect 52606 41376 52922 41377
rect 52606 41312 52612 41376
rect 52676 41312 52692 41376
rect 52756 41312 52772 41376
rect 52836 41312 52852 41376
rect 52916 41312 52922 41376
rect 52606 41311 52922 41312
rect 57606 41376 57922 41377
rect 57606 41312 57612 41376
rect 57676 41312 57692 41376
rect 57756 41312 57772 41376
rect 57836 41312 57852 41376
rect 57916 41312 57922 41376
rect 57606 41311 57922 41312
rect 58525 40898 58591 40901
rect 59200 40898 60000 40928
rect 58525 40896 60000 40898
rect 58525 40840 58530 40896
rect 58586 40840 60000 40896
rect 58525 40838 60000 40840
rect 58525 40835 58591 40838
rect 1946 40832 2262 40833
rect 1946 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2262 40832
rect 1946 40767 2262 40768
rect 6946 40832 7262 40833
rect 6946 40768 6952 40832
rect 7016 40768 7032 40832
rect 7096 40768 7112 40832
rect 7176 40768 7192 40832
rect 7256 40768 7262 40832
rect 6946 40767 7262 40768
rect 11946 40832 12262 40833
rect 11946 40768 11952 40832
rect 12016 40768 12032 40832
rect 12096 40768 12112 40832
rect 12176 40768 12192 40832
rect 12256 40768 12262 40832
rect 11946 40767 12262 40768
rect 16946 40832 17262 40833
rect 16946 40768 16952 40832
rect 17016 40768 17032 40832
rect 17096 40768 17112 40832
rect 17176 40768 17192 40832
rect 17256 40768 17262 40832
rect 16946 40767 17262 40768
rect 21946 40832 22262 40833
rect 21946 40768 21952 40832
rect 22016 40768 22032 40832
rect 22096 40768 22112 40832
rect 22176 40768 22192 40832
rect 22256 40768 22262 40832
rect 21946 40767 22262 40768
rect 26946 40832 27262 40833
rect 26946 40768 26952 40832
rect 27016 40768 27032 40832
rect 27096 40768 27112 40832
rect 27176 40768 27192 40832
rect 27256 40768 27262 40832
rect 26946 40767 27262 40768
rect 31946 40832 32262 40833
rect 31946 40768 31952 40832
rect 32016 40768 32032 40832
rect 32096 40768 32112 40832
rect 32176 40768 32192 40832
rect 32256 40768 32262 40832
rect 31946 40767 32262 40768
rect 36946 40832 37262 40833
rect 36946 40768 36952 40832
rect 37016 40768 37032 40832
rect 37096 40768 37112 40832
rect 37176 40768 37192 40832
rect 37256 40768 37262 40832
rect 36946 40767 37262 40768
rect 41946 40832 42262 40833
rect 41946 40768 41952 40832
rect 42016 40768 42032 40832
rect 42096 40768 42112 40832
rect 42176 40768 42192 40832
rect 42256 40768 42262 40832
rect 41946 40767 42262 40768
rect 46946 40832 47262 40833
rect 46946 40768 46952 40832
rect 47016 40768 47032 40832
rect 47096 40768 47112 40832
rect 47176 40768 47192 40832
rect 47256 40768 47262 40832
rect 46946 40767 47262 40768
rect 51946 40832 52262 40833
rect 51946 40768 51952 40832
rect 52016 40768 52032 40832
rect 52096 40768 52112 40832
rect 52176 40768 52192 40832
rect 52256 40768 52262 40832
rect 51946 40767 52262 40768
rect 56946 40832 57262 40833
rect 56946 40768 56952 40832
rect 57016 40768 57032 40832
rect 57096 40768 57112 40832
rect 57176 40768 57192 40832
rect 57256 40768 57262 40832
rect 59200 40808 60000 40838
rect 56946 40767 57262 40768
rect 2606 40288 2922 40289
rect 2606 40224 2612 40288
rect 2676 40224 2692 40288
rect 2756 40224 2772 40288
rect 2836 40224 2852 40288
rect 2916 40224 2922 40288
rect 2606 40223 2922 40224
rect 7606 40288 7922 40289
rect 7606 40224 7612 40288
rect 7676 40224 7692 40288
rect 7756 40224 7772 40288
rect 7836 40224 7852 40288
rect 7916 40224 7922 40288
rect 7606 40223 7922 40224
rect 12606 40288 12922 40289
rect 12606 40224 12612 40288
rect 12676 40224 12692 40288
rect 12756 40224 12772 40288
rect 12836 40224 12852 40288
rect 12916 40224 12922 40288
rect 12606 40223 12922 40224
rect 17606 40288 17922 40289
rect 17606 40224 17612 40288
rect 17676 40224 17692 40288
rect 17756 40224 17772 40288
rect 17836 40224 17852 40288
rect 17916 40224 17922 40288
rect 17606 40223 17922 40224
rect 22606 40288 22922 40289
rect 22606 40224 22612 40288
rect 22676 40224 22692 40288
rect 22756 40224 22772 40288
rect 22836 40224 22852 40288
rect 22916 40224 22922 40288
rect 22606 40223 22922 40224
rect 27606 40288 27922 40289
rect 27606 40224 27612 40288
rect 27676 40224 27692 40288
rect 27756 40224 27772 40288
rect 27836 40224 27852 40288
rect 27916 40224 27922 40288
rect 27606 40223 27922 40224
rect 32606 40288 32922 40289
rect 32606 40224 32612 40288
rect 32676 40224 32692 40288
rect 32756 40224 32772 40288
rect 32836 40224 32852 40288
rect 32916 40224 32922 40288
rect 32606 40223 32922 40224
rect 37606 40288 37922 40289
rect 37606 40224 37612 40288
rect 37676 40224 37692 40288
rect 37756 40224 37772 40288
rect 37836 40224 37852 40288
rect 37916 40224 37922 40288
rect 37606 40223 37922 40224
rect 42606 40288 42922 40289
rect 42606 40224 42612 40288
rect 42676 40224 42692 40288
rect 42756 40224 42772 40288
rect 42836 40224 42852 40288
rect 42916 40224 42922 40288
rect 42606 40223 42922 40224
rect 47606 40288 47922 40289
rect 47606 40224 47612 40288
rect 47676 40224 47692 40288
rect 47756 40224 47772 40288
rect 47836 40224 47852 40288
rect 47916 40224 47922 40288
rect 47606 40223 47922 40224
rect 52606 40288 52922 40289
rect 52606 40224 52612 40288
rect 52676 40224 52692 40288
rect 52756 40224 52772 40288
rect 52836 40224 52852 40288
rect 52916 40224 52922 40288
rect 52606 40223 52922 40224
rect 57606 40288 57922 40289
rect 57606 40224 57612 40288
rect 57676 40224 57692 40288
rect 57756 40224 57772 40288
rect 57836 40224 57852 40288
rect 57916 40224 57922 40288
rect 57606 40223 57922 40224
rect 58525 40082 58591 40085
rect 59200 40082 60000 40112
rect 58525 40080 60000 40082
rect 58525 40024 58530 40080
rect 58586 40024 60000 40080
rect 58525 40022 60000 40024
rect 58525 40019 58591 40022
rect 59200 39992 60000 40022
rect 1946 39744 2262 39745
rect 1946 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2262 39744
rect 1946 39679 2262 39680
rect 6946 39744 7262 39745
rect 6946 39680 6952 39744
rect 7016 39680 7032 39744
rect 7096 39680 7112 39744
rect 7176 39680 7192 39744
rect 7256 39680 7262 39744
rect 6946 39679 7262 39680
rect 11946 39744 12262 39745
rect 11946 39680 11952 39744
rect 12016 39680 12032 39744
rect 12096 39680 12112 39744
rect 12176 39680 12192 39744
rect 12256 39680 12262 39744
rect 11946 39679 12262 39680
rect 16946 39744 17262 39745
rect 16946 39680 16952 39744
rect 17016 39680 17032 39744
rect 17096 39680 17112 39744
rect 17176 39680 17192 39744
rect 17256 39680 17262 39744
rect 16946 39679 17262 39680
rect 21946 39744 22262 39745
rect 21946 39680 21952 39744
rect 22016 39680 22032 39744
rect 22096 39680 22112 39744
rect 22176 39680 22192 39744
rect 22256 39680 22262 39744
rect 21946 39679 22262 39680
rect 26946 39744 27262 39745
rect 26946 39680 26952 39744
rect 27016 39680 27032 39744
rect 27096 39680 27112 39744
rect 27176 39680 27192 39744
rect 27256 39680 27262 39744
rect 26946 39679 27262 39680
rect 31946 39744 32262 39745
rect 31946 39680 31952 39744
rect 32016 39680 32032 39744
rect 32096 39680 32112 39744
rect 32176 39680 32192 39744
rect 32256 39680 32262 39744
rect 31946 39679 32262 39680
rect 36946 39744 37262 39745
rect 36946 39680 36952 39744
rect 37016 39680 37032 39744
rect 37096 39680 37112 39744
rect 37176 39680 37192 39744
rect 37256 39680 37262 39744
rect 36946 39679 37262 39680
rect 41946 39744 42262 39745
rect 41946 39680 41952 39744
rect 42016 39680 42032 39744
rect 42096 39680 42112 39744
rect 42176 39680 42192 39744
rect 42256 39680 42262 39744
rect 41946 39679 42262 39680
rect 46946 39744 47262 39745
rect 46946 39680 46952 39744
rect 47016 39680 47032 39744
rect 47096 39680 47112 39744
rect 47176 39680 47192 39744
rect 47256 39680 47262 39744
rect 46946 39679 47262 39680
rect 51946 39744 52262 39745
rect 51946 39680 51952 39744
rect 52016 39680 52032 39744
rect 52096 39680 52112 39744
rect 52176 39680 52192 39744
rect 52256 39680 52262 39744
rect 51946 39679 52262 39680
rect 56946 39744 57262 39745
rect 56946 39680 56952 39744
rect 57016 39680 57032 39744
rect 57096 39680 57112 39744
rect 57176 39680 57192 39744
rect 57256 39680 57262 39744
rect 56946 39679 57262 39680
rect 58525 39266 58591 39269
rect 59200 39266 60000 39296
rect 58525 39264 60000 39266
rect 58525 39208 58530 39264
rect 58586 39208 60000 39264
rect 58525 39206 60000 39208
rect 58525 39203 58591 39206
rect 2606 39200 2922 39201
rect 2606 39136 2612 39200
rect 2676 39136 2692 39200
rect 2756 39136 2772 39200
rect 2836 39136 2852 39200
rect 2916 39136 2922 39200
rect 2606 39135 2922 39136
rect 7606 39200 7922 39201
rect 7606 39136 7612 39200
rect 7676 39136 7692 39200
rect 7756 39136 7772 39200
rect 7836 39136 7852 39200
rect 7916 39136 7922 39200
rect 7606 39135 7922 39136
rect 12606 39200 12922 39201
rect 12606 39136 12612 39200
rect 12676 39136 12692 39200
rect 12756 39136 12772 39200
rect 12836 39136 12852 39200
rect 12916 39136 12922 39200
rect 12606 39135 12922 39136
rect 17606 39200 17922 39201
rect 17606 39136 17612 39200
rect 17676 39136 17692 39200
rect 17756 39136 17772 39200
rect 17836 39136 17852 39200
rect 17916 39136 17922 39200
rect 17606 39135 17922 39136
rect 22606 39200 22922 39201
rect 22606 39136 22612 39200
rect 22676 39136 22692 39200
rect 22756 39136 22772 39200
rect 22836 39136 22852 39200
rect 22916 39136 22922 39200
rect 22606 39135 22922 39136
rect 27606 39200 27922 39201
rect 27606 39136 27612 39200
rect 27676 39136 27692 39200
rect 27756 39136 27772 39200
rect 27836 39136 27852 39200
rect 27916 39136 27922 39200
rect 27606 39135 27922 39136
rect 32606 39200 32922 39201
rect 32606 39136 32612 39200
rect 32676 39136 32692 39200
rect 32756 39136 32772 39200
rect 32836 39136 32852 39200
rect 32916 39136 32922 39200
rect 32606 39135 32922 39136
rect 37606 39200 37922 39201
rect 37606 39136 37612 39200
rect 37676 39136 37692 39200
rect 37756 39136 37772 39200
rect 37836 39136 37852 39200
rect 37916 39136 37922 39200
rect 37606 39135 37922 39136
rect 42606 39200 42922 39201
rect 42606 39136 42612 39200
rect 42676 39136 42692 39200
rect 42756 39136 42772 39200
rect 42836 39136 42852 39200
rect 42916 39136 42922 39200
rect 42606 39135 42922 39136
rect 47606 39200 47922 39201
rect 47606 39136 47612 39200
rect 47676 39136 47692 39200
rect 47756 39136 47772 39200
rect 47836 39136 47852 39200
rect 47916 39136 47922 39200
rect 47606 39135 47922 39136
rect 52606 39200 52922 39201
rect 52606 39136 52612 39200
rect 52676 39136 52692 39200
rect 52756 39136 52772 39200
rect 52836 39136 52852 39200
rect 52916 39136 52922 39200
rect 52606 39135 52922 39136
rect 57606 39200 57922 39201
rect 57606 39136 57612 39200
rect 57676 39136 57692 39200
rect 57756 39136 57772 39200
rect 57836 39136 57852 39200
rect 57916 39136 57922 39200
rect 59200 39176 60000 39206
rect 57606 39135 57922 39136
rect 1946 38656 2262 38657
rect 1946 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2262 38656
rect 1946 38591 2262 38592
rect 6946 38656 7262 38657
rect 6946 38592 6952 38656
rect 7016 38592 7032 38656
rect 7096 38592 7112 38656
rect 7176 38592 7192 38656
rect 7256 38592 7262 38656
rect 6946 38591 7262 38592
rect 11946 38656 12262 38657
rect 11946 38592 11952 38656
rect 12016 38592 12032 38656
rect 12096 38592 12112 38656
rect 12176 38592 12192 38656
rect 12256 38592 12262 38656
rect 11946 38591 12262 38592
rect 16946 38656 17262 38657
rect 16946 38592 16952 38656
rect 17016 38592 17032 38656
rect 17096 38592 17112 38656
rect 17176 38592 17192 38656
rect 17256 38592 17262 38656
rect 16946 38591 17262 38592
rect 21946 38656 22262 38657
rect 21946 38592 21952 38656
rect 22016 38592 22032 38656
rect 22096 38592 22112 38656
rect 22176 38592 22192 38656
rect 22256 38592 22262 38656
rect 21946 38591 22262 38592
rect 26946 38656 27262 38657
rect 26946 38592 26952 38656
rect 27016 38592 27032 38656
rect 27096 38592 27112 38656
rect 27176 38592 27192 38656
rect 27256 38592 27262 38656
rect 26946 38591 27262 38592
rect 31946 38656 32262 38657
rect 31946 38592 31952 38656
rect 32016 38592 32032 38656
rect 32096 38592 32112 38656
rect 32176 38592 32192 38656
rect 32256 38592 32262 38656
rect 31946 38591 32262 38592
rect 36946 38656 37262 38657
rect 36946 38592 36952 38656
rect 37016 38592 37032 38656
rect 37096 38592 37112 38656
rect 37176 38592 37192 38656
rect 37256 38592 37262 38656
rect 36946 38591 37262 38592
rect 41946 38656 42262 38657
rect 41946 38592 41952 38656
rect 42016 38592 42032 38656
rect 42096 38592 42112 38656
rect 42176 38592 42192 38656
rect 42256 38592 42262 38656
rect 41946 38591 42262 38592
rect 46946 38656 47262 38657
rect 46946 38592 46952 38656
rect 47016 38592 47032 38656
rect 47096 38592 47112 38656
rect 47176 38592 47192 38656
rect 47256 38592 47262 38656
rect 46946 38591 47262 38592
rect 51946 38656 52262 38657
rect 51946 38592 51952 38656
rect 52016 38592 52032 38656
rect 52096 38592 52112 38656
rect 52176 38592 52192 38656
rect 52256 38592 52262 38656
rect 51946 38591 52262 38592
rect 56946 38656 57262 38657
rect 56946 38592 56952 38656
rect 57016 38592 57032 38656
rect 57096 38592 57112 38656
rect 57176 38592 57192 38656
rect 57256 38592 57262 38656
rect 56946 38591 57262 38592
rect 58525 38450 58591 38453
rect 59200 38450 60000 38480
rect 58525 38448 60000 38450
rect 58525 38392 58530 38448
rect 58586 38392 60000 38448
rect 58525 38390 60000 38392
rect 58525 38387 58591 38390
rect 59200 38360 60000 38390
rect 2606 38112 2922 38113
rect 2606 38048 2612 38112
rect 2676 38048 2692 38112
rect 2756 38048 2772 38112
rect 2836 38048 2852 38112
rect 2916 38048 2922 38112
rect 2606 38047 2922 38048
rect 7606 38112 7922 38113
rect 7606 38048 7612 38112
rect 7676 38048 7692 38112
rect 7756 38048 7772 38112
rect 7836 38048 7852 38112
rect 7916 38048 7922 38112
rect 7606 38047 7922 38048
rect 12606 38112 12922 38113
rect 12606 38048 12612 38112
rect 12676 38048 12692 38112
rect 12756 38048 12772 38112
rect 12836 38048 12852 38112
rect 12916 38048 12922 38112
rect 12606 38047 12922 38048
rect 17606 38112 17922 38113
rect 17606 38048 17612 38112
rect 17676 38048 17692 38112
rect 17756 38048 17772 38112
rect 17836 38048 17852 38112
rect 17916 38048 17922 38112
rect 17606 38047 17922 38048
rect 22606 38112 22922 38113
rect 22606 38048 22612 38112
rect 22676 38048 22692 38112
rect 22756 38048 22772 38112
rect 22836 38048 22852 38112
rect 22916 38048 22922 38112
rect 22606 38047 22922 38048
rect 27606 38112 27922 38113
rect 27606 38048 27612 38112
rect 27676 38048 27692 38112
rect 27756 38048 27772 38112
rect 27836 38048 27852 38112
rect 27916 38048 27922 38112
rect 27606 38047 27922 38048
rect 32606 38112 32922 38113
rect 32606 38048 32612 38112
rect 32676 38048 32692 38112
rect 32756 38048 32772 38112
rect 32836 38048 32852 38112
rect 32916 38048 32922 38112
rect 32606 38047 32922 38048
rect 37606 38112 37922 38113
rect 37606 38048 37612 38112
rect 37676 38048 37692 38112
rect 37756 38048 37772 38112
rect 37836 38048 37852 38112
rect 37916 38048 37922 38112
rect 37606 38047 37922 38048
rect 42606 38112 42922 38113
rect 42606 38048 42612 38112
rect 42676 38048 42692 38112
rect 42756 38048 42772 38112
rect 42836 38048 42852 38112
rect 42916 38048 42922 38112
rect 42606 38047 42922 38048
rect 47606 38112 47922 38113
rect 47606 38048 47612 38112
rect 47676 38048 47692 38112
rect 47756 38048 47772 38112
rect 47836 38048 47852 38112
rect 47916 38048 47922 38112
rect 47606 38047 47922 38048
rect 52606 38112 52922 38113
rect 52606 38048 52612 38112
rect 52676 38048 52692 38112
rect 52756 38048 52772 38112
rect 52836 38048 52852 38112
rect 52916 38048 52922 38112
rect 52606 38047 52922 38048
rect 57606 38112 57922 38113
rect 57606 38048 57612 38112
rect 57676 38048 57692 38112
rect 57756 38048 57772 38112
rect 57836 38048 57852 38112
rect 57916 38048 57922 38112
rect 57606 38047 57922 38048
rect 58525 37634 58591 37637
rect 59200 37634 60000 37664
rect 58525 37632 60000 37634
rect 58525 37576 58530 37632
rect 58586 37576 60000 37632
rect 58525 37574 60000 37576
rect 58525 37571 58591 37574
rect 1946 37568 2262 37569
rect 1946 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2262 37568
rect 1946 37503 2262 37504
rect 6946 37568 7262 37569
rect 6946 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7262 37568
rect 6946 37503 7262 37504
rect 11946 37568 12262 37569
rect 11946 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12262 37568
rect 11946 37503 12262 37504
rect 16946 37568 17262 37569
rect 16946 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17262 37568
rect 16946 37503 17262 37504
rect 21946 37568 22262 37569
rect 21946 37504 21952 37568
rect 22016 37504 22032 37568
rect 22096 37504 22112 37568
rect 22176 37504 22192 37568
rect 22256 37504 22262 37568
rect 21946 37503 22262 37504
rect 26946 37568 27262 37569
rect 26946 37504 26952 37568
rect 27016 37504 27032 37568
rect 27096 37504 27112 37568
rect 27176 37504 27192 37568
rect 27256 37504 27262 37568
rect 26946 37503 27262 37504
rect 31946 37568 32262 37569
rect 31946 37504 31952 37568
rect 32016 37504 32032 37568
rect 32096 37504 32112 37568
rect 32176 37504 32192 37568
rect 32256 37504 32262 37568
rect 31946 37503 32262 37504
rect 36946 37568 37262 37569
rect 36946 37504 36952 37568
rect 37016 37504 37032 37568
rect 37096 37504 37112 37568
rect 37176 37504 37192 37568
rect 37256 37504 37262 37568
rect 36946 37503 37262 37504
rect 41946 37568 42262 37569
rect 41946 37504 41952 37568
rect 42016 37504 42032 37568
rect 42096 37504 42112 37568
rect 42176 37504 42192 37568
rect 42256 37504 42262 37568
rect 41946 37503 42262 37504
rect 46946 37568 47262 37569
rect 46946 37504 46952 37568
rect 47016 37504 47032 37568
rect 47096 37504 47112 37568
rect 47176 37504 47192 37568
rect 47256 37504 47262 37568
rect 46946 37503 47262 37504
rect 51946 37568 52262 37569
rect 51946 37504 51952 37568
rect 52016 37504 52032 37568
rect 52096 37504 52112 37568
rect 52176 37504 52192 37568
rect 52256 37504 52262 37568
rect 51946 37503 52262 37504
rect 56946 37568 57262 37569
rect 56946 37504 56952 37568
rect 57016 37504 57032 37568
rect 57096 37504 57112 37568
rect 57176 37504 57192 37568
rect 57256 37504 57262 37568
rect 59200 37544 60000 37574
rect 56946 37503 57262 37504
rect 2606 37024 2922 37025
rect 2606 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2922 37024
rect 2606 36959 2922 36960
rect 7606 37024 7922 37025
rect 7606 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7922 37024
rect 7606 36959 7922 36960
rect 12606 37024 12922 37025
rect 12606 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12922 37024
rect 12606 36959 12922 36960
rect 17606 37024 17922 37025
rect 17606 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17922 37024
rect 17606 36959 17922 36960
rect 22606 37024 22922 37025
rect 22606 36960 22612 37024
rect 22676 36960 22692 37024
rect 22756 36960 22772 37024
rect 22836 36960 22852 37024
rect 22916 36960 22922 37024
rect 22606 36959 22922 36960
rect 27606 37024 27922 37025
rect 27606 36960 27612 37024
rect 27676 36960 27692 37024
rect 27756 36960 27772 37024
rect 27836 36960 27852 37024
rect 27916 36960 27922 37024
rect 27606 36959 27922 36960
rect 32606 37024 32922 37025
rect 32606 36960 32612 37024
rect 32676 36960 32692 37024
rect 32756 36960 32772 37024
rect 32836 36960 32852 37024
rect 32916 36960 32922 37024
rect 32606 36959 32922 36960
rect 37606 37024 37922 37025
rect 37606 36960 37612 37024
rect 37676 36960 37692 37024
rect 37756 36960 37772 37024
rect 37836 36960 37852 37024
rect 37916 36960 37922 37024
rect 37606 36959 37922 36960
rect 42606 37024 42922 37025
rect 42606 36960 42612 37024
rect 42676 36960 42692 37024
rect 42756 36960 42772 37024
rect 42836 36960 42852 37024
rect 42916 36960 42922 37024
rect 42606 36959 42922 36960
rect 47606 37024 47922 37025
rect 47606 36960 47612 37024
rect 47676 36960 47692 37024
rect 47756 36960 47772 37024
rect 47836 36960 47852 37024
rect 47916 36960 47922 37024
rect 47606 36959 47922 36960
rect 52606 37024 52922 37025
rect 52606 36960 52612 37024
rect 52676 36960 52692 37024
rect 52756 36960 52772 37024
rect 52836 36960 52852 37024
rect 52916 36960 52922 37024
rect 52606 36959 52922 36960
rect 57606 37024 57922 37025
rect 57606 36960 57612 37024
rect 57676 36960 57692 37024
rect 57756 36960 57772 37024
rect 57836 36960 57852 37024
rect 57916 36960 57922 37024
rect 57606 36959 57922 36960
rect 58525 36818 58591 36821
rect 59200 36818 60000 36848
rect 58525 36816 60000 36818
rect 58525 36760 58530 36816
rect 58586 36760 60000 36816
rect 58525 36758 60000 36760
rect 58525 36755 58591 36758
rect 59200 36728 60000 36758
rect 1946 36480 2262 36481
rect 1946 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2262 36480
rect 1946 36415 2262 36416
rect 6946 36480 7262 36481
rect 6946 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7262 36480
rect 6946 36415 7262 36416
rect 11946 36480 12262 36481
rect 11946 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12262 36480
rect 11946 36415 12262 36416
rect 16946 36480 17262 36481
rect 16946 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17262 36480
rect 16946 36415 17262 36416
rect 21946 36480 22262 36481
rect 21946 36416 21952 36480
rect 22016 36416 22032 36480
rect 22096 36416 22112 36480
rect 22176 36416 22192 36480
rect 22256 36416 22262 36480
rect 21946 36415 22262 36416
rect 26946 36480 27262 36481
rect 26946 36416 26952 36480
rect 27016 36416 27032 36480
rect 27096 36416 27112 36480
rect 27176 36416 27192 36480
rect 27256 36416 27262 36480
rect 26946 36415 27262 36416
rect 31946 36480 32262 36481
rect 31946 36416 31952 36480
rect 32016 36416 32032 36480
rect 32096 36416 32112 36480
rect 32176 36416 32192 36480
rect 32256 36416 32262 36480
rect 31946 36415 32262 36416
rect 36946 36480 37262 36481
rect 36946 36416 36952 36480
rect 37016 36416 37032 36480
rect 37096 36416 37112 36480
rect 37176 36416 37192 36480
rect 37256 36416 37262 36480
rect 36946 36415 37262 36416
rect 41946 36480 42262 36481
rect 41946 36416 41952 36480
rect 42016 36416 42032 36480
rect 42096 36416 42112 36480
rect 42176 36416 42192 36480
rect 42256 36416 42262 36480
rect 41946 36415 42262 36416
rect 46946 36480 47262 36481
rect 46946 36416 46952 36480
rect 47016 36416 47032 36480
rect 47096 36416 47112 36480
rect 47176 36416 47192 36480
rect 47256 36416 47262 36480
rect 46946 36415 47262 36416
rect 51946 36480 52262 36481
rect 51946 36416 51952 36480
rect 52016 36416 52032 36480
rect 52096 36416 52112 36480
rect 52176 36416 52192 36480
rect 52256 36416 52262 36480
rect 51946 36415 52262 36416
rect 56946 36480 57262 36481
rect 56946 36416 56952 36480
rect 57016 36416 57032 36480
rect 57096 36416 57112 36480
rect 57176 36416 57192 36480
rect 57256 36416 57262 36480
rect 56946 36415 57262 36416
rect 58525 36002 58591 36005
rect 59200 36002 60000 36032
rect 58525 36000 60000 36002
rect 58525 35944 58530 36000
rect 58586 35944 60000 36000
rect 58525 35942 60000 35944
rect 58525 35939 58591 35942
rect 2606 35936 2922 35937
rect 2606 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2922 35936
rect 2606 35871 2922 35872
rect 7606 35936 7922 35937
rect 7606 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7922 35936
rect 7606 35871 7922 35872
rect 12606 35936 12922 35937
rect 12606 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12922 35936
rect 12606 35871 12922 35872
rect 17606 35936 17922 35937
rect 17606 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17922 35936
rect 17606 35871 17922 35872
rect 22606 35936 22922 35937
rect 22606 35872 22612 35936
rect 22676 35872 22692 35936
rect 22756 35872 22772 35936
rect 22836 35872 22852 35936
rect 22916 35872 22922 35936
rect 22606 35871 22922 35872
rect 27606 35936 27922 35937
rect 27606 35872 27612 35936
rect 27676 35872 27692 35936
rect 27756 35872 27772 35936
rect 27836 35872 27852 35936
rect 27916 35872 27922 35936
rect 27606 35871 27922 35872
rect 32606 35936 32922 35937
rect 32606 35872 32612 35936
rect 32676 35872 32692 35936
rect 32756 35872 32772 35936
rect 32836 35872 32852 35936
rect 32916 35872 32922 35936
rect 32606 35871 32922 35872
rect 37606 35936 37922 35937
rect 37606 35872 37612 35936
rect 37676 35872 37692 35936
rect 37756 35872 37772 35936
rect 37836 35872 37852 35936
rect 37916 35872 37922 35936
rect 37606 35871 37922 35872
rect 42606 35936 42922 35937
rect 42606 35872 42612 35936
rect 42676 35872 42692 35936
rect 42756 35872 42772 35936
rect 42836 35872 42852 35936
rect 42916 35872 42922 35936
rect 42606 35871 42922 35872
rect 47606 35936 47922 35937
rect 47606 35872 47612 35936
rect 47676 35872 47692 35936
rect 47756 35872 47772 35936
rect 47836 35872 47852 35936
rect 47916 35872 47922 35936
rect 47606 35871 47922 35872
rect 52606 35936 52922 35937
rect 52606 35872 52612 35936
rect 52676 35872 52692 35936
rect 52756 35872 52772 35936
rect 52836 35872 52852 35936
rect 52916 35872 52922 35936
rect 52606 35871 52922 35872
rect 57606 35936 57922 35937
rect 57606 35872 57612 35936
rect 57676 35872 57692 35936
rect 57756 35872 57772 35936
rect 57836 35872 57852 35936
rect 57916 35872 57922 35936
rect 59200 35912 60000 35942
rect 57606 35871 57922 35872
rect 1946 35392 2262 35393
rect 1946 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2262 35392
rect 1946 35327 2262 35328
rect 6946 35392 7262 35393
rect 6946 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7262 35392
rect 6946 35327 7262 35328
rect 11946 35392 12262 35393
rect 11946 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12262 35392
rect 11946 35327 12262 35328
rect 16946 35392 17262 35393
rect 16946 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17262 35392
rect 16946 35327 17262 35328
rect 21946 35392 22262 35393
rect 21946 35328 21952 35392
rect 22016 35328 22032 35392
rect 22096 35328 22112 35392
rect 22176 35328 22192 35392
rect 22256 35328 22262 35392
rect 21946 35327 22262 35328
rect 26946 35392 27262 35393
rect 26946 35328 26952 35392
rect 27016 35328 27032 35392
rect 27096 35328 27112 35392
rect 27176 35328 27192 35392
rect 27256 35328 27262 35392
rect 26946 35327 27262 35328
rect 31946 35392 32262 35393
rect 31946 35328 31952 35392
rect 32016 35328 32032 35392
rect 32096 35328 32112 35392
rect 32176 35328 32192 35392
rect 32256 35328 32262 35392
rect 31946 35327 32262 35328
rect 36946 35392 37262 35393
rect 36946 35328 36952 35392
rect 37016 35328 37032 35392
rect 37096 35328 37112 35392
rect 37176 35328 37192 35392
rect 37256 35328 37262 35392
rect 36946 35327 37262 35328
rect 41946 35392 42262 35393
rect 41946 35328 41952 35392
rect 42016 35328 42032 35392
rect 42096 35328 42112 35392
rect 42176 35328 42192 35392
rect 42256 35328 42262 35392
rect 41946 35327 42262 35328
rect 46946 35392 47262 35393
rect 46946 35328 46952 35392
rect 47016 35328 47032 35392
rect 47096 35328 47112 35392
rect 47176 35328 47192 35392
rect 47256 35328 47262 35392
rect 46946 35327 47262 35328
rect 51946 35392 52262 35393
rect 51946 35328 51952 35392
rect 52016 35328 52032 35392
rect 52096 35328 52112 35392
rect 52176 35328 52192 35392
rect 52256 35328 52262 35392
rect 51946 35327 52262 35328
rect 56946 35392 57262 35393
rect 56946 35328 56952 35392
rect 57016 35328 57032 35392
rect 57096 35328 57112 35392
rect 57176 35328 57192 35392
rect 57256 35328 57262 35392
rect 56946 35327 57262 35328
rect 58525 35186 58591 35189
rect 59200 35186 60000 35216
rect 58525 35184 60000 35186
rect 58525 35128 58530 35184
rect 58586 35128 60000 35184
rect 58525 35126 60000 35128
rect 58525 35123 58591 35126
rect 59200 35096 60000 35126
rect 2606 34848 2922 34849
rect 2606 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2922 34848
rect 2606 34783 2922 34784
rect 7606 34848 7922 34849
rect 7606 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7922 34848
rect 7606 34783 7922 34784
rect 12606 34848 12922 34849
rect 12606 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12922 34848
rect 12606 34783 12922 34784
rect 17606 34848 17922 34849
rect 17606 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17922 34848
rect 17606 34783 17922 34784
rect 22606 34848 22922 34849
rect 22606 34784 22612 34848
rect 22676 34784 22692 34848
rect 22756 34784 22772 34848
rect 22836 34784 22852 34848
rect 22916 34784 22922 34848
rect 22606 34783 22922 34784
rect 27606 34848 27922 34849
rect 27606 34784 27612 34848
rect 27676 34784 27692 34848
rect 27756 34784 27772 34848
rect 27836 34784 27852 34848
rect 27916 34784 27922 34848
rect 27606 34783 27922 34784
rect 32606 34848 32922 34849
rect 32606 34784 32612 34848
rect 32676 34784 32692 34848
rect 32756 34784 32772 34848
rect 32836 34784 32852 34848
rect 32916 34784 32922 34848
rect 32606 34783 32922 34784
rect 37606 34848 37922 34849
rect 37606 34784 37612 34848
rect 37676 34784 37692 34848
rect 37756 34784 37772 34848
rect 37836 34784 37852 34848
rect 37916 34784 37922 34848
rect 37606 34783 37922 34784
rect 42606 34848 42922 34849
rect 42606 34784 42612 34848
rect 42676 34784 42692 34848
rect 42756 34784 42772 34848
rect 42836 34784 42852 34848
rect 42916 34784 42922 34848
rect 42606 34783 42922 34784
rect 47606 34848 47922 34849
rect 47606 34784 47612 34848
rect 47676 34784 47692 34848
rect 47756 34784 47772 34848
rect 47836 34784 47852 34848
rect 47916 34784 47922 34848
rect 47606 34783 47922 34784
rect 52606 34848 52922 34849
rect 52606 34784 52612 34848
rect 52676 34784 52692 34848
rect 52756 34784 52772 34848
rect 52836 34784 52852 34848
rect 52916 34784 52922 34848
rect 52606 34783 52922 34784
rect 57606 34848 57922 34849
rect 57606 34784 57612 34848
rect 57676 34784 57692 34848
rect 57756 34784 57772 34848
rect 57836 34784 57852 34848
rect 57916 34784 57922 34848
rect 57606 34783 57922 34784
rect 58525 34370 58591 34373
rect 59200 34370 60000 34400
rect 58525 34368 60000 34370
rect 58525 34312 58530 34368
rect 58586 34312 60000 34368
rect 58525 34310 60000 34312
rect 58525 34307 58591 34310
rect 1946 34304 2262 34305
rect 1946 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2262 34304
rect 1946 34239 2262 34240
rect 6946 34304 7262 34305
rect 6946 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7262 34304
rect 6946 34239 7262 34240
rect 11946 34304 12262 34305
rect 11946 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12262 34304
rect 11946 34239 12262 34240
rect 16946 34304 17262 34305
rect 16946 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17262 34304
rect 16946 34239 17262 34240
rect 21946 34304 22262 34305
rect 21946 34240 21952 34304
rect 22016 34240 22032 34304
rect 22096 34240 22112 34304
rect 22176 34240 22192 34304
rect 22256 34240 22262 34304
rect 21946 34239 22262 34240
rect 26946 34304 27262 34305
rect 26946 34240 26952 34304
rect 27016 34240 27032 34304
rect 27096 34240 27112 34304
rect 27176 34240 27192 34304
rect 27256 34240 27262 34304
rect 26946 34239 27262 34240
rect 31946 34304 32262 34305
rect 31946 34240 31952 34304
rect 32016 34240 32032 34304
rect 32096 34240 32112 34304
rect 32176 34240 32192 34304
rect 32256 34240 32262 34304
rect 31946 34239 32262 34240
rect 36946 34304 37262 34305
rect 36946 34240 36952 34304
rect 37016 34240 37032 34304
rect 37096 34240 37112 34304
rect 37176 34240 37192 34304
rect 37256 34240 37262 34304
rect 36946 34239 37262 34240
rect 41946 34304 42262 34305
rect 41946 34240 41952 34304
rect 42016 34240 42032 34304
rect 42096 34240 42112 34304
rect 42176 34240 42192 34304
rect 42256 34240 42262 34304
rect 41946 34239 42262 34240
rect 46946 34304 47262 34305
rect 46946 34240 46952 34304
rect 47016 34240 47032 34304
rect 47096 34240 47112 34304
rect 47176 34240 47192 34304
rect 47256 34240 47262 34304
rect 46946 34239 47262 34240
rect 51946 34304 52262 34305
rect 51946 34240 51952 34304
rect 52016 34240 52032 34304
rect 52096 34240 52112 34304
rect 52176 34240 52192 34304
rect 52256 34240 52262 34304
rect 51946 34239 52262 34240
rect 56946 34304 57262 34305
rect 56946 34240 56952 34304
rect 57016 34240 57032 34304
rect 57096 34240 57112 34304
rect 57176 34240 57192 34304
rect 57256 34240 57262 34304
rect 59200 34280 60000 34310
rect 56946 34239 57262 34240
rect 2606 33760 2922 33761
rect 2606 33696 2612 33760
rect 2676 33696 2692 33760
rect 2756 33696 2772 33760
rect 2836 33696 2852 33760
rect 2916 33696 2922 33760
rect 2606 33695 2922 33696
rect 7606 33760 7922 33761
rect 7606 33696 7612 33760
rect 7676 33696 7692 33760
rect 7756 33696 7772 33760
rect 7836 33696 7852 33760
rect 7916 33696 7922 33760
rect 7606 33695 7922 33696
rect 12606 33760 12922 33761
rect 12606 33696 12612 33760
rect 12676 33696 12692 33760
rect 12756 33696 12772 33760
rect 12836 33696 12852 33760
rect 12916 33696 12922 33760
rect 12606 33695 12922 33696
rect 17606 33760 17922 33761
rect 17606 33696 17612 33760
rect 17676 33696 17692 33760
rect 17756 33696 17772 33760
rect 17836 33696 17852 33760
rect 17916 33696 17922 33760
rect 17606 33695 17922 33696
rect 22606 33760 22922 33761
rect 22606 33696 22612 33760
rect 22676 33696 22692 33760
rect 22756 33696 22772 33760
rect 22836 33696 22852 33760
rect 22916 33696 22922 33760
rect 22606 33695 22922 33696
rect 27606 33760 27922 33761
rect 27606 33696 27612 33760
rect 27676 33696 27692 33760
rect 27756 33696 27772 33760
rect 27836 33696 27852 33760
rect 27916 33696 27922 33760
rect 27606 33695 27922 33696
rect 32606 33760 32922 33761
rect 32606 33696 32612 33760
rect 32676 33696 32692 33760
rect 32756 33696 32772 33760
rect 32836 33696 32852 33760
rect 32916 33696 32922 33760
rect 32606 33695 32922 33696
rect 37606 33760 37922 33761
rect 37606 33696 37612 33760
rect 37676 33696 37692 33760
rect 37756 33696 37772 33760
rect 37836 33696 37852 33760
rect 37916 33696 37922 33760
rect 37606 33695 37922 33696
rect 42606 33760 42922 33761
rect 42606 33696 42612 33760
rect 42676 33696 42692 33760
rect 42756 33696 42772 33760
rect 42836 33696 42852 33760
rect 42916 33696 42922 33760
rect 42606 33695 42922 33696
rect 47606 33760 47922 33761
rect 47606 33696 47612 33760
rect 47676 33696 47692 33760
rect 47756 33696 47772 33760
rect 47836 33696 47852 33760
rect 47916 33696 47922 33760
rect 47606 33695 47922 33696
rect 52606 33760 52922 33761
rect 52606 33696 52612 33760
rect 52676 33696 52692 33760
rect 52756 33696 52772 33760
rect 52836 33696 52852 33760
rect 52916 33696 52922 33760
rect 52606 33695 52922 33696
rect 57606 33760 57922 33761
rect 57606 33696 57612 33760
rect 57676 33696 57692 33760
rect 57756 33696 57772 33760
rect 57836 33696 57852 33760
rect 57916 33696 57922 33760
rect 57606 33695 57922 33696
rect 58525 33554 58591 33557
rect 59200 33554 60000 33584
rect 58525 33552 60000 33554
rect 58525 33496 58530 33552
rect 58586 33496 60000 33552
rect 58525 33494 60000 33496
rect 58525 33491 58591 33494
rect 59200 33464 60000 33494
rect 1946 33216 2262 33217
rect 1946 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2262 33216
rect 1946 33151 2262 33152
rect 6946 33216 7262 33217
rect 6946 33152 6952 33216
rect 7016 33152 7032 33216
rect 7096 33152 7112 33216
rect 7176 33152 7192 33216
rect 7256 33152 7262 33216
rect 6946 33151 7262 33152
rect 11946 33216 12262 33217
rect 11946 33152 11952 33216
rect 12016 33152 12032 33216
rect 12096 33152 12112 33216
rect 12176 33152 12192 33216
rect 12256 33152 12262 33216
rect 11946 33151 12262 33152
rect 16946 33216 17262 33217
rect 16946 33152 16952 33216
rect 17016 33152 17032 33216
rect 17096 33152 17112 33216
rect 17176 33152 17192 33216
rect 17256 33152 17262 33216
rect 16946 33151 17262 33152
rect 21946 33216 22262 33217
rect 21946 33152 21952 33216
rect 22016 33152 22032 33216
rect 22096 33152 22112 33216
rect 22176 33152 22192 33216
rect 22256 33152 22262 33216
rect 21946 33151 22262 33152
rect 26946 33216 27262 33217
rect 26946 33152 26952 33216
rect 27016 33152 27032 33216
rect 27096 33152 27112 33216
rect 27176 33152 27192 33216
rect 27256 33152 27262 33216
rect 26946 33151 27262 33152
rect 31946 33216 32262 33217
rect 31946 33152 31952 33216
rect 32016 33152 32032 33216
rect 32096 33152 32112 33216
rect 32176 33152 32192 33216
rect 32256 33152 32262 33216
rect 31946 33151 32262 33152
rect 36946 33216 37262 33217
rect 36946 33152 36952 33216
rect 37016 33152 37032 33216
rect 37096 33152 37112 33216
rect 37176 33152 37192 33216
rect 37256 33152 37262 33216
rect 36946 33151 37262 33152
rect 41946 33216 42262 33217
rect 41946 33152 41952 33216
rect 42016 33152 42032 33216
rect 42096 33152 42112 33216
rect 42176 33152 42192 33216
rect 42256 33152 42262 33216
rect 41946 33151 42262 33152
rect 46946 33216 47262 33217
rect 46946 33152 46952 33216
rect 47016 33152 47032 33216
rect 47096 33152 47112 33216
rect 47176 33152 47192 33216
rect 47256 33152 47262 33216
rect 46946 33151 47262 33152
rect 51946 33216 52262 33217
rect 51946 33152 51952 33216
rect 52016 33152 52032 33216
rect 52096 33152 52112 33216
rect 52176 33152 52192 33216
rect 52256 33152 52262 33216
rect 51946 33151 52262 33152
rect 56946 33216 57262 33217
rect 56946 33152 56952 33216
rect 57016 33152 57032 33216
rect 57096 33152 57112 33216
rect 57176 33152 57192 33216
rect 57256 33152 57262 33216
rect 56946 33151 57262 33152
rect 58525 32738 58591 32741
rect 59200 32738 60000 32768
rect 58525 32736 60000 32738
rect 58525 32680 58530 32736
rect 58586 32680 60000 32736
rect 58525 32678 60000 32680
rect 58525 32675 58591 32678
rect 2606 32672 2922 32673
rect 2606 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2922 32672
rect 2606 32607 2922 32608
rect 7606 32672 7922 32673
rect 7606 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7922 32672
rect 7606 32607 7922 32608
rect 12606 32672 12922 32673
rect 12606 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12922 32672
rect 12606 32607 12922 32608
rect 17606 32672 17922 32673
rect 17606 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17922 32672
rect 17606 32607 17922 32608
rect 22606 32672 22922 32673
rect 22606 32608 22612 32672
rect 22676 32608 22692 32672
rect 22756 32608 22772 32672
rect 22836 32608 22852 32672
rect 22916 32608 22922 32672
rect 22606 32607 22922 32608
rect 27606 32672 27922 32673
rect 27606 32608 27612 32672
rect 27676 32608 27692 32672
rect 27756 32608 27772 32672
rect 27836 32608 27852 32672
rect 27916 32608 27922 32672
rect 27606 32607 27922 32608
rect 32606 32672 32922 32673
rect 32606 32608 32612 32672
rect 32676 32608 32692 32672
rect 32756 32608 32772 32672
rect 32836 32608 32852 32672
rect 32916 32608 32922 32672
rect 32606 32607 32922 32608
rect 37606 32672 37922 32673
rect 37606 32608 37612 32672
rect 37676 32608 37692 32672
rect 37756 32608 37772 32672
rect 37836 32608 37852 32672
rect 37916 32608 37922 32672
rect 37606 32607 37922 32608
rect 42606 32672 42922 32673
rect 42606 32608 42612 32672
rect 42676 32608 42692 32672
rect 42756 32608 42772 32672
rect 42836 32608 42852 32672
rect 42916 32608 42922 32672
rect 42606 32607 42922 32608
rect 47606 32672 47922 32673
rect 47606 32608 47612 32672
rect 47676 32608 47692 32672
rect 47756 32608 47772 32672
rect 47836 32608 47852 32672
rect 47916 32608 47922 32672
rect 47606 32607 47922 32608
rect 52606 32672 52922 32673
rect 52606 32608 52612 32672
rect 52676 32608 52692 32672
rect 52756 32608 52772 32672
rect 52836 32608 52852 32672
rect 52916 32608 52922 32672
rect 52606 32607 52922 32608
rect 57606 32672 57922 32673
rect 57606 32608 57612 32672
rect 57676 32608 57692 32672
rect 57756 32608 57772 32672
rect 57836 32608 57852 32672
rect 57916 32608 57922 32672
rect 59200 32648 60000 32678
rect 57606 32607 57922 32608
rect 1946 32128 2262 32129
rect 1946 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2262 32128
rect 1946 32063 2262 32064
rect 6946 32128 7262 32129
rect 6946 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7262 32128
rect 6946 32063 7262 32064
rect 11946 32128 12262 32129
rect 11946 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12262 32128
rect 11946 32063 12262 32064
rect 16946 32128 17262 32129
rect 16946 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17262 32128
rect 16946 32063 17262 32064
rect 21946 32128 22262 32129
rect 21946 32064 21952 32128
rect 22016 32064 22032 32128
rect 22096 32064 22112 32128
rect 22176 32064 22192 32128
rect 22256 32064 22262 32128
rect 21946 32063 22262 32064
rect 26946 32128 27262 32129
rect 26946 32064 26952 32128
rect 27016 32064 27032 32128
rect 27096 32064 27112 32128
rect 27176 32064 27192 32128
rect 27256 32064 27262 32128
rect 26946 32063 27262 32064
rect 31946 32128 32262 32129
rect 31946 32064 31952 32128
rect 32016 32064 32032 32128
rect 32096 32064 32112 32128
rect 32176 32064 32192 32128
rect 32256 32064 32262 32128
rect 31946 32063 32262 32064
rect 36946 32128 37262 32129
rect 36946 32064 36952 32128
rect 37016 32064 37032 32128
rect 37096 32064 37112 32128
rect 37176 32064 37192 32128
rect 37256 32064 37262 32128
rect 36946 32063 37262 32064
rect 41946 32128 42262 32129
rect 41946 32064 41952 32128
rect 42016 32064 42032 32128
rect 42096 32064 42112 32128
rect 42176 32064 42192 32128
rect 42256 32064 42262 32128
rect 41946 32063 42262 32064
rect 46946 32128 47262 32129
rect 46946 32064 46952 32128
rect 47016 32064 47032 32128
rect 47096 32064 47112 32128
rect 47176 32064 47192 32128
rect 47256 32064 47262 32128
rect 46946 32063 47262 32064
rect 51946 32128 52262 32129
rect 51946 32064 51952 32128
rect 52016 32064 52032 32128
rect 52096 32064 52112 32128
rect 52176 32064 52192 32128
rect 52256 32064 52262 32128
rect 51946 32063 52262 32064
rect 56946 32128 57262 32129
rect 56946 32064 56952 32128
rect 57016 32064 57032 32128
rect 57096 32064 57112 32128
rect 57176 32064 57192 32128
rect 57256 32064 57262 32128
rect 56946 32063 57262 32064
rect 58525 31922 58591 31925
rect 59200 31922 60000 31952
rect 58525 31920 60000 31922
rect 58525 31864 58530 31920
rect 58586 31864 60000 31920
rect 58525 31862 60000 31864
rect 58525 31859 58591 31862
rect 59200 31832 60000 31862
rect 2606 31584 2922 31585
rect 2606 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2922 31584
rect 2606 31519 2922 31520
rect 7606 31584 7922 31585
rect 7606 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7922 31584
rect 7606 31519 7922 31520
rect 12606 31584 12922 31585
rect 12606 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12922 31584
rect 12606 31519 12922 31520
rect 17606 31584 17922 31585
rect 17606 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17922 31584
rect 17606 31519 17922 31520
rect 22606 31584 22922 31585
rect 22606 31520 22612 31584
rect 22676 31520 22692 31584
rect 22756 31520 22772 31584
rect 22836 31520 22852 31584
rect 22916 31520 22922 31584
rect 22606 31519 22922 31520
rect 27606 31584 27922 31585
rect 27606 31520 27612 31584
rect 27676 31520 27692 31584
rect 27756 31520 27772 31584
rect 27836 31520 27852 31584
rect 27916 31520 27922 31584
rect 27606 31519 27922 31520
rect 32606 31584 32922 31585
rect 32606 31520 32612 31584
rect 32676 31520 32692 31584
rect 32756 31520 32772 31584
rect 32836 31520 32852 31584
rect 32916 31520 32922 31584
rect 32606 31519 32922 31520
rect 37606 31584 37922 31585
rect 37606 31520 37612 31584
rect 37676 31520 37692 31584
rect 37756 31520 37772 31584
rect 37836 31520 37852 31584
rect 37916 31520 37922 31584
rect 37606 31519 37922 31520
rect 42606 31584 42922 31585
rect 42606 31520 42612 31584
rect 42676 31520 42692 31584
rect 42756 31520 42772 31584
rect 42836 31520 42852 31584
rect 42916 31520 42922 31584
rect 42606 31519 42922 31520
rect 47606 31584 47922 31585
rect 47606 31520 47612 31584
rect 47676 31520 47692 31584
rect 47756 31520 47772 31584
rect 47836 31520 47852 31584
rect 47916 31520 47922 31584
rect 47606 31519 47922 31520
rect 52606 31584 52922 31585
rect 52606 31520 52612 31584
rect 52676 31520 52692 31584
rect 52756 31520 52772 31584
rect 52836 31520 52852 31584
rect 52916 31520 52922 31584
rect 52606 31519 52922 31520
rect 57606 31584 57922 31585
rect 57606 31520 57612 31584
rect 57676 31520 57692 31584
rect 57756 31520 57772 31584
rect 57836 31520 57852 31584
rect 57916 31520 57922 31584
rect 57606 31519 57922 31520
rect 58525 31106 58591 31109
rect 59200 31106 60000 31136
rect 58525 31104 60000 31106
rect 58525 31048 58530 31104
rect 58586 31048 60000 31104
rect 58525 31046 60000 31048
rect 58525 31043 58591 31046
rect 1946 31040 2262 31041
rect 1946 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2262 31040
rect 1946 30975 2262 30976
rect 6946 31040 7262 31041
rect 6946 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7262 31040
rect 6946 30975 7262 30976
rect 11946 31040 12262 31041
rect 11946 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12262 31040
rect 11946 30975 12262 30976
rect 16946 31040 17262 31041
rect 16946 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17262 31040
rect 16946 30975 17262 30976
rect 21946 31040 22262 31041
rect 21946 30976 21952 31040
rect 22016 30976 22032 31040
rect 22096 30976 22112 31040
rect 22176 30976 22192 31040
rect 22256 30976 22262 31040
rect 21946 30975 22262 30976
rect 26946 31040 27262 31041
rect 26946 30976 26952 31040
rect 27016 30976 27032 31040
rect 27096 30976 27112 31040
rect 27176 30976 27192 31040
rect 27256 30976 27262 31040
rect 26946 30975 27262 30976
rect 31946 31040 32262 31041
rect 31946 30976 31952 31040
rect 32016 30976 32032 31040
rect 32096 30976 32112 31040
rect 32176 30976 32192 31040
rect 32256 30976 32262 31040
rect 31946 30975 32262 30976
rect 36946 31040 37262 31041
rect 36946 30976 36952 31040
rect 37016 30976 37032 31040
rect 37096 30976 37112 31040
rect 37176 30976 37192 31040
rect 37256 30976 37262 31040
rect 36946 30975 37262 30976
rect 41946 31040 42262 31041
rect 41946 30976 41952 31040
rect 42016 30976 42032 31040
rect 42096 30976 42112 31040
rect 42176 30976 42192 31040
rect 42256 30976 42262 31040
rect 41946 30975 42262 30976
rect 46946 31040 47262 31041
rect 46946 30976 46952 31040
rect 47016 30976 47032 31040
rect 47096 30976 47112 31040
rect 47176 30976 47192 31040
rect 47256 30976 47262 31040
rect 46946 30975 47262 30976
rect 51946 31040 52262 31041
rect 51946 30976 51952 31040
rect 52016 30976 52032 31040
rect 52096 30976 52112 31040
rect 52176 30976 52192 31040
rect 52256 30976 52262 31040
rect 51946 30975 52262 30976
rect 56946 31040 57262 31041
rect 56946 30976 56952 31040
rect 57016 30976 57032 31040
rect 57096 30976 57112 31040
rect 57176 30976 57192 31040
rect 57256 30976 57262 31040
rect 59200 31016 60000 31046
rect 56946 30975 57262 30976
rect 2606 30496 2922 30497
rect 2606 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2922 30496
rect 2606 30431 2922 30432
rect 7606 30496 7922 30497
rect 7606 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7922 30496
rect 7606 30431 7922 30432
rect 12606 30496 12922 30497
rect 12606 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12922 30496
rect 12606 30431 12922 30432
rect 17606 30496 17922 30497
rect 17606 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17922 30496
rect 17606 30431 17922 30432
rect 22606 30496 22922 30497
rect 22606 30432 22612 30496
rect 22676 30432 22692 30496
rect 22756 30432 22772 30496
rect 22836 30432 22852 30496
rect 22916 30432 22922 30496
rect 22606 30431 22922 30432
rect 27606 30496 27922 30497
rect 27606 30432 27612 30496
rect 27676 30432 27692 30496
rect 27756 30432 27772 30496
rect 27836 30432 27852 30496
rect 27916 30432 27922 30496
rect 27606 30431 27922 30432
rect 32606 30496 32922 30497
rect 32606 30432 32612 30496
rect 32676 30432 32692 30496
rect 32756 30432 32772 30496
rect 32836 30432 32852 30496
rect 32916 30432 32922 30496
rect 32606 30431 32922 30432
rect 37606 30496 37922 30497
rect 37606 30432 37612 30496
rect 37676 30432 37692 30496
rect 37756 30432 37772 30496
rect 37836 30432 37852 30496
rect 37916 30432 37922 30496
rect 37606 30431 37922 30432
rect 42606 30496 42922 30497
rect 42606 30432 42612 30496
rect 42676 30432 42692 30496
rect 42756 30432 42772 30496
rect 42836 30432 42852 30496
rect 42916 30432 42922 30496
rect 42606 30431 42922 30432
rect 47606 30496 47922 30497
rect 47606 30432 47612 30496
rect 47676 30432 47692 30496
rect 47756 30432 47772 30496
rect 47836 30432 47852 30496
rect 47916 30432 47922 30496
rect 47606 30431 47922 30432
rect 52606 30496 52922 30497
rect 52606 30432 52612 30496
rect 52676 30432 52692 30496
rect 52756 30432 52772 30496
rect 52836 30432 52852 30496
rect 52916 30432 52922 30496
rect 52606 30431 52922 30432
rect 57606 30496 57922 30497
rect 57606 30432 57612 30496
rect 57676 30432 57692 30496
rect 57756 30432 57772 30496
rect 57836 30432 57852 30496
rect 57916 30432 57922 30496
rect 57606 30431 57922 30432
rect 58525 30290 58591 30293
rect 59200 30290 60000 30320
rect 58525 30288 60000 30290
rect 58525 30232 58530 30288
rect 58586 30232 60000 30288
rect 58525 30230 60000 30232
rect 58525 30227 58591 30230
rect 59200 30200 60000 30230
rect 0 29928 800 30048
rect 1946 29952 2262 29953
rect 1946 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2262 29952
rect 1946 29887 2262 29888
rect 6946 29952 7262 29953
rect 6946 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7262 29952
rect 6946 29887 7262 29888
rect 11946 29952 12262 29953
rect 11946 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12262 29952
rect 11946 29887 12262 29888
rect 16946 29952 17262 29953
rect 16946 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17262 29952
rect 16946 29887 17262 29888
rect 21946 29952 22262 29953
rect 21946 29888 21952 29952
rect 22016 29888 22032 29952
rect 22096 29888 22112 29952
rect 22176 29888 22192 29952
rect 22256 29888 22262 29952
rect 21946 29887 22262 29888
rect 26946 29952 27262 29953
rect 26946 29888 26952 29952
rect 27016 29888 27032 29952
rect 27096 29888 27112 29952
rect 27176 29888 27192 29952
rect 27256 29888 27262 29952
rect 26946 29887 27262 29888
rect 31946 29952 32262 29953
rect 31946 29888 31952 29952
rect 32016 29888 32032 29952
rect 32096 29888 32112 29952
rect 32176 29888 32192 29952
rect 32256 29888 32262 29952
rect 31946 29887 32262 29888
rect 36946 29952 37262 29953
rect 36946 29888 36952 29952
rect 37016 29888 37032 29952
rect 37096 29888 37112 29952
rect 37176 29888 37192 29952
rect 37256 29888 37262 29952
rect 36946 29887 37262 29888
rect 41946 29952 42262 29953
rect 41946 29888 41952 29952
rect 42016 29888 42032 29952
rect 42096 29888 42112 29952
rect 42176 29888 42192 29952
rect 42256 29888 42262 29952
rect 41946 29887 42262 29888
rect 46946 29952 47262 29953
rect 46946 29888 46952 29952
rect 47016 29888 47032 29952
rect 47096 29888 47112 29952
rect 47176 29888 47192 29952
rect 47256 29888 47262 29952
rect 46946 29887 47262 29888
rect 51946 29952 52262 29953
rect 51946 29888 51952 29952
rect 52016 29888 52032 29952
rect 52096 29888 52112 29952
rect 52176 29888 52192 29952
rect 52256 29888 52262 29952
rect 51946 29887 52262 29888
rect 56946 29952 57262 29953
rect 56946 29888 56952 29952
rect 57016 29888 57032 29952
rect 57096 29888 57112 29952
rect 57176 29888 57192 29952
rect 57256 29888 57262 29952
rect 56946 29887 57262 29888
rect 58525 29474 58591 29477
rect 59200 29474 60000 29504
rect 58525 29472 60000 29474
rect 58525 29416 58530 29472
rect 58586 29416 60000 29472
rect 58525 29414 60000 29416
rect 58525 29411 58591 29414
rect 2606 29408 2922 29409
rect 2606 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2922 29408
rect 2606 29343 2922 29344
rect 7606 29408 7922 29409
rect 7606 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7922 29408
rect 7606 29343 7922 29344
rect 12606 29408 12922 29409
rect 12606 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12922 29408
rect 12606 29343 12922 29344
rect 17606 29408 17922 29409
rect 17606 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17922 29408
rect 17606 29343 17922 29344
rect 22606 29408 22922 29409
rect 22606 29344 22612 29408
rect 22676 29344 22692 29408
rect 22756 29344 22772 29408
rect 22836 29344 22852 29408
rect 22916 29344 22922 29408
rect 22606 29343 22922 29344
rect 27606 29408 27922 29409
rect 27606 29344 27612 29408
rect 27676 29344 27692 29408
rect 27756 29344 27772 29408
rect 27836 29344 27852 29408
rect 27916 29344 27922 29408
rect 27606 29343 27922 29344
rect 32606 29408 32922 29409
rect 32606 29344 32612 29408
rect 32676 29344 32692 29408
rect 32756 29344 32772 29408
rect 32836 29344 32852 29408
rect 32916 29344 32922 29408
rect 32606 29343 32922 29344
rect 37606 29408 37922 29409
rect 37606 29344 37612 29408
rect 37676 29344 37692 29408
rect 37756 29344 37772 29408
rect 37836 29344 37852 29408
rect 37916 29344 37922 29408
rect 37606 29343 37922 29344
rect 42606 29408 42922 29409
rect 42606 29344 42612 29408
rect 42676 29344 42692 29408
rect 42756 29344 42772 29408
rect 42836 29344 42852 29408
rect 42916 29344 42922 29408
rect 42606 29343 42922 29344
rect 47606 29408 47922 29409
rect 47606 29344 47612 29408
rect 47676 29344 47692 29408
rect 47756 29344 47772 29408
rect 47836 29344 47852 29408
rect 47916 29344 47922 29408
rect 47606 29343 47922 29344
rect 52606 29408 52922 29409
rect 52606 29344 52612 29408
rect 52676 29344 52692 29408
rect 52756 29344 52772 29408
rect 52836 29344 52852 29408
rect 52916 29344 52922 29408
rect 52606 29343 52922 29344
rect 57606 29408 57922 29409
rect 57606 29344 57612 29408
rect 57676 29344 57692 29408
rect 57756 29344 57772 29408
rect 57836 29344 57852 29408
rect 57916 29344 57922 29408
rect 59200 29384 60000 29414
rect 57606 29343 57922 29344
rect 1946 28864 2262 28865
rect 1946 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2262 28864
rect 1946 28799 2262 28800
rect 6946 28864 7262 28865
rect 6946 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7262 28864
rect 6946 28799 7262 28800
rect 11946 28864 12262 28865
rect 11946 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12262 28864
rect 11946 28799 12262 28800
rect 16946 28864 17262 28865
rect 16946 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17262 28864
rect 16946 28799 17262 28800
rect 21946 28864 22262 28865
rect 21946 28800 21952 28864
rect 22016 28800 22032 28864
rect 22096 28800 22112 28864
rect 22176 28800 22192 28864
rect 22256 28800 22262 28864
rect 21946 28799 22262 28800
rect 26946 28864 27262 28865
rect 26946 28800 26952 28864
rect 27016 28800 27032 28864
rect 27096 28800 27112 28864
rect 27176 28800 27192 28864
rect 27256 28800 27262 28864
rect 26946 28799 27262 28800
rect 31946 28864 32262 28865
rect 31946 28800 31952 28864
rect 32016 28800 32032 28864
rect 32096 28800 32112 28864
rect 32176 28800 32192 28864
rect 32256 28800 32262 28864
rect 31946 28799 32262 28800
rect 36946 28864 37262 28865
rect 36946 28800 36952 28864
rect 37016 28800 37032 28864
rect 37096 28800 37112 28864
rect 37176 28800 37192 28864
rect 37256 28800 37262 28864
rect 36946 28799 37262 28800
rect 41946 28864 42262 28865
rect 41946 28800 41952 28864
rect 42016 28800 42032 28864
rect 42096 28800 42112 28864
rect 42176 28800 42192 28864
rect 42256 28800 42262 28864
rect 41946 28799 42262 28800
rect 46946 28864 47262 28865
rect 46946 28800 46952 28864
rect 47016 28800 47032 28864
rect 47096 28800 47112 28864
rect 47176 28800 47192 28864
rect 47256 28800 47262 28864
rect 46946 28799 47262 28800
rect 51946 28864 52262 28865
rect 51946 28800 51952 28864
rect 52016 28800 52032 28864
rect 52096 28800 52112 28864
rect 52176 28800 52192 28864
rect 52256 28800 52262 28864
rect 51946 28799 52262 28800
rect 56946 28864 57262 28865
rect 56946 28800 56952 28864
rect 57016 28800 57032 28864
rect 57096 28800 57112 28864
rect 57176 28800 57192 28864
rect 57256 28800 57262 28864
rect 56946 28799 57262 28800
rect 58525 28658 58591 28661
rect 59200 28658 60000 28688
rect 58525 28656 60000 28658
rect 58525 28600 58530 28656
rect 58586 28600 60000 28656
rect 58525 28598 60000 28600
rect 58525 28595 58591 28598
rect 59200 28568 60000 28598
rect 2606 28320 2922 28321
rect 2606 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2922 28320
rect 2606 28255 2922 28256
rect 7606 28320 7922 28321
rect 7606 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7922 28320
rect 7606 28255 7922 28256
rect 12606 28320 12922 28321
rect 12606 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12922 28320
rect 12606 28255 12922 28256
rect 17606 28320 17922 28321
rect 17606 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17922 28320
rect 17606 28255 17922 28256
rect 22606 28320 22922 28321
rect 22606 28256 22612 28320
rect 22676 28256 22692 28320
rect 22756 28256 22772 28320
rect 22836 28256 22852 28320
rect 22916 28256 22922 28320
rect 22606 28255 22922 28256
rect 27606 28320 27922 28321
rect 27606 28256 27612 28320
rect 27676 28256 27692 28320
rect 27756 28256 27772 28320
rect 27836 28256 27852 28320
rect 27916 28256 27922 28320
rect 27606 28255 27922 28256
rect 32606 28320 32922 28321
rect 32606 28256 32612 28320
rect 32676 28256 32692 28320
rect 32756 28256 32772 28320
rect 32836 28256 32852 28320
rect 32916 28256 32922 28320
rect 32606 28255 32922 28256
rect 37606 28320 37922 28321
rect 37606 28256 37612 28320
rect 37676 28256 37692 28320
rect 37756 28256 37772 28320
rect 37836 28256 37852 28320
rect 37916 28256 37922 28320
rect 37606 28255 37922 28256
rect 42606 28320 42922 28321
rect 42606 28256 42612 28320
rect 42676 28256 42692 28320
rect 42756 28256 42772 28320
rect 42836 28256 42852 28320
rect 42916 28256 42922 28320
rect 42606 28255 42922 28256
rect 47606 28320 47922 28321
rect 47606 28256 47612 28320
rect 47676 28256 47692 28320
rect 47756 28256 47772 28320
rect 47836 28256 47852 28320
rect 47916 28256 47922 28320
rect 47606 28255 47922 28256
rect 52606 28320 52922 28321
rect 52606 28256 52612 28320
rect 52676 28256 52692 28320
rect 52756 28256 52772 28320
rect 52836 28256 52852 28320
rect 52916 28256 52922 28320
rect 52606 28255 52922 28256
rect 57606 28320 57922 28321
rect 57606 28256 57612 28320
rect 57676 28256 57692 28320
rect 57756 28256 57772 28320
rect 57836 28256 57852 28320
rect 57916 28256 57922 28320
rect 57606 28255 57922 28256
rect 58525 27842 58591 27845
rect 59200 27842 60000 27872
rect 58525 27840 60000 27842
rect 58525 27784 58530 27840
rect 58586 27784 60000 27840
rect 58525 27782 60000 27784
rect 58525 27779 58591 27782
rect 1946 27776 2262 27777
rect 1946 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2262 27776
rect 1946 27711 2262 27712
rect 6946 27776 7262 27777
rect 6946 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7262 27776
rect 6946 27711 7262 27712
rect 11946 27776 12262 27777
rect 11946 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12262 27776
rect 11946 27711 12262 27712
rect 16946 27776 17262 27777
rect 16946 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17262 27776
rect 16946 27711 17262 27712
rect 21946 27776 22262 27777
rect 21946 27712 21952 27776
rect 22016 27712 22032 27776
rect 22096 27712 22112 27776
rect 22176 27712 22192 27776
rect 22256 27712 22262 27776
rect 21946 27711 22262 27712
rect 26946 27776 27262 27777
rect 26946 27712 26952 27776
rect 27016 27712 27032 27776
rect 27096 27712 27112 27776
rect 27176 27712 27192 27776
rect 27256 27712 27262 27776
rect 26946 27711 27262 27712
rect 31946 27776 32262 27777
rect 31946 27712 31952 27776
rect 32016 27712 32032 27776
rect 32096 27712 32112 27776
rect 32176 27712 32192 27776
rect 32256 27712 32262 27776
rect 31946 27711 32262 27712
rect 36946 27776 37262 27777
rect 36946 27712 36952 27776
rect 37016 27712 37032 27776
rect 37096 27712 37112 27776
rect 37176 27712 37192 27776
rect 37256 27712 37262 27776
rect 36946 27711 37262 27712
rect 41946 27776 42262 27777
rect 41946 27712 41952 27776
rect 42016 27712 42032 27776
rect 42096 27712 42112 27776
rect 42176 27712 42192 27776
rect 42256 27712 42262 27776
rect 41946 27711 42262 27712
rect 46946 27776 47262 27777
rect 46946 27712 46952 27776
rect 47016 27712 47032 27776
rect 47096 27712 47112 27776
rect 47176 27712 47192 27776
rect 47256 27712 47262 27776
rect 46946 27711 47262 27712
rect 51946 27776 52262 27777
rect 51946 27712 51952 27776
rect 52016 27712 52032 27776
rect 52096 27712 52112 27776
rect 52176 27712 52192 27776
rect 52256 27712 52262 27776
rect 51946 27711 52262 27712
rect 56946 27776 57262 27777
rect 56946 27712 56952 27776
rect 57016 27712 57032 27776
rect 57096 27712 57112 27776
rect 57176 27712 57192 27776
rect 57256 27712 57262 27776
rect 59200 27752 60000 27782
rect 56946 27711 57262 27712
rect 2606 27232 2922 27233
rect 2606 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2922 27232
rect 2606 27167 2922 27168
rect 7606 27232 7922 27233
rect 7606 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7922 27232
rect 7606 27167 7922 27168
rect 12606 27232 12922 27233
rect 12606 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12922 27232
rect 12606 27167 12922 27168
rect 17606 27232 17922 27233
rect 17606 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17922 27232
rect 17606 27167 17922 27168
rect 22606 27232 22922 27233
rect 22606 27168 22612 27232
rect 22676 27168 22692 27232
rect 22756 27168 22772 27232
rect 22836 27168 22852 27232
rect 22916 27168 22922 27232
rect 22606 27167 22922 27168
rect 27606 27232 27922 27233
rect 27606 27168 27612 27232
rect 27676 27168 27692 27232
rect 27756 27168 27772 27232
rect 27836 27168 27852 27232
rect 27916 27168 27922 27232
rect 27606 27167 27922 27168
rect 32606 27232 32922 27233
rect 32606 27168 32612 27232
rect 32676 27168 32692 27232
rect 32756 27168 32772 27232
rect 32836 27168 32852 27232
rect 32916 27168 32922 27232
rect 32606 27167 32922 27168
rect 37606 27232 37922 27233
rect 37606 27168 37612 27232
rect 37676 27168 37692 27232
rect 37756 27168 37772 27232
rect 37836 27168 37852 27232
rect 37916 27168 37922 27232
rect 37606 27167 37922 27168
rect 42606 27232 42922 27233
rect 42606 27168 42612 27232
rect 42676 27168 42692 27232
rect 42756 27168 42772 27232
rect 42836 27168 42852 27232
rect 42916 27168 42922 27232
rect 42606 27167 42922 27168
rect 47606 27232 47922 27233
rect 47606 27168 47612 27232
rect 47676 27168 47692 27232
rect 47756 27168 47772 27232
rect 47836 27168 47852 27232
rect 47916 27168 47922 27232
rect 47606 27167 47922 27168
rect 52606 27232 52922 27233
rect 52606 27168 52612 27232
rect 52676 27168 52692 27232
rect 52756 27168 52772 27232
rect 52836 27168 52852 27232
rect 52916 27168 52922 27232
rect 52606 27167 52922 27168
rect 57606 27232 57922 27233
rect 57606 27168 57612 27232
rect 57676 27168 57692 27232
rect 57756 27168 57772 27232
rect 57836 27168 57852 27232
rect 57916 27168 57922 27232
rect 57606 27167 57922 27168
rect 58525 27026 58591 27029
rect 59200 27026 60000 27056
rect 58525 27024 60000 27026
rect 58525 26968 58530 27024
rect 58586 26968 60000 27024
rect 58525 26966 60000 26968
rect 58525 26963 58591 26966
rect 59200 26936 60000 26966
rect 1946 26688 2262 26689
rect 1946 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2262 26688
rect 1946 26623 2262 26624
rect 6946 26688 7262 26689
rect 6946 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7262 26688
rect 6946 26623 7262 26624
rect 11946 26688 12262 26689
rect 11946 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12262 26688
rect 11946 26623 12262 26624
rect 16946 26688 17262 26689
rect 16946 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17262 26688
rect 16946 26623 17262 26624
rect 21946 26688 22262 26689
rect 21946 26624 21952 26688
rect 22016 26624 22032 26688
rect 22096 26624 22112 26688
rect 22176 26624 22192 26688
rect 22256 26624 22262 26688
rect 21946 26623 22262 26624
rect 26946 26688 27262 26689
rect 26946 26624 26952 26688
rect 27016 26624 27032 26688
rect 27096 26624 27112 26688
rect 27176 26624 27192 26688
rect 27256 26624 27262 26688
rect 26946 26623 27262 26624
rect 31946 26688 32262 26689
rect 31946 26624 31952 26688
rect 32016 26624 32032 26688
rect 32096 26624 32112 26688
rect 32176 26624 32192 26688
rect 32256 26624 32262 26688
rect 31946 26623 32262 26624
rect 36946 26688 37262 26689
rect 36946 26624 36952 26688
rect 37016 26624 37032 26688
rect 37096 26624 37112 26688
rect 37176 26624 37192 26688
rect 37256 26624 37262 26688
rect 36946 26623 37262 26624
rect 41946 26688 42262 26689
rect 41946 26624 41952 26688
rect 42016 26624 42032 26688
rect 42096 26624 42112 26688
rect 42176 26624 42192 26688
rect 42256 26624 42262 26688
rect 41946 26623 42262 26624
rect 46946 26688 47262 26689
rect 46946 26624 46952 26688
rect 47016 26624 47032 26688
rect 47096 26624 47112 26688
rect 47176 26624 47192 26688
rect 47256 26624 47262 26688
rect 46946 26623 47262 26624
rect 51946 26688 52262 26689
rect 51946 26624 51952 26688
rect 52016 26624 52032 26688
rect 52096 26624 52112 26688
rect 52176 26624 52192 26688
rect 52256 26624 52262 26688
rect 51946 26623 52262 26624
rect 56946 26688 57262 26689
rect 56946 26624 56952 26688
rect 57016 26624 57032 26688
rect 57096 26624 57112 26688
rect 57176 26624 57192 26688
rect 57256 26624 57262 26688
rect 56946 26623 57262 26624
rect 58341 26210 58407 26213
rect 59200 26210 60000 26240
rect 58341 26208 60000 26210
rect 58341 26152 58346 26208
rect 58402 26152 60000 26208
rect 58341 26150 60000 26152
rect 58341 26147 58407 26150
rect 2606 26144 2922 26145
rect 2606 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2922 26144
rect 2606 26079 2922 26080
rect 7606 26144 7922 26145
rect 7606 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7922 26144
rect 7606 26079 7922 26080
rect 12606 26144 12922 26145
rect 12606 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12922 26144
rect 12606 26079 12922 26080
rect 17606 26144 17922 26145
rect 17606 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17922 26144
rect 17606 26079 17922 26080
rect 22606 26144 22922 26145
rect 22606 26080 22612 26144
rect 22676 26080 22692 26144
rect 22756 26080 22772 26144
rect 22836 26080 22852 26144
rect 22916 26080 22922 26144
rect 22606 26079 22922 26080
rect 27606 26144 27922 26145
rect 27606 26080 27612 26144
rect 27676 26080 27692 26144
rect 27756 26080 27772 26144
rect 27836 26080 27852 26144
rect 27916 26080 27922 26144
rect 27606 26079 27922 26080
rect 32606 26144 32922 26145
rect 32606 26080 32612 26144
rect 32676 26080 32692 26144
rect 32756 26080 32772 26144
rect 32836 26080 32852 26144
rect 32916 26080 32922 26144
rect 32606 26079 32922 26080
rect 37606 26144 37922 26145
rect 37606 26080 37612 26144
rect 37676 26080 37692 26144
rect 37756 26080 37772 26144
rect 37836 26080 37852 26144
rect 37916 26080 37922 26144
rect 37606 26079 37922 26080
rect 42606 26144 42922 26145
rect 42606 26080 42612 26144
rect 42676 26080 42692 26144
rect 42756 26080 42772 26144
rect 42836 26080 42852 26144
rect 42916 26080 42922 26144
rect 42606 26079 42922 26080
rect 47606 26144 47922 26145
rect 47606 26080 47612 26144
rect 47676 26080 47692 26144
rect 47756 26080 47772 26144
rect 47836 26080 47852 26144
rect 47916 26080 47922 26144
rect 47606 26079 47922 26080
rect 52606 26144 52922 26145
rect 52606 26080 52612 26144
rect 52676 26080 52692 26144
rect 52756 26080 52772 26144
rect 52836 26080 52852 26144
rect 52916 26080 52922 26144
rect 52606 26079 52922 26080
rect 57606 26144 57922 26145
rect 57606 26080 57612 26144
rect 57676 26080 57692 26144
rect 57756 26080 57772 26144
rect 57836 26080 57852 26144
rect 57916 26080 57922 26144
rect 59200 26120 60000 26150
rect 57606 26079 57922 26080
rect 1946 25600 2262 25601
rect 1946 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2262 25600
rect 1946 25535 2262 25536
rect 6946 25600 7262 25601
rect 6946 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7262 25600
rect 6946 25535 7262 25536
rect 11946 25600 12262 25601
rect 11946 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12262 25600
rect 11946 25535 12262 25536
rect 16946 25600 17262 25601
rect 16946 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17262 25600
rect 16946 25535 17262 25536
rect 21946 25600 22262 25601
rect 21946 25536 21952 25600
rect 22016 25536 22032 25600
rect 22096 25536 22112 25600
rect 22176 25536 22192 25600
rect 22256 25536 22262 25600
rect 21946 25535 22262 25536
rect 26946 25600 27262 25601
rect 26946 25536 26952 25600
rect 27016 25536 27032 25600
rect 27096 25536 27112 25600
rect 27176 25536 27192 25600
rect 27256 25536 27262 25600
rect 26946 25535 27262 25536
rect 31946 25600 32262 25601
rect 31946 25536 31952 25600
rect 32016 25536 32032 25600
rect 32096 25536 32112 25600
rect 32176 25536 32192 25600
rect 32256 25536 32262 25600
rect 31946 25535 32262 25536
rect 36946 25600 37262 25601
rect 36946 25536 36952 25600
rect 37016 25536 37032 25600
rect 37096 25536 37112 25600
rect 37176 25536 37192 25600
rect 37256 25536 37262 25600
rect 36946 25535 37262 25536
rect 41946 25600 42262 25601
rect 41946 25536 41952 25600
rect 42016 25536 42032 25600
rect 42096 25536 42112 25600
rect 42176 25536 42192 25600
rect 42256 25536 42262 25600
rect 41946 25535 42262 25536
rect 46946 25600 47262 25601
rect 46946 25536 46952 25600
rect 47016 25536 47032 25600
rect 47096 25536 47112 25600
rect 47176 25536 47192 25600
rect 47256 25536 47262 25600
rect 46946 25535 47262 25536
rect 51946 25600 52262 25601
rect 51946 25536 51952 25600
rect 52016 25536 52032 25600
rect 52096 25536 52112 25600
rect 52176 25536 52192 25600
rect 52256 25536 52262 25600
rect 51946 25535 52262 25536
rect 56946 25600 57262 25601
rect 56946 25536 56952 25600
rect 57016 25536 57032 25600
rect 57096 25536 57112 25600
rect 57176 25536 57192 25600
rect 57256 25536 57262 25600
rect 56946 25535 57262 25536
rect 58525 25394 58591 25397
rect 59200 25394 60000 25424
rect 58525 25392 60000 25394
rect 58525 25336 58530 25392
rect 58586 25336 60000 25392
rect 58525 25334 60000 25336
rect 58525 25331 58591 25334
rect 59200 25304 60000 25334
rect 2606 25056 2922 25057
rect 2606 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2922 25056
rect 2606 24991 2922 24992
rect 7606 25056 7922 25057
rect 7606 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7922 25056
rect 7606 24991 7922 24992
rect 12606 25056 12922 25057
rect 12606 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12922 25056
rect 12606 24991 12922 24992
rect 17606 25056 17922 25057
rect 17606 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17922 25056
rect 17606 24991 17922 24992
rect 22606 25056 22922 25057
rect 22606 24992 22612 25056
rect 22676 24992 22692 25056
rect 22756 24992 22772 25056
rect 22836 24992 22852 25056
rect 22916 24992 22922 25056
rect 22606 24991 22922 24992
rect 27606 25056 27922 25057
rect 27606 24992 27612 25056
rect 27676 24992 27692 25056
rect 27756 24992 27772 25056
rect 27836 24992 27852 25056
rect 27916 24992 27922 25056
rect 27606 24991 27922 24992
rect 32606 25056 32922 25057
rect 32606 24992 32612 25056
rect 32676 24992 32692 25056
rect 32756 24992 32772 25056
rect 32836 24992 32852 25056
rect 32916 24992 32922 25056
rect 32606 24991 32922 24992
rect 37606 25056 37922 25057
rect 37606 24992 37612 25056
rect 37676 24992 37692 25056
rect 37756 24992 37772 25056
rect 37836 24992 37852 25056
rect 37916 24992 37922 25056
rect 37606 24991 37922 24992
rect 42606 25056 42922 25057
rect 42606 24992 42612 25056
rect 42676 24992 42692 25056
rect 42756 24992 42772 25056
rect 42836 24992 42852 25056
rect 42916 24992 42922 25056
rect 42606 24991 42922 24992
rect 47606 25056 47922 25057
rect 47606 24992 47612 25056
rect 47676 24992 47692 25056
rect 47756 24992 47772 25056
rect 47836 24992 47852 25056
rect 47916 24992 47922 25056
rect 47606 24991 47922 24992
rect 52606 25056 52922 25057
rect 52606 24992 52612 25056
rect 52676 24992 52692 25056
rect 52756 24992 52772 25056
rect 52836 24992 52852 25056
rect 52916 24992 52922 25056
rect 52606 24991 52922 24992
rect 57606 25056 57922 25057
rect 57606 24992 57612 25056
rect 57676 24992 57692 25056
rect 57756 24992 57772 25056
rect 57836 24992 57852 25056
rect 57916 24992 57922 25056
rect 57606 24991 57922 24992
rect 58525 24578 58591 24581
rect 59200 24578 60000 24608
rect 58525 24576 60000 24578
rect 58525 24520 58530 24576
rect 58586 24520 60000 24576
rect 58525 24518 60000 24520
rect 58525 24515 58591 24518
rect 1946 24512 2262 24513
rect 1946 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2262 24512
rect 1946 24447 2262 24448
rect 6946 24512 7262 24513
rect 6946 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7262 24512
rect 6946 24447 7262 24448
rect 11946 24512 12262 24513
rect 11946 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12262 24512
rect 11946 24447 12262 24448
rect 16946 24512 17262 24513
rect 16946 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17262 24512
rect 16946 24447 17262 24448
rect 21946 24512 22262 24513
rect 21946 24448 21952 24512
rect 22016 24448 22032 24512
rect 22096 24448 22112 24512
rect 22176 24448 22192 24512
rect 22256 24448 22262 24512
rect 21946 24447 22262 24448
rect 26946 24512 27262 24513
rect 26946 24448 26952 24512
rect 27016 24448 27032 24512
rect 27096 24448 27112 24512
rect 27176 24448 27192 24512
rect 27256 24448 27262 24512
rect 26946 24447 27262 24448
rect 31946 24512 32262 24513
rect 31946 24448 31952 24512
rect 32016 24448 32032 24512
rect 32096 24448 32112 24512
rect 32176 24448 32192 24512
rect 32256 24448 32262 24512
rect 31946 24447 32262 24448
rect 36946 24512 37262 24513
rect 36946 24448 36952 24512
rect 37016 24448 37032 24512
rect 37096 24448 37112 24512
rect 37176 24448 37192 24512
rect 37256 24448 37262 24512
rect 36946 24447 37262 24448
rect 41946 24512 42262 24513
rect 41946 24448 41952 24512
rect 42016 24448 42032 24512
rect 42096 24448 42112 24512
rect 42176 24448 42192 24512
rect 42256 24448 42262 24512
rect 41946 24447 42262 24448
rect 46946 24512 47262 24513
rect 46946 24448 46952 24512
rect 47016 24448 47032 24512
rect 47096 24448 47112 24512
rect 47176 24448 47192 24512
rect 47256 24448 47262 24512
rect 46946 24447 47262 24448
rect 51946 24512 52262 24513
rect 51946 24448 51952 24512
rect 52016 24448 52032 24512
rect 52096 24448 52112 24512
rect 52176 24448 52192 24512
rect 52256 24448 52262 24512
rect 51946 24447 52262 24448
rect 56946 24512 57262 24513
rect 56946 24448 56952 24512
rect 57016 24448 57032 24512
rect 57096 24448 57112 24512
rect 57176 24448 57192 24512
rect 57256 24448 57262 24512
rect 59200 24488 60000 24518
rect 56946 24447 57262 24448
rect 2606 23968 2922 23969
rect 2606 23904 2612 23968
rect 2676 23904 2692 23968
rect 2756 23904 2772 23968
rect 2836 23904 2852 23968
rect 2916 23904 2922 23968
rect 2606 23903 2922 23904
rect 7606 23968 7922 23969
rect 7606 23904 7612 23968
rect 7676 23904 7692 23968
rect 7756 23904 7772 23968
rect 7836 23904 7852 23968
rect 7916 23904 7922 23968
rect 7606 23903 7922 23904
rect 12606 23968 12922 23969
rect 12606 23904 12612 23968
rect 12676 23904 12692 23968
rect 12756 23904 12772 23968
rect 12836 23904 12852 23968
rect 12916 23904 12922 23968
rect 12606 23903 12922 23904
rect 17606 23968 17922 23969
rect 17606 23904 17612 23968
rect 17676 23904 17692 23968
rect 17756 23904 17772 23968
rect 17836 23904 17852 23968
rect 17916 23904 17922 23968
rect 17606 23903 17922 23904
rect 22606 23968 22922 23969
rect 22606 23904 22612 23968
rect 22676 23904 22692 23968
rect 22756 23904 22772 23968
rect 22836 23904 22852 23968
rect 22916 23904 22922 23968
rect 22606 23903 22922 23904
rect 27606 23968 27922 23969
rect 27606 23904 27612 23968
rect 27676 23904 27692 23968
rect 27756 23904 27772 23968
rect 27836 23904 27852 23968
rect 27916 23904 27922 23968
rect 27606 23903 27922 23904
rect 32606 23968 32922 23969
rect 32606 23904 32612 23968
rect 32676 23904 32692 23968
rect 32756 23904 32772 23968
rect 32836 23904 32852 23968
rect 32916 23904 32922 23968
rect 32606 23903 32922 23904
rect 37606 23968 37922 23969
rect 37606 23904 37612 23968
rect 37676 23904 37692 23968
rect 37756 23904 37772 23968
rect 37836 23904 37852 23968
rect 37916 23904 37922 23968
rect 37606 23903 37922 23904
rect 42606 23968 42922 23969
rect 42606 23904 42612 23968
rect 42676 23904 42692 23968
rect 42756 23904 42772 23968
rect 42836 23904 42852 23968
rect 42916 23904 42922 23968
rect 42606 23903 42922 23904
rect 47606 23968 47922 23969
rect 47606 23904 47612 23968
rect 47676 23904 47692 23968
rect 47756 23904 47772 23968
rect 47836 23904 47852 23968
rect 47916 23904 47922 23968
rect 47606 23903 47922 23904
rect 52606 23968 52922 23969
rect 52606 23904 52612 23968
rect 52676 23904 52692 23968
rect 52756 23904 52772 23968
rect 52836 23904 52852 23968
rect 52916 23904 52922 23968
rect 52606 23903 52922 23904
rect 57606 23968 57922 23969
rect 57606 23904 57612 23968
rect 57676 23904 57692 23968
rect 57756 23904 57772 23968
rect 57836 23904 57852 23968
rect 57916 23904 57922 23968
rect 57606 23903 57922 23904
rect 58525 23762 58591 23765
rect 59200 23762 60000 23792
rect 58525 23760 60000 23762
rect 58525 23704 58530 23760
rect 58586 23704 60000 23760
rect 58525 23702 60000 23704
rect 58525 23699 58591 23702
rect 59200 23672 60000 23702
rect 1946 23424 2262 23425
rect 1946 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2262 23424
rect 1946 23359 2262 23360
rect 6946 23424 7262 23425
rect 6946 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7262 23424
rect 6946 23359 7262 23360
rect 11946 23424 12262 23425
rect 11946 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12262 23424
rect 11946 23359 12262 23360
rect 16946 23424 17262 23425
rect 16946 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17262 23424
rect 16946 23359 17262 23360
rect 21946 23424 22262 23425
rect 21946 23360 21952 23424
rect 22016 23360 22032 23424
rect 22096 23360 22112 23424
rect 22176 23360 22192 23424
rect 22256 23360 22262 23424
rect 21946 23359 22262 23360
rect 26946 23424 27262 23425
rect 26946 23360 26952 23424
rect 27016 23360 27032 23424
rect 27096 23360 27112 23424
rect 27176 23360 27192 23424
rect 27256 23360 27262 23424
rect 26946 23359 27262 23360
rect 31946 23424 32262 23425
rect 31946 23360 31952 23424
rect 32016 23360 32032 23424
rect 32096 23360 32112 23424
rect 32176 23360 32192 23424
rect 32256 23360 32262 23424
rect 31946 23359 32262 23360
rect 36946 23424 37262 23425
rect 36946 23360 36952 23424
rect 37016 23360 37032 23424
rect 37096 23360 37112 23424
rect 37176 23360 37192 23424
rect 37256 23360 37262 23424
rect 36946 23359 37262 23360
rect 41946 23424 42262 23425
rect 41946 23360 41952 23424
rect 42016 23360 42032 23424
rect 42096 23360 42112 23424
rect 42176 23360 42192 23424
rect 42256 23360 42262 23424
rect 41946 23359 42262 23360
rect 46946 23424 47262 23425
rect 46946 23360 46952 23424
rect 47016 23360 47032 23424
rect 47096 23360 47112 23424
rect 47176 23360 47192 23424
rect 47256 23360 47262 23424
rect 46946 23359 47262 23360
rect 51946 23424 52262 23425
rect 51946 23360 51952 23424
rect 52016 23360 52032 23424
rect 52096 23360 52112 23424
rect 52176 23360 52192 23424
rect 52256 23360 52262 23424
rect 51946 23359 52262 23360
rect 56946 23424 57262 23425
rect 56946 23360 56952 23424
rect 57016 23360 57032 23424
rect 57096 23360 57112 23424
rect 57176 23360 57192 23424
rect 57256 23360 57262 23424
rect 56946 23359 57262 23360
rect 58525 22946 58591 22949
rect 59200 22946 60000 22976
rect 58525 22944 60000 22946
rect 58525 22888 58530 22944
rect 58586 22888 60000 22944
rect 58525 22886 60000 22888
rect 58525 22883 58591 22886
rect 2606 22880 2922 22881
rect 2606 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2922 22880
rect 2606 22815 2922 22816
rect 7606 22880 7922 22881
rect 7606 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7922 22880
rect 7606 22815 7922 22816
rect 12606 22880 12922 22881
rect 12606 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12922 22880
rect 12606 22815 12922 22816
rect 17606 22880 17922 22881
rect 17606 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17922 22880
rect 17606 22815 17922 22816
rect 22606 22880 22922 22881
rect 22606 22816 22612 22880
rect 22676 22816 22692 22880
rect 22756 22816 22772 22880
rect 22836 22816 22852 22880
rect 22916 22816 22922 22880
rect 22606 22815 22922 22816
rect 27606 22880 27922 22881
rect 27606 22816 27612 22880
rect 27676 22816 27692 22880
rect 27756 22816 27772 22880
rect 27836 22816 27852 22880
rect 27916 22816 27922 22880
rect 27606 22815 27922 22816
rect 32606 22880 32922 22881
rect 32606 22816 32612 22880
rect 32676 22816 32692 22880
rect 32756 22816 32772 22880
rect 32836 22816 32852 22880
rect 32916 22816 32922 22880
rect 32606 22815 32922 22816
rect 37606 22880 37922 22881
rect 37606 22816 37612 22880
rect 37676 22816 37692 22880
rect 37756 22816 37772 22880
rect 37836 22816 37852 22880
rect 37916 22816 37922 22880
rect 37606 22815 37922 22816
rect 42606 22880 42922 22881
rect 42606 22816 42612 22880
rect 42676 22816 42692 22880
rect 42756 22816 42772 22880
rect 42836 22816 42852 22880
rect 42916 22816 42922 22880
rect 42606 22815 42922 22816
rect 47606 22880 47922 22881
rect 47606 22816 47612 22880
rect 47676 22816 47692 22880
rect 47756 22816 47772 22880
rect 47836 22816 47852 22880
rect 47916 22816 47922 22880
rect 47606 22815 47922 22816
rect 52606 22880 52922 22881
rect 52606 22816 52612 22880
rect 52676 22816 52692 22880
rect 52756 22816 52772 22880
rect 52836 22816 52852 22880
rect 52916 22816 52922 22880
rect 52606 22815 52922 22816
rect 57606 22880 57922 22881
rect 57606 22816 57612 22880
rect 57676 22816 57692 22880
rect 57756 22816 57772 22880
rect 57836 22816 57852 22880
rect 57916 22816 57922 22880
rect 59200 22856 60000 22886
rect 57606 22815 57922 22816
rect 1946 22336 2262 22337
rect 1946 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2262 22336
rect 1946 22271 2262 22272
rect 6946 22336 7262 22337
rect 6946 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7262 22336
rect 6946 22271 7262 22272
rect 11946 22336 12262 22337
rect 11946 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12262 22336
rect 11946 22271 12262 22272
rect 16946 22336 17262 22337
rect 16946 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17262 22336
rect 16946 22271 17262 22272
rect 21946 22336 22262 22337
rect 21946 22272 21952 22336
rect 22016 22272 22032 22336
rect 22096 22272 22112 22336
rect 22176 22272 22192 22336
rect 22256 22272 22262 22336
rect 21946 22271 22262 22272
rect 26946 22336 27262 22337
rect 26946 22272 26952 22336
rect 27016 22272 27032 22336
rect 27096 22272 27112 22336
rect 27176 22272 27192 22336
rect 27256 22272 27262 22336
rect 26946 22271 27262 22272
rect 31946 22336 32262 22337
rect 31946 22272 31952 22336
rect 32016 22272 32032 22336
rect 32096 22272 32112 22336
rect 32176 22272 32192 22336
rect 32256 22272 32262 22336
rect 31946 22271 32262 22272
rect 36946 22336 37262 22337
rect 36946 22272 36952 22336
rect 37016 22272 37032 22336
rect 37096 22272 37112 22336
rect 37176 22272 37192 22336
rect 37256 22272 37262 22336
rect 36946 22271 37262 22272
rect 41946 22336 42262 22337
rect 41946 22272 41952 22336
rect 42016 22272 42032 22336
rect 42096 22272 42112 22336
rect 42176 22272 42192 22336
rect 42256 22272 42262 22336
rect 41946 22271 42262 22272
rect 46946 22336 47262 22337
rect 46946 22272 46952 22336
rect 47016 22272 47032 22336
rect 47096 22272 47112 22336
rect 47176 22272 47192 22336
rect 47256 22272 47262 22336
rect 46946 22271 47262 22272
rect 51946 22336 52262 22337
rect 51946 22272 51952 22336
rect 52016 22272 52032 22336
rect 52096 22272 52112 22336
rect 52176 22272 52192 22336
rect 52256 22272 52262 22336
rect 51946 22271 52262 22272
rect 56946 22336 57262 22337
rect 56946 22272 56952 22336
rect 57016 22272 57032 22336
rect 57096 22272 57112 22336
rect 57176 22272 57192 22336
rect 57256 22272 57262 22336
rect 56946 22271 57262 22272
rect 58525 22130 58591 22133
rect 59200 22130 60000 22160
rect 58525 22128 60000 22130
rect 58525 22072 58530 22128
rect 58586 22072 60000 22128
rect 58525 22070 60000 22072
rect 58525 22067 58591 22070
rect 59200 22040 60000 22070
rect 2606 21792 2922 21793
rect 2606 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2922 21792
rect 2606 21727 2922 21728
rect 7606 21792 7922 21793
rect 7606 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7922 21792
rect 7606 21727 7922 21728
rect 12606 21792 12922 21793
rect 12606 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12922 21792
rect 12606 21727 12922 21728
rect 17606 21792 17922 21793
rect 17606 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17922 21792
rect 17606 21727 17922 21728
rect 22606 21792 22922 21793
rect 22606 21728 22612 21792
rect 22676 21728 22692 21792
rect 22756 21728 22772 21792
rect 22836 21728 22852 21792
rect 22916 21728 22922 21792
rect 22606 21727 22922 21728
rect 27606 21792 27922 21793
rect 27606 21728 27612 21792
rect 27676 21728 27692 21792
rect 27756 21728 27772 21792
rect 27836 21728 27852 21792
rect 27916 21728 27922 21792
rect 27606 21727 27922 21728
rect 32606 21792 32922 21793
rect 32606 21728 32612 21792
rect 32676 21728 32692 21792
rect 32756 21728 32772 21792
rect 32836 21728 32852 21792
rect 32916 21728 32922 21792
rect 32606 21727 32922 21728
rect 37606 21792 37922 21793
rect 37606 21728 37612 21792
rect 37676 21728 37692 21792
rect 37756 21728 37772 21792
rect 37836 21728 37852 21792
rect 37916 21728 37922 21792
rect 37606 21727 37922 21728
rect 42606 21792 42922 21793
rect 42606 21728 42612 21792
rect 42676 21728 42692 21792
rect 42756 21728 42772 21792
rect 42836 21728 42852 21792
rect 42916 21728 42922 21792
rect 42606 21727 42922 21728
rect 47606 21792 47922 21793
rect 47606 21728 47612 21792
rect 47676 21728 47692 21792
rect 47756 21728 47772 21792
rect 47836 21728 47852 21792
rect 47916 21728 47922 21792
rect 47606 21727 47922 21728
rect 52606 21792 52922 21793
rect 52606 21728 52612 21792
rect 52676 21728 52692 21792
rect 52756 21728 52772 21792
rect 52836 21728 52852 21792
rect 52916 21728 52922 21792
rect 52606 21727 52922 21728
rect 57606 21792 57922 21793
rect 57606 21728 57612 21792
rect 57676 21728 57692 21792
rect 57756 21728 57772 21792
rect 57836 21728 57852 21792
rect 57916 21728 57922 21792
rect 57606 21727 57922 21728
rect 58525 21314 58591 21317
rect 59200 21314 60000 21344
rect 58525 21312 60000 21314
rect 58525 21256 58530 21312
rect 58586 21256 60000 21312
rect 58525 21254 60000 21256
rect 58525 21251 58591 21254
rect 1946 21248 2262 21249
rect 1946 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2262 21248
rect 1946 21183 2262 21184
rect 6946 21248 7262 21249
rect 6946 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7262 21248
rect 6946 21183 7262 21184
rect 11946 21248 12262 21249
rect 11946 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12262 21248
rect 11946 21183 12262 21184
rect 16946 21248 17262 21249
rect 16946 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17262 21248
rect 16946 21183 17262 21184
rect 21946 21248 22262 21249
rect 21946 21184 21952 21248
rect 22016 21184 22032 21248
rect 22096 21184 22112 21248
rect 22176 21184 22192 21248
rect 22256 21184 22262 21248
rect 21946 21183 22262 21184
rect 26946 21248 27262 21249
rect 26946 21184 26952 21248
rect 27016 21184 27032 21248
rect 27096 21184 27112 21248
rect 27176 21184 27192 21248
rect 27256 21184 27262 21248
rect 26946 21183 27262 21184
rect 31946 21248 32262 21249
rect 31946 21184 31952 21248
rect 32016 21184 32032 21248
rect 32096 21184 32112 21248
rect 32176 21184 32192 21248
rect 32256 21184 32262 21248
rect 31946 21183 32262 21184
rect 36946 21248 37262 21249
rect 36946 21184 36952 21248
rect 37016 21184 37032 21248
rect 37096 21184 37112 21248
rect 37176 21184 37192 21248
rect 37256 21184 37262 21248
rect 36946 21183 37262 21184
rect 41946 21248 42262 21249
rect 41946 21184 41952 21248
rect 42016 21184 42032 21248
rect 42096 21184 42112 21248
rect 42176 21184 42192 21248
rect 42256 21184 42262 21248
rect 41946 21183 42262 21184
rect 46946 21248 47262 21249
rect 46946 21184 46952 21248
rect 47016 21184 47032 21248
rect 47096 21184 47112 21248
rect 47176 21184 47192 21248
rect 47256 21184 47262 21248
rect 46946 21183 47262 21184
rect 51946 21248 52262 21249
rect 51946 21184 51952 21248
rect 52016 21184 52032 21248
rect 52096 21184 52112 21248
rect 52176 21184 52192 21248
rect 52256 21184 52262 21248
rect 51946 21183 52262 21184
rect 56946 21248 57262 21249
rect 56946 21184 56952 21248
rect 57016 21184 57032 21248
rect 57096 21184 57112 21248
rect 57176 21184 57192 21248
rect 57256 21184 57262 21248
rect 59200 21224 60000 21254
rect 56946 21183 57262 21184
rect 2606 20704 2922 20705
rect 2606 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2922 20704
rect 2606 20639 2922 20640
rect 7606 20704 7922 20705
rect 7606 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7922 20704
rect 7606 20639 7922 20640
rect 12606 20704 12922 20705
rect 12606 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12922 20704
rect 12606 20639 12922 20640
rect 17606 20704 17922 20705
rect 17606 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17922 20704
rect 17606 20639 17922 20640
rect 22606 20704 22922 20705
rect 22606 20640 22612 20704
rect 22676 20640 22692 20704
rect 22756 20640 22772 20704
rect 22836 20640 22852 20704
rect 22916 20640 22922 20704
rect 22606 20639 22922 20640
rect 27606 20704 27922 20705
rect 27606 20640 27612 20704
rect 27676 20640 27692 20704
rect 27756 20640 27772 20704
rect 27836 20640 27852 20704
rect 27916 20640 27922 20704
rect 27606 20639 27922 20640
rect 32606 20704 32922 20705
rect 32606 20640 32612 20704
rect 32676 20640 32692 20704
rect 32756 20640 32772 20704
rect 32836 20640 32852 20704
rect 32916 20640 32922 20704
rect 32606 20639 32922 20640
rect 37606 20704 37922 20705
rect 37606 20640 37612 20704
rect 37676 20640 37692 20704
rect 37756 20640 37772 20704
rect 37836 20640 37852 20704
rect 37916 20640 37922 20704
rect 37606 20639 37922 20640
rect 42606 20704 42922 20705
rect 42606 20640 42612 20704
rect 42676 20640 42692 20704
rect 42756 20640 42772 20704
rect 42836 20640 42852 20704
rect 42916 20640 42922 20704
rect 42606 20639 42922 20640
rect 47606 20704 47922 20705
rect 47606 20640 47612 20704
rect 47676 20640 47692 20704
rect 47756 20640 47772 20704
rect 47836 20640 47852 20704
rect 47916 20640 47922 20704
rect 47606 20639 47922 20640
rect 52606 20704 52922 20705
rect 52606 20640 52612 20704
rect 52676 20640 52692 20704
rect 52756 20640 52772 20704
rect 52836 20640 52852 20704
rect 52916 20640 52922 20704
rect 52606 20639 52922 20640
rect 57606 20704 57922 20705
rect 57606 20640 57612 20704
rect 57676 20640 57692 20704
rect 57756 20640 57772 20704
rect 57836 20640 57852 20704
rect 57916 20640 57922 20704
rect 57606 20639 57922 20640
rect 58525 20498 58591 20501
rect 59200 20498 60000 20528
rect 58525 20496 60000 20498
rect 58525 20440 58530 20496
rect 58586 20440 60000 20496
rect 58525 20438 60000 20440
rect 58525 20435 58591 20438
rect 59200 20408 60000 20438
rect 1946 20160 2262 20161
rect 1946 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2262 20160
rect 1946 20095 2262 20096
rect 6946 20160 7262 20161
rect 6946 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7262 20160
rect 6946 20095 7262 20096
rect 11946 20160 12262 20161
rect 11946 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12262 20160
rect 11946 20095 12262 20096
rect 16946 20160 17262 20161
rect 16946 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17262 20160
rect 16946 20095 17262 20096
rect 21946 20160 22262 20161
rect 21946 20096 21952 20160
rect 22016 20096 22032 20160
rect 22096 20096 22112 20160
rect 22176 20096 22192 20160
rect 22256 20096 22262 20160
rect 21946 20095 22262 20096
rect 26946 20160 27262 20161
rect 26946 20096 26952 20160
rect 27016 20096 27032 20160
rect 27096 20096 27112 20160
rect 27176 20096 27192 20160
rect 27256 20096 27262 20160
rect 26946 20095 27262 20096
rect 31946 20160 32262 20161
rect 31946 20096 31952 20160
rect 32016 20096 32032 20160
rect 32096 20096 32112 20160
rect 32176 20096 32192 20160
rect 32256 20096 32262 20160
rect 31946 20095 32262 20096
rect 36946 20160 37262 20161
rect 36946 20096 36952 20160
rect 37016 20096 37032 20160
rect 37096 20096 37112 20160
rect 37176 20096 37192 20160
rect 37256 20096 37262 20160
rect 36946 20095 37262 20096
rect 41946 20160 42262 20161
rect 41946 20096 41952 20160
rect 42016 20096 42032 20160
rect 42096 20096 42112 20160
rect 42176 20096 42192 20160
rect 42256 20096 42262 20160
rect 41946 20095 42262 20096
rect 46946 20160 47262 20161
rect 46946 20096 46952 20160
rect 47016 20096 47032 20160
rect 47096 20096 47112 20160
rect 47176 20096 47192 20160
rect 47256 20096 47262 20160
rect 46946 20095 47262 20096
rect 51946 20160 52262 20161
rect 51946 20096 51952 20160
rect 52016 20096 52032 20160
rect 52096 20096 52112 20160
rect 52176 20096 52192 20160
rect 52256 20096 52262 20160
rect 51946 20095 52262 20096
rect 56946 20160 57262 20161
rect 56946 20096 56952 20160
rect 57016 20096 57032 20160
rect 57096 20096 57112 20160
rect 57176 20096 57192 20160
rect 57256 20096 57262 20160
rect 56946 20095 57262 20096
rect 58525 19682 58591 19685
rect 59200 19682 60000 19712
rect 58525 19680 60000 19682
rect 58525 19624 58530 19680
rect 58586 19624 60000 19680
rect 58525 19622 60000 19624
rect 58525 19619 58591 19622
rect 2606 19616 2922 19617
rect 2606 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2922 19616
rect 2606 19551 2922 19552
rect 7606 19616 7922 19617
rect 7606 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7922 19616
rect 7606 19551 7922 19552
rect 12606 19616 12922 19617
rect 12606 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12922 19616
rect 12606 19551 12922 19552
rect 17606 19616 17922 19617
rect 17606 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17922 19616
rect 17606 19551 17922 19552
rect 22606 19616 22922 19617
rect 22606 19552 22612 19616
rect 22676 19552 22692 19616
rect 22756 19552 22772 19616
rect 22836 19552 22852 19616
rect 22916 19552 22922 19616
rect 22606 19551 22922 19552
rect 27606 19616 27922 19617
rect 27606 19552 27612 19616
rect 27676 19552 27692 19616
rect 27756 19552 27772 19616
rect 27836 19552 27852 19616
rect 27916 19552 27922 19616
rect 27606 19551 27922 19552
rect 32606 19616 32922 19617
rect 32606 19552 32612 19616
rect 32676 19552 32692 19616
rect 32756 19552 32772 19616
rect 32836 19552 32852 19616
rect 32916 19552 32922 19616
rect 32606 19551 32922 19552
rect 37606 19616 37922 19617
rect 37606 19552 37612 19616
rect 37676 19552 37692 19616
rect 37756 19552 37772 19616
rect 37836 19552 37852 19616
rect 37916 19552 37922 19616
rect 37606 19551 37922 19552
rect 42606 19616 42922 19617
rect 42606 19552 42612 19616
rect 42676 19552 42692 19616
rect 42756 19552 42772 19616
rect 42836 19552 42852 19616
rect 42916 19552 42922 19616
rect 42606 19551 42922 19552
rect 47606 19616 47922 19617
rect 47606 19552 47612 19616
rect 47676 19552 47692 19616
rect 47756 19552 47772 19616
rect 47836 19552 47852 19616
rect 47916 19552 47922 19616
rect 47606 19551 47922 19552
rect 52606 19616 52922 19617
rect 52606 19552 52612 19616
rect 52676 19552 52692 19616
rect 52756 19552 52772 19616
rect 52836 19552 52852 19616
rect 52916 19552 52922 19616
rect 52606 19551 52922 19552
rect 57606 19616 57922 19617
rect 57606 19552 57612 19616
rect 57676 19552 57692 19616
rect 57756 19552 57772 19616
rect 57836 19552 57852 19616
rect 57916 19552 57922 19616
rect 59200 19592 60000 19622
rect 57606 19551 57922 19552
rect 1946 19072 2262 19073
rect 1946 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2262 19072
rect 1946 19007 2262 19008
rect 6946 19072 7262 19073
rect 6946 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7262 19072
rect 6946 19007 7262 19008
rect 11946 19072 12262 19073
rect 11946 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12262 19072
rect 11946 19007 12262 19008
rect 16946 19072 17262 19073
rect 16946 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17262 19072
rect 16946 19007 17262 19008
rect 21946 19072 22262 19073
rect 21946 19008 21952 19072
rect 22016 19008 22032 19072
rect 22096 19008 22112 19072
rect 22176 19008 22192 19072
rect 22256 19008 22262 19072
rect 21946 19007 22262 19008
rect 26946 19072 27262 19073
rect 26946 19008 26952 19072
rect 27016 19008 27032 19072
rect 27096 19008 27112 19072
rect 27176 19008 27192 19072
rect 27256 19008 27262 19072
rect 26946 19007 27262 19008
rect 31946 19072 32262 19073
rect 31946 19008 31952 19072
rect 32016 19008 32032 19072
rect 32096 19008 32112 19072
rect 32176 19008 32192 19072
rect 32256 19008 32262 19072
rect 31946 19007 32262 19008
rect 36946 19072 37262 19073
rect 36946 19008 36952 19072
rect 37016 19008 37032 19072
rect 37096 19008 37112 19072
rect 37176 19008 37192 19072
rect 37256 19008 37262 19072
rect 36946 19007 37262 19008
rect 41946 19072 42262 19073
rect 41946 19008 41952 19072
rect 42016 19008 42032 19072
rect 42096 19008 42112 19072
rect 42176 19008 42192 19072
rect 42256 19008 42262 19072
rect 41946 19007 42262 19008
rect 46946 19072 47262 19073
rect 46946 19008 46952 19072
rect 47016 19008 47032 19072
rect 47096 19008 47112 19072
rect 47176 19008 47192 19072
rect 47256 19008 47262 19072
rect 46946 19007 47262 19008
rect 51946 19072 52262 19073
rect 51946 19008 51952 19072
rect 52016 19008 52032 19072
rect 52096 19008 52112 19072
rect 52176 19008 52192 19072
rect 52256 19008 52262 19072
rect 51946 19007 52262 19008
rect 56946 19072 57262 19073
rect 56946 19008 56952 19072
rect 57016 19008 57032 19072
rect 57096 19008 57112 19072
rect 57176 19008 57192 19072
rect 57256 19008 57262 19072
rect 56946 19007 57262 19008
rect 58525 18866 58591 18869
rect 59200 18866 60000 18896
rect 58525 18864 60000 18866
rect 58525 18808 58530 18864
rect 58586 18808 60000 18864
rect 58525 18806 60000 18808
rect 58525 18803 58591 18806
rect 59200 18776 60000 18806
rect 2606 18528 2922 18529
rect 2606 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2922 18528
rect 2606 18463 2922 18464
rect 7606 18528 7922 18529
rect 7606 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7922 18528
rect 7606 18463 7922 18464
rect 12606 18528 12922 18529
rect 12606 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12922 18528
rect 12606 18463 12922 18464
rect 17606 18528 17922 18529
rect 17606 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17922 18528
rect 17606 18463 17922 18464
rect 22606 18528 22922 18529
rect 22606 18464 22612 18528
rect 22676 18464 22692 18528
rect 22756 18464 22772 18528
rect 22836 18464 22852 18528
rect 22916 18464 22922 18528
rect 22606 18463 22922 18464
rect 27606 18528 27922 18529
rect 27606 18464 27612 18528
rect 27676 18464 27692 18528
rect 27756 18464 27772 18528
rect 27836 18464 27852 18528
rect 27916 18464 27922 18528
rect 27606 18463 27922 18464
rect 32606 18528 32922 18529
rect 32606 18464 32612 18528
rect 32676 18464 32692 18528
rect 32756 18464 32772 18528
rect 32836 18464 32852 18528
rect 32916 18464 32922 18528
rect 32606 18463 32922 18464
rect 37606 18528 37922 18529
rect 37606 18464 37612 18528
rect 37676 18464 37692 18528
rect 37756 18464 37772 18528
rect 37836 18464 37852 18528
rect 37916 18464 37922 18528
rect 37606 18463 37922 18464
rect 42606 18528 42922 18529
rect 42606 18464 42612 18528
rect 42676 18464 42692 18528
rect 42756 18464 42772 18528
rect 42836 18464 42852 18528
rect 42916 18464 42922 18528
rect 42606 18463 42922 18464
rect 47606 18528 47922 18529
rect 47606 18464 47612 18528
rect 47676 18464 47692 18528
rect 47756 18464 47772 18528
rect 47836 18464 47852 18528
rect 47916 18464 47922 18528
rect 47606 18463 47922 18464
rect 52606 18528 52922 18529
rect 52606 18464 52612 18528
rect 52676 18464 52692 18528
rect 52756 18464 52772 18528
rect 52836 18464 52852 18528
rect 52916 18464 52922 18528
rect 52606 18463 52922 18464
rect 57606 18528 57922 18529
rect 57606 18464 57612 18528
rect 57676 18464 57692 18528
rect 57756 18464 57772 18528
rect 57836 18464 57852 18528
rect 57916 18464 57922 18528
rect 57606 18463 57922 18464
rect 58525 18050 58591 18053
rect 59200 18050 60000 18080
rect 58525 18048 60000 18050
rect 58525 17992 58530 18048
rect 58586 17992 60000 18048
rect 58525 17990 60000 17992
rect 58525 17987 58591 17990
rect 1946 17984 2262 17985
rect 1946 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2262 17984
rect 1946 17919 2262 17920
rect 6946 17984 7262 17985
rect 6946 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7262 17984
rect 6946 17919 7262 17920
rect 11946 17984 12262 17985
rect 11946 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12262 17984
rect 11946 17919 12262 17920
rect 16946 17984 17262 17985
rect 16946 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17262 17984
rect 16946 17919 17262 17920
rect 21946 17984 22262 17985
rect 21946 17920 21952 17984
rect 22016 17920 22032 17984
rect 22096 17920 22112 17984
rect 22176 17920 22192 17984
rect 22256 17920 22262 17984
rect 21946 17919 22262 17920
rect 26946 17984 27262 17985
rect 26946 17920 26952 17984
rect 27016 17920 27032 17984
rect 27096 17920 27112 17984
rect 27176 17920 27192 17984
rect 27256 17920 27262 17984
rect 26946 17919 27262 17920
rect 31946 17984 32262 17985
rect 31946 17920 31952 17984
rect 32016 17920 32032 17984
rect 32096 17920 32112 17984
rect 32176 17920 32192 17984
rect 32256 17920 32262 17984
rect 31946 17919 32262 17920
rect 36946 17984 37262 17985
rect 36946 17920 36952 17984
rect 37016 17920 37032 17984
rect 37096 17920 37112 17984
rect 37176 17920 37192 17984
rect 37256 17920 37262 17984
rect 36946 17919 37262 17920
rect 41946 17984 42262 17985
rect 41946 17920 41952 17984
rect 42016 17920 42032 17984
rect 42096 17920 42112 17984
rect 42176 17920 42192 17984
rect 42256 17920 42262 17984
rect 41946 17919 42262 17920
rect 46946 17984 47262 17985
rect 46946 17920 46952 17984
rect 47016 17920 47032 17984
rect 47096 17920 47112 17984
rect 47176 17920 47192 17984
rect 47256 17920 47262 17984
rect 46946 17919 47262 17920
rect 51946 17984 52262 17985
rect 51946 17920 51952 17984
rect 52016 17920 52032 17984
rect 52096 17920 52112 17984
rect 52176 17920 52192 17984
rect 52256 17920 52262 17984
rect 51946 17919 52262 17920
rect 56946 17984 57262 17985
rect 56946 17920 56952 17984
rect 57016 17920 57032 17984
rect 57096 17920 57112 17984
rect 57176 17920 57192 17984
rect 57256 17920 57262 17984
rect 59200 17960 60000 17990
rect 56946 17919 57262 17920
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 17606 17375 17922 17376
rect 22606 17440 22922 17441
rect 22606 17376 22612 17440
rect 22676 17376 22692 17440
rect 22756 17376 22772 17440
rect 22836 17376 22852 17440
rect 22916 17376 22922 17440
rect 22606 17375 22922 17376
rect 27606 17440 27922 17441
rect 27606 17376 27612 17440
rect 27676 17376 27692 17440
rect 27756 17376 27772 17440
rect 27836 17376 27852 17440
rect 27916 17376 27922 17440
rect 27606 17375 27922 17376
rect 32606 17440 32922 17441
rect 32606 17376 32612 17440
rect 32676 17376 32692 17440
rect 32756 17376 32772 17440
rect 32836 17376 32852 17440
rect 32916 17376 32922 17440
rect 32606 17375 32922 17376
rect 37606 17440 37922 17441
rect 37606 17376 37612 17440
rect 37676 17376 37692 17440
rect 37756 17376 37772 17440
rect 37836 17376 37852 17440
rect 37916 17376 37922 17440
rect 37606 17375 37922 17376
rect 42606 17440 42922 17441
rect 42606 17376 42612 17440
rect 42676 17376 42692 17440
rect 42756 17376 42772 17440
rect 42836 17376 42852 17440
rect 42916 17376 42922 17440
rect 42606 17375 42922 17376
rect 47606 17440 47922 17441
rect 47606 17376 47612 17440
rect 47676 17376 47692 17440
rect 47756 17376 47772 17440
rect 47836 17376 47852 17440
rect 47916 17376 47922 17440
rect 47606 17375 47922 17376
rect 52606 17440 52922 17441
rect 52606 17376 52612 17440
rect 52676 17376 52692 17440
rect 52756 17376 52772 17440
rect 52836 17376 52852 17440
rect 52916 17376 52922 17440
rect 52606 17375 52922 17376
rect 57606 17440 57922 17441
rect 57606 17376 57612 17440
rect 57676 17376 57692 17440
rect 57756 17376 57772 17440
rect 57836 17376 57852 17440
rect 57916 17376 57922 17440
rect 57606 17375 57922 17376
rect 58525 17234 58591 17237
rect 59200 17234 60000 17264
rect 58525 17232 60000 17234
rect 58525 17176 58530 17232
rect 58586 17176 60000 17232
rect 58525 17174 60000 17176
rect 58525 17171 58591 17174
rect 59200 17144 60000 17174
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 21946 16896 22262 16897
rect 21946 16832 21952 16896
rect 22016 16832 22032 16896
rect 22096 16832 22112 16896
rect 22176 16832 22192 16896
rect 22256 16832 22262 16896
rect 21946 16831 22262 16832
rect 26946 16896 27262 16897
rect 26946 16832 26952 16896
rect 27016 16832 27032 16896
rect 27096 16832 27112 16896
rect 27176 16832 27192 16896
rect 27256 16832 27262 16896
rect 26946 16831 27262 16832
rect 31946 16896 32262 16897
rect 31946 16832 31952 16896
rect 32016 16832 32032 16896
rect 32096 16832 32112 16896
rect 32176 16832 32192 16896
rect 32256 16832 32262 16896
rect 31946 16831 32262 16832
rect 36946 16896 37262 16897
rect 36946 16832 36952 16896
rect 37016 16832 37032 16896
rect 37096 16832 37112 16896
rect 37176 16832 37192 16896
rect 37256 16832 37262 16896
rect 36946 16831 37262 16832
rect 41946 16896 42262 16897
rect 41946 16832 41952 16896
rect 42016 16832 42032 16896
rect 42096 16832 42112 16896
rect 42176 16832 42192 16896
rect 42256 16832 42262 16896
rect 41946 16831 42262 16832
rect 46946 16896 47262 16897
rect 46946 16832 46952 16896
rect 47016 16832 47032 16896
rect 47096 16832 47112 16896
rect 47176 16832 47192 16896
rect 47256 16832 47262 16896
rect 46946 16831 47262 16832
rect 51946 16896 52262 16897
rect 51946 16832 51952 16896
rect 52016 16832 52032 16896
rect 52096 16832 52112 16896
rect 52176 16832 52192 16896
rect 52256 16832 52262 16896
rect 51946 16831 52262 16832
rect 56946 16896 57262 16897
rect 56946 16832 56952 16896
rect 57016 16832 57032 16896
rect 57096 16832 57112 16896
rect 57176 16832 57192 16896
rect 57256 16832 57262 16896
rect 56946 16831 57262 16832
rect 57881 16554 57947 16557
rect 57881 16552 58082 16554
rect 57881 16496 57886 16552
rect 57942 16496 58082 16552
rect 57881 16494 58082 16496
rect 57881 16491 57947 16494
rect 58022 16418 58082 16494
rect 59200 16418 60000 16448
rect 58022 16358 60000 16418
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 17606 16287 17922 16288
rect 22606 16352 22922 16353
rect 22606 16288 22612 16352
rect 22676 16288 22692 16352
rect 22756 16288 22772 16352
rect 22836 16288 22852 16352
rect 22916 16288 22922 16352
rect 22606 16287 22922 16288
rect 27606 16352 27922 16353
rect 27606 16288 27612 16352
rect 27676 16288 27692 16352
rect 27756 16288 27772 16352
rect 27836 16288 27852 16352
rect 27916 16288 27922 16352
rect 27606 16287 27922 16288
rect 32606 16352 32922 16353
rect 32606 16288 32612 16352
rect 32676 16288 32692 16352
rect 32756 16288 32772 16352
rect 32836 16288 32852 16352
rect 32916 16288 32922 16352
rect 32606 16287 32922 16288
rect 37606 16352 37922 16353
rect 37606 16288 37612 16352
rect 37676 16288 37692 16352
rect 37756 16288 37772 16352
rect 37836 16288 37852 16352
rect 37916 16288 37922 16352
rect 37606 16287 37922 16288
rect 42606 16352 42922 16353
rect 42606 16288 42612 16352
rect 42676 16288 42692 16352
rect 42756 16288 42772 16352
rect 42836 16288 42852 16352
rect 42916 16288 42922 16352
rect 42606 16287 42922 16288
rect 47606 16352 47922 16353
rect 47606 16288 47612 16352
rect 47676 16288 47692 16352
rect 47756 16288 47772 16352
rect 47836 16288 47852 16352
rect 47916 16288 47922 16352
rect 47606 16287 47922 16288
rect 52606 16352 52922 16353
rect 52606 16288 52612 16352
rect 52676 16288 52692 16352
rect 52756 16288 52772 16352
rect 52836 16288 52852 16352
rect 52916 16288 52922 16352
rect 52606 16287 52922 16288
rect 57606 16352 57922 16353
rect 57606 16288 57612 16352
rect 57676 16288 57692 16352
rect 57756 16288 57772 16352
rect 57836 16288 57852 16352
rect 57916 16288 57922 16352
rect 59200 16328 60000 16358
rect 57606 16287 57922 16288
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 21946 15808 22262 15809
rect 21946 15744 21952 15808
rect 22016 15744 22032 15808
rect 22096 15744 22112 15808
rect 22176 15744 22192 15808
rect 22256 15744 22262 15808
rect 21946 15743 22262 15744
rect 26946 15808 27262 15809
rect 26946 15744 26952 15808
rect 27016 15744 27032 15808
rect 27096 15744 27112 15808
rect 27176 15744 27192 15808
rect 27256 15744 27262 15808
rect 26946 15743 27262 15744
rect 31946 15808 32262 15809
rect 31946 15744 31952 15808
rect 32016 15744 32032 15808
rect 32096 15744 32112 15808
rect 32176 15744 32192 15808
rect 32256 15744 32262 15808
rect 31946 15743 32262 15744
rect 36946 15808 37262 15809
rect 36946 15744 36952 15808
rect 37016 15744 37032 15808
rect 37096 15744 37112 15808
rect 37176 15744 37192 15808
rect 37256 15744 37262 15808
rect 36946 15743 37262 15744
rect 41946 15808 42262 15809
rect 41946 15744 41952 15808
rect 42016 15744 42032 15808
rect 42096 15744 42112 15808
rect 42176 15744 42192 15808
rect 42256 15744 42262 15808
rect 41946 15743 42262 15744
rect 46946 15808 47262 15809
rect 46946 15744 46952 15808
rect 47016 15744 47032 15808
rect 47096 15744 47112 15808
rect 47176 15744 47192 15808
rect 47256 15744 47262 15808
rect 46946 15743 47262 15744
rect 51946 15808 52262 15809
rect 51946 15744 51952 15808
rect 52016 15744 52032 15808
rect 52096 15744 52112 15808
rect 52176 15744 52192 15808
rect 52256 15744 52262 15808
rect 51946 15743 52262 15744
rect 56946 15808 57262 15809
rect 56946 15744 56952 15808
rect 57016 15744 57032 15808
rect 57096 15744 57112 15808
rect 57176 15744 57192 15808
rect 57256 15744 57262 15808
rect 56946 15743 57262 15744
rect 58525 15602 58591 15605
rect 59200 15602 60000 15632
rect 58525 15600 60000 15602
rect 58525 15544 58530 15600
rect 58586 15544 60000 15600
rect 58525 15542 60000 15544
rect 58525 15539 58591 15542
rect 59200 15512 60000 15542
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 17606 15199 17922 15200
rect 22606 15264 22922 15265
rect 22606 15200 22612 15264
rect 22676 15200 22692 15264
rect 22756 15200 22772 15264
rect 22836 15200 22852 15264
rect 22916 15200 22922 15264
rect 22606 15199 22922 15200
rect 27606 15264 27922 15265
rect 27606 15200 27612 15264
rect 27676 15200 27692 15264
rect 27756 15200 27772 15264
rect 27836 15200 27852 15264
rect 27916 15200 27922 15264
rect 27606 15199 27922 15200
rect 32606 15264 32922 15265
rect 32606 15200 32612 15264
rect 32676 15200 32692 15264
rect 32756 15200 32772 15264
rect 32836 15200 32852 15264
rect 32916 15200 32922 15264
rect 32606 15199 32922 15200
rect 37606 15264 37922 15265
rect 37606 15200 37612 15264
rect 37676 15200 37692 15264
rect 37756 15200 37772 15264
rect 37836 15200 37852 15264
rect 37916 15200 37922 15264
rect 37606 15199 37922 15200
rect 42606 15264 42922 15265
rect 42606 15200 42612 15264
rect 42676 15200 42692 15264
rect 42756 15200 42772 15264
rect 42836 15200 42852 15264
rect 42916 15200 42922 15264
rect 42606 15199 42922 15200
rect 47606 15264 47922 15265
rect 47606 15200 47612 15264
rect 47676 15200 47692 15264
rect 47756 15200 47772 15264
rect 47836 15200 47852 15264
rect 47916 15200 47922 15264
rect 47606 15199 47922 15200
rect 52606 15264 52922 15265
rect 52606 15200 52612 15264
rect 52676 15200 52692 15264
rect 52756 15200 52772 15264
rect 52836 15200 52852 15264
rect 52916 15200 52922 15264
rect 52606 15199 52922 15200
rect 57606 15264 57922 15265
rect 57606 15200 57612 15264
rect 57676 15200 57692 15264
rect 57756 15200 57772 15264
rect 57836 15200 57852 15264
rect 57916 15200 57922 15264
rect 57606 15199 57922 15200
rect 58525 14786 58591 14789
rect 59200 14786 60000 14816
rect 58525 14784 60000 14786
rect 58525 14728 58530 14784
rect 58586 14728 60000 14784
rect 58525 14726 60000 14728
rect 58525 14723 58591 14726
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 21946 14720 22262 14721
rect 21946 14656 21952 14720
rect 22016 14656 22032 14720
rect 22096 14656 22112 14720
rect 22176 14656 22192 14720
rect 22256 14656 22262 14720
rect 21946 14655 22262 14656
rect 26946 14720 27262 14721
rect 26946 14656 26952 14720
rect 27016 14656 27032 14720
rect 27096 14656 27112 14720
rect 27176 14656 27192 14720
rect 27256 14656 27262 14720
rect 26946 14655 27262 14656
rect 31946 14720 32262 14721
rect 31946 14656 31952 14720
rect 32016 14656 32032 14720
rect 32096 14656 32112 14720
rect 32176 14656 32192 14720
rect 32256 14656 32262 14720
rect 31946 14655 32262 14656
rect 36946 14720 37262 14721
rect 36946 14656 36952 14720
rect 37016 14656 37032 14720
rect 37096 14656 37112 14720
rect 37176 14656 37192 14720
rect 37256 14656 37262 14720
rect 36946 14655 37262 14656
rect 41946 14720 42262 14721
rect 41946 14656 41952 14720
rect 42016 14656 42032 14720
rect 42096 14656 42112 14720
rect 42176 14656 42192 14720
rect 42256 14656 42262 14720
rect 41946 14655 42262 14656
rect 46946 14720 47262 14721
rect 46946 14656 46952 14720
rect 47016 14656 47032 14720
rect 47096 14656 47112 14720
rect 47176 14656 47192 14720
rect 47256 14656 47262 14720
rect 46946 14655 47262 14656
rect 51946 14720 52262 14721
rect 51946 14656 51952 14720
rect 52016 14656 52032 14720
rect 52096 14656 52112 14720
rect 52176 14656 52192 14720
rect 52256 14656 52262 14720
rect 51946 14655 52262 14656
rect 56946 14720 57262 14721
rect 56946 14656 56952 14720
rect 57016 14656 57032 14720
rect 57096 14656 57112 14720
rect 57176 14656 57192 14720
rect 57256 14656 57262 14720
rect 59200 14696 60000 14726
rect 56946 14655 57262 14656
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 17606 14111 17922 14112
rect 22606 14176 22922 14177
rect 22606 14112 22612 14176
rect 22676 14112 22692 14176
rect 22756 14112 22772 14176
rect 22836 14112 22852 14176
rect 22916 14112 22922 14176
rect 22606 14111 22922 14112
rect 27606 14176 27922 14177
rect 27606 14112 27612 14176
rect 27676 14112 27692 14176
rect 27756 14112 27772 14176
rect 27836 14112 27852 14176
rect 27916 14112 27922 14176
rect 27606 14111 27922 14112
rect 32606 14176 32922 14177
rect 32606 14112 32612 14176
rect 32676 14112 32692 14176
rect 32756 14112 32772 14176
rect 32836 14112 32852 14176
rect 32916 14112 32922 14176
rect 32606 14111 32922 14112
rect 37606 14176 37922 14177
rect 37606 14112 37612 14176
rect 37676 14112 37692 14176
rect 37756 14112 37772 14176
rect 37836 14112 37852 14176
rect 37916 14112 37922 14176
rect 37606 14111 37922 14112
rect 42606 14176 42922 14177
rect 42606 14112 42612 14176
rect 42676 14112 42692 14176
rect 42756 14112 42772 14176
rect 42836 14112 42852 14176
rect 42916 14112 42922 14176
rect 42606 14111 42922 14112
rect 47606 14176 47922 14177
rect 47606 14112 47612 14176
rect 47676 14112 47692 14176
rect 47756 14112 47772 14176
rect 47836 14112 47852 14176
rect 47916 14112 47922 14176
rect 47606 14111 47922 14112
rect 52606 14176 52922 14177
rect 52606 14112 52612 14176
rect 52676 14112 52692 14176
rect 52756 14112 52772 14176
rect 52836 14112 52852 14176
rect 52916 14112 52922 14176
rect 52606 14111 52922 14112
rect 57606 14176 57922 14177
rect 57606 14112 57612 14176
rect 57676 14112 57692 14176
rect 57756 14112 57772 14176
rect 57836 14112 57852 14176
rect 57916 14112 57922 14176
rect 57606 14111 57922 14112
rect 58525 13970 58591 13973
rect 59200 13970 60000 14000
rect 58525 13968 60000 13970
rect 58525 13912 58530 13968
rect 58586 13912 60000 13968
rect 58525 13910 60000 13912
rect 58525 13907 58591 13910
rect 59200 13880 60000 13910
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 16946 13567 17262 13568
rect 21946 13632 22262 13633
rect 21946 13568 21952 13632
rect 22016 13568 22032 13632
rect 22096 13568 22112 13632
rect 22176 13568 22192 13632
rect 22256 13568 22262 13632
rect 21946 13567 22262 13568
rect 26946 13632 27262 13633
rect 26946 13568 26952 13632
rect 27016 13568 27032 13632
rect 27096 13568 27112 13632
rect 27176 13568 27192 13632
rect 27256 13568 27262 13632
rect 26946 13567 27262 13568
rect 31946 13632 32262 13633
rect 31946 13568 31952 13632
rect 32016 13568 32032 13632
rect 32096 13568 32112 13632
rect 32176 13568 32192 13632
rect 32256 13568 32262 13632
rect 31946 13567 32262 13568
rect 36946 13632 37262 13633
rect 36946 13568 36952 13632
rect 37016 13568 37032 13632
rect 37096 13568 37112 13632
rect 37176 13568 37192 13632
rect 37256 13568 37262 13632
rect 36946 13567 37262 13568
rect 41946 13632 42262 13633
rect 41946 13568 41952 13632
rect 42016 13568 42032 13632
rect 42096 13568 42112 13632
rect 42176 13568 42192 13632
rect 42256 13568 42262 13632
rect 41946 13567 42262 13568
rect 46946 13632 47262 13633
rect 46946 13568 46952 13632
rect 47016 13568 47032 13632
rect 47096 13568 47112 13632
rect 47176 13568 47192 13632
rect 47256 13568 47262 13632
rect 46946 13567 47262 13568
rect 51946 13632 52262 13633
rect 51946 13568 51952 13632
rect 52016 13568 52032 13632
rect 52096 13568 52112 13632
rect 52176 13568 52192 13632
rect 52256 13568 52262 13632
rect 51946 13567 52262 13568
rect 56946 13632 57262 13633
rect 56946 13568 56952 13632
rect 57016 13568 57032 13632
rect 57096 13568 57112 13632
rect 57176 13568 57192 13632
rect 57256 13568 57262 13632
rect 56946 13567 57262 13568
rect 58525 13154 58591 13157
rect 59200 13154 60000 13184
rect 58525 13152 60000 13154
rect 58525 13096 58530 13152
rect 58586 13096 60000 13152
rect 58525 13094 60000 13096
rect 58525 13091 58591 13094
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 17606 13023 17922 13024
rect 22606 13088 22922 13089
rect 22606 13024 22612 13088
rect 22676 13024 22692 13088
rect 22756 13024 22772 13088
rect 22836 13024 22852 13088
rect 22916 13024 22922 13088
rect 22606 13023 22922 13024
rect 27606 13088 27922 13089
rect 27606 13024 27612 13088
rect 27676 13024 27692 13088
rect 27756 13024 27772 13088
rect 27836 13024 27852 13088
rect 27916 13024 27922 13088
rect 27606 13023 27922 13024
rect 32606 13088 32922 13089
rect 32606 13024 32612 13088
rect 32676 13024 32692 13088
rect 32756 13024 32772 13088
rect 32836 13024 32852 13088
rect 32916 13024 32922 13088
rect 32606 13023 32922 13024
rect 37606 13088 37922 13089
rect 37606 13024 37612 13088
rect 37676 13024 37692 13088
rect 37756 13024 37772 13088
rect 37836 13024 37852 13088
rect 37916 13024 37922 13088
rect 37606 13023 37922 13024
rect 42606 13088 42922 13089
rect 42606 13024 42612 13088
rect 42676 13024 42692 13088
rect 42756 13024 42772 13088
rect 42836 13024 42852 13088
rect 42916 13024 42922 13088
rect 42606 13023 42922 13024
rect 47606 13088 47922 13089
rect 47606 13024 47612 13088
rect 47676 13024 47692 13088
rect 47756 13024 47772 13088
rect 47836 13024 47852 13088
rect 47916 13024 47922 13088
rect 47606 13023 47922 13024
rect 52606 13088 52922 13089
rect 52606 13024 52612 13088
rect 52676 13024 52692 13088
rect 52756 13024 52772 13088
rect 52836 13024 52852 13088
rect 52916 13024 52922 13088
rect 52606 13023 52922 13024
rect 57606 13088 57922 13089
rect 57606 13024 57612 13088
rect 57676 13024 57692 13088
rect 57756 13024 57772 13088
rect 57836 13024 57852 13088
rect 57916 13024 57922 13088
rect 59200 13064 60000 13094
rect 57606 13023 57922 13024
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 21946 12544 22262 12545
rect 21946 12480 21952 12544
rect 22016 12480 22032 12544
rect 22096 12480 22112 12544
rect 22176 12480 22192 12544
rect 22256 12480 22262 12544
rect 21946 12479 22262 12480
rect 26946 12544 27262 12545
rect 26946 12480 26952 12544
rect 27016 12480 27032 12544
rect 27096 12480 27112 12544
rect 27176 12480 27192 12544
rect 27256 12480 27262 12544
rect 26946 12479 27262 12480
rect 31946 12544 32262 12545
rect 31946 12480 31952 12544
rect 32016 12480 32032 12544
rect 32096 12480 32112 12544
rect 32176 12480 32192 12544
rect 32256 12480 32262 12544
rect 31946 12479 32262 12480
rect 36946 12544 37262 12545
rect 36946 12480 36952 12544
rect 37016 12480 37032 12544
rect 37096 12480 37112 12544
rect 37176 12480 37192 12544
rect 37256 12480 37262 12544
rect 36946 12479 37262 12480
rect 41946 12544 42262 12545
rect 41946 12480 41952 12544
rect 42016 12480 42032 12544
rect 42096 12480 42112 12544
rect 42176 12480 42192 12544
rect 42256 12480 42262 12544
rect 41946 12479 42262 12480
rect 46946 12544 47262 12545
rect 46946 12480 46952 12544
rect 47016 12480 47032 12544
rect 47096 12480 47112 12544
rect 47176 12480 47192 12544
rect 47256 12480 47262 12544
rect 46946 12479 47262 12480
rect 51946 12544 52262 12545
rect 51946 12480 51952 12544
rect 52016 12480 52032 12544
rect 52096 12480 52112 12544
rect 52176 12480 52192 12544
rect 52256 12480 52262 12544
rect 51946 12479 52262 12480
rect 56946 12544 57262 12545
rect 56946 12480 56952 12544
rect 57016 12480 57032 12544
rect 57096 12480 57112 12544
rect 57176 12480 57192 12544
rect 57256 12480 57262 12544
rect 56946 12479 57262 12480
rect 58525 12338 58591 12341
rect 59200 12338 60000 12368
rect 58525 12336 60000 12338
rect 58525 12280 58530 12336
rect 58586 12280 60000 12336
rect 58525 12278 60000 12280
rect 58525 12275 58591 12278
rect 59200 12248 60000 12278
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 17606 11935 17922 11936
rect 22606 12000 22922 12001
rect 22606 11936 22612 12000
rect 22676 11936 22692 12000
rect 22756 11936 22772 12000
rect 22836 11936 22852 12000
rect 22916 11936 22922 12000
rect 22606 11935 22922 11936
rect 27606 12000 27922 12001
rect 27606 11936 27612 12000
rect 27676 11936 27692 12000
rect 27756 11936 27772 12000
rect 27836 11936 27852 12000
rect 27916 11936 27922 12000
rect 27606 11935 27922 11936
rect 32606 12000 32922 12001
rect 32606 11936 32612 12000
rect 32676 11936 32692 12000
rect 32756 11936 32772 12000
rect 32836 11936 32852 12000
rect 32916 11936 32922 12000
rect 32606 11935 32922 11936
rect 37606 12000 37922 12001
rect 37606 11936 37612 12000
rect 37676 11936 37692 12000
rect 37756 11936 37772 12000
rect 37836 11936 37852 12000
rect 37916 11936 37922 12000
rect 37606 11935 37922 11936
rect 42606 12000 42922 12001
rect 42606 11936 42612 12000
rect 42676 11936 42692 12000
rect 42756 11936 42772 12000
rect 42836 11936 42852 12000
rect 42916 11936 42922 12000
rect 42606 11935 42922 11936
rect 47606 12000 47922 12001
rect 47606 11936 47612 12000
rect 47676 11936 47692 12000
rect 47756 11936 47772 12000
rect 47836 11936 47852 12000
rect 47916 11936 47922 12000
rect 47606 11935 47922 11936
rect 52606 12000 52922 12001
rect 52606 11936 52612 12000
rect 52676 11936 52692 12000
rect 52756 11936 52772 12000
rect 52836 11936 52852 12000
rect 52916 11936 52922 12000
rect 52606 11935 52922 11936
rect 57606 12000 57922 12001
rect 57606 11936 57612 12000
rect 57676 11936 57692 12000
rect 57756 11936 57772 12000
rect 57836 11936 57852 12000
rect 57916 11936 57922 12000
rect 57606 11935 57922 11936
rect 58525 11522 58591 11525
rect 59200 11522 60000 11552
rect 58525 11520 60000 11522
rect 58525 11464 58530 11520
rect 58586 11464 60000 11520
rect 58525 11462 60000 11464
rect 58525 11459 58591 11462
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 21946 11456 22262 11457
rect 21946 11392 21952 11456
rect 22016 11392 22032 11456
rect 22096 11392 22112 11456
rect 22176 11392 22192 11456
rect 22256 11392 22262 11456
rect 21946 11391 22262 11392
rect 26946 11456 27262 11457
rect 26946 11392 26952 11456
rect 27016 11392 27032 11456
rect 27096 11392 27112 11456
rect 27176 11392 27192 11456
rect 27256 11392 27262 11456
rect 26946 11391 27262 11392
rect 31946 11456 32262 11457
rect 31946 11392 31952 11456
rect 32016 11392 32032 11456
rect 32096 11392 32112 11456
rect 32176 11392 32192 11456
rect 32256 11392 32262 11456
rect 31946 11391 32262 11392
rect 36946 11456 37262 11457
rect 36946 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37262 11456
rect 36946 11391 37262 11392
rect 41946 11456 42262 11457
rect 41946 11392 41952 11456
rect 42016 11392 42032 11456
rect 42096 11392 42112 11456
rect 42176 11392 42192 11456
rect 42256 11392 42262 11456
rect 41946 11391 42262 11392
rect 46946 11456 47262 11457
rect 46946 11392 46952 11456
rect 47016 11392 47032 11456
rect 47096 11392 47112 11456
rect 47176 11392 47192 11456
rect 47256 11392 47262 11456
rect 46946 11391 47262 11392
rect 51946 11456 52262 11457
rect 51946 11392 51952 11456
rect 52016 11392 52032 11456
rect 52096 11392 52112 11456
rect 52176 11392 52192 11456
rect 52256 11392 52262 11456
rect 51946 11391 52262 11392
rect 56946 11456 57262 11457
rect 56946 11392 56952 11456
rect 57016 11392 57032 11456
rect 57096 11392 57112 11456
rect 57176 11392 57192 11456
rect 57256 11392 57262 11456
rect 59200 11432 60000 11462
rect 56946 11391 57262 11392
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 17606 10847 17922 10848
rect 22606 10912 22922 10913
rect 22606 10848 22612 10912
rect 22676 10848 22692 10912
rect 22756 10848 22772 10912
rect 22836 10848 22852 10912
rect 22916 10848 22922 10912
rect 22606 10847 22922 10848
rect 27606 10912 27922 10913
rect 27606 10848 27612 10912
rect 27676 10848 27692 10912
rect 27756 10848 27772 10912
rect 27836 10848 27852 10912
rect 27916 10848 27922 10912
rect 27606 10847 27922 10848
rect 32606 10912 32922 10913
rect 32606 10848 32612 10912
rect 32676 10848 32692 10912
rect 32756 10848 32772 10912
rect 32836 10848 32852 10912
rect 32916 10848 32922 10912
rect 32606 10847 32922 10848
rect 37606 10912 37922 10913
rect 37606 10848 37612 10912
rect 37676 10848 37692 10912
rect 37756 10848 37772 10912
rect 37836 10848 37852 10912
rect 37916 10848 37922 10912
rect 37606 10847 37922 10848
rect 42606 10912 42922 10913
rect 42606 10848 42612 10912
rect 42676 10848 42692 10912
rect 42756 10848 42772 10912
rect 42836 10848 42852 10912
rect 42916 10848 42922 10912
rect 42606 10847 42922 10848
rect 47606 10912 47922 10913
rect 47606 10848 47612 10912
rect 47676 10848 47692 10912
rect 47756 10848 47772 10912
rect 47836 10848 47852 10912
rect 47916 10848 47922 10912
rect 47606 10847 47922 10848
rect 52606 10912 52922 10913
rect 52606 10848 52612 10912
rect 52676 10848 52692 10912
rect 52756 10848 52772 10912
rect 52836 10848 52852 10912
rect 52916 10848 52922 10912
rect 52606 10847 52922 10848
rect 57606 10912 57922 10913
rect 57606 10848 57612 10912
rect 57676 10848 57692 10912
rect 57756 10848 57772 10912
rect 57836 10848 57852 10912
rect 57916 10848 57922 10912
rect 57606 10847 57922 10848
rect 58525 10706 58591 10709
rect 59200 10706 60000 10736
rect 58525 10704 60000 10706
rect 58525 10648 58530 10704
rect 58586 10648 60000 10704
rect 58525 10646 60000 10648
rect 58525 10643 58591 10646
rect 59200 10616 60000 10646
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 16946 10303 17262 10304
rect 21946 10368 22262 10369
rect 21946 10304 21952 10368
rect 22016 10304 22032 10368
rect 22096 10304 22112 10368
rect 22176 10304 22192 10368
rect 22256 10304 22262 10368
rect 21946 10303 22262 10304
rect 26946 10368 27262 10369
rect 26946 10304 26952 10368
rect 27016 10304 27032 10368
rect 27096 10304 27112 10368
rect 27176 10304 27192 10368
rect 27256 10304 27262 10368
rect 26946 10303 27262 10304
rect 31946 10368 32262 10369
rect 31946 10304 31952 10368
rect 32016 10304 32032 10368
rect 32096 10304 32112 10368
rect 32176 10304 32192 10368
rect 32256 10304 32262 10368
rect 31946 10303 32262 10304
rect 36946 10368 37262 10369
rect 36946 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37262 10368
rect 36946 10303 37262 10304
rect 41946 10368 42262 10369
rect 41946 10304 41952 10368
rect 42016 10304 42032 10368
rect 42096 10304 42112 10368
rect 42176 10304 42192 10368
rect 42256 10304 42262 10368
rect 41946 10303 42262 10304
rect 46946 10368 47262 10369
rect 46946 10304 46952 10368
rect 47016 10304 47032 10368
rect 47096 10304 47112 10368
rect 47176 10304 47192 10368
rect 47256 10304 47262 10368
rect 46946 10303 47262 10304
rect 51946 10368 52262 10369
rect 51946 10304 51952 10368
rect 52016 10304 52032 10368
rect 52096 10304 52112 10368
rect 52176 10304 52192 10368
rect 52256 10304 52262 10368
rect 51946 10303 52262 10304
rect 56946 10368 57262 10369
rect 56946 10304 56952 10368
rect 57016 10304 57032 10368
rect 57096 10304 57112 10368
rect 57176 10304 57192 10368
rect 57256 10304 57262 10368
rect 56946 10303 57262 10304
rect 0 10072 800 10192
rect 58525 9890 58591 9893
rect 59200 9890 60000 9920
rect 58525 9888 60000 9890
rect 58525 9832 58530 9888
rect 58586 9832 60000 9888
rect 58525 9830 60000 9832
rect 58525 9827 58591 9830
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 17606 9759 17922 9760
rect 22606 9824 22922 9825
rect 22606 9760 22612 9824
rect 22676 9760 22692 9824
rect 22756 9760 22772 9824
rect 22836 9760 22852 9824
rect 22916 9760 22922 9824
rect 22606 9759 22922 9760
rect 27606 9824 27922 9825
rect 27606 9760 27612 9824
rect 27676 9760 27692 9824
rect 27756 9760 27772 9824
rect 27836 9760 27852 9824
rect 27916 9760 27922 9824
rect 27606 9759 27922 9760
rect 32606 9824 32922 9825
rect 32606 9760 32612 9824
rect 32676 9760 32692 9824
rect 32756 9760 32772 9824
rect 32836 9760 32852 9824
rect 32916 9760 32922 9824
rect 32606 9759 32922 9760
rect 37606 9824 37922 9825
rect 37606 9760 37612 9824
rect 37676 9760 37692 9824
rect 37756 9760 37772 9824
rect 37836 9760 37852 9824
rect 37916 9760 37922 9824
rect 37606 9759 37922 9760
rect 42606 9824 42922 9825
rect 42606 9760 42612 9824
rect 42676 9760 42692 9824
rect 42756 9760 42772 9824
rect 42836 9760 42852 9824
rect 42916 9760 42922 9824
rect 42606 9759 42922 9760
rect 47606 9824 47922 9825
rect 47606 9760 47612 9824
rect 47676 9760 47692 9824
rect 47756 9760 47772 9824
rect 47836 9760 47852 9824
rect 47916 9760 47922 9824
rect 47606 9759 47922 9760
rect 52606 9824 52922 9825
rect 52606 9760 52612 9824
rect 52676 9760 52692 9824
rect 52756 9760 52772 9824
rect 52836 9760 52852 9824
rect 52916 9760 52922 9824
rect 52606 9759 52922 9760
rect 57606 9824 57922 9825
rect 57606 9760 57612 9824
rect 57676 9760 57692 9824
rect 57756 9760 57772 9824
rect 57836 9760 57852 9824
rect 57916 9760 57922 9824
rect 59200 9800 60000 9830
rect 57606 9759 57922 9760
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 21946 9280 22262 9281
rect 21946 9216 21952 9280
rect 22016 9216 22032 9280
rect 22096 9216 22112 9280
rect 22176 9216 22192 9280
rect 22256 9216 22262 9280
rect 21946 9215 22262 9216
rect 26946 9280 27262 9281
rect 26946 9216 26952 9280
rect 27016 9216 27032 9280
rect 27096 9216 27112 9280
rect 27176 9216 27192 9280
rect 27256 9216 27262 9280
rect 26946 9215 27262 9216
rect 31946 9280 32262 9281
rect 31946 9216 31952 9280
rect 32016 9216 32032 9280
rect 32096 9216 32112 9280
rect 32176 9216 32192 9280
rect 32256 9216 32262 9280
rect 31946 9215 32262 9216
rect 36946 9280 37262 9281
rect 36946 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37262 9280
rect 36946 9215 37262 9216
rect 41946 9280 42262 9281
rect 41946 9216 41952 9280
rect 42016 9216 42032 9280
rect 42096 9216 42112 9280
rect 42176 9216 42192 9280
rect 42256 9216 42262 9280
rect 41946 9215 42262 9216
rect 46946 9280 47262 9281
rect 46946 9216 46952 9280
rect 47016 9216 47032 9280
rect 47096 9216 47112 9280
rect 47176 9216 47192 9280
rect 47256 9216 47262 9280
rect 46946 9215 47262 9216
rect 51946 9280 52262 9281
rect 51946 9216 51952 9280
rect 52016 9216 52032 9280
rect 52096 9216 52112 9280
rect 52176 9216 52192 9280
rect 52256 9216 52262 9280
rect 51946 9215 52262 9216
rect 56946 9280 57262 9281
rect 56946 9216 56952 9280
rect 57016 9216 57032 9280
rect 57096 9216 57112 9280
rect 57176 9216 57192 9280
rect 57256 9216 57262 9280
rect 56946 9215 57262 9216
rect 58525 9074 58591 9077
rect 59200 9074 60000 9104
rect 58525 9072 60000 9074
rect 58525 9016 58530 9072
rect 58586 9016 60000 9072
rect 58525 9014 60000 9016
rect 58525 9011 58591 9014
rect 59200 8984 60000 9014
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 17606 8671 17922 8672
rect 22606 8736 22922 8737
rect 22606 8672 22612 8736
rect 22676 8672 22692 8736
rect 22756 8672 22772 8736
rect 22836 8672 22852 8736
rect 22916 8672 22922 8736
rect 22606 8671 22922 8672
rect 27606 8736 27922 8737
rect 27606 8672 27612 8736
rect 27676 8672 27692 8736
rect 27756 8672 27772 8736
rect 27836 8672 27852 8736
rect 27916 8672 27922 8736
rect 27606 8671 27922 8672
rect 32606 8736 32922 8737
rect 32606 8672 32612 8736
rect 32676 8672 32692 8736
rect 32756 8672 32772 8736
rect 32836 8672 32852 8736
rect 32916 8672 32922 8736
rect 32606 8671 32922 8672
rect 37606 8736 37922 8737
rect 37606 8672 37612 8736
rect 37676 8672 37692 8736
rect 37756 8672 37772 8736
rect 37836 8672 37852 8736
rect 37916 8672 37922 8736
rect 37606 8671 37922 8672
rect 42606 8736 42922 8737
rect 42606 8672 42612 8736
rect 42676 8672 42692 8736
rect 42756 8672 42772 8736
rect 42836 8672 42852 8736
rect 42916 8672 42922 8736
rect 42606 8671 42922 8672
rect 47606 8736 47922 8737
rect 47606 8672 47612 8736
rect 47676 8672 47692 8736
rect 47756 8672 47772 8736
rect 47836 8672 47852 8736
rect 47916 8672 47922 8736
rect 47606 8671 47922 8672
rect 52606 8736 52922 8737
rect 52606 8672 52612 8736
rect 52676 8672 52692 8736
rect 52756 8672 52772 8736
rect 52836 8672 52852 8736
rect 52916 8672 52922 8736
rect 52606 8671 52922 8672
rect 57606 8736 57922 8737
rect 57606 8672 57612 8736
rect 57676 8672 57692 8736
rect 57756 8672 57772 8736
rect 57836 8672 57852 8736
rect 57916 8672 57922 8736
rect 57606 8671 57922 8672
rect 58525 8258 58591 8261
rect 59200 8258 60000 8288
rect 58525 8256 60000 8258
rect 58525 8200 58530 8256
rect 58586 8200 60000 8256
rect 58525 8198 60000 8200
rect 58525 8195 58591 8198
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 21946 8192 22262 8193
rect 21946 8128 21952 8192
rect 22016 8128 22032 8192
rect 22096 8128 22112 8192
rect 22176 8128 22192 8192
rect 22256 8128 22262 8192
rect 21946 8127 22262 8128
rect 26946 8192 27262 8193
rect 26946 8128 26952 8192
rect 27016 8128 27032 8192
rect 27096 8128 27112 8192
rect 27176 8128 27192 8192
rect 27256 8128 27262 8192
rect 26946 8127 27262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 36946 8192 37262 8193
rect 36946 8128 36952 8192
rect 37016 8128 37032 8192
rect 37096 8128 37112 8192
rect 37176 8128 37192 8192
rect 37256 8128 37262 8192
rect 36946 8127 37262 8128
rect 41946 8192 42262 8193
rect 41946 8128 41952 8192
rect 42016 8128 42032 8192
rect 42096 8128 42112 8192
rect 42176 8128 42192 8192
rect 42256 8128 42262 8192
rect 41946 8127 42262 8128
rect 46946 8192 47262 8193
rect 46946 8128 46952 8192
rect 47016 8128 47032 8192
rect 47096 8128 47112 8192
rect 47176 8128 47192 8192
rect 47256 8128 47262 8192
rect 46946 8127 47262 8128
rect 51946 8192 52262 8193
rect 51946 8128 51952 8192
rect 52016 8128 52032 8192
rect 52096 8128 52112 8192
rect 52176 8128 52192 8192
rect 52256 8128 52262 8192
rect 51946 8127 52262 8128
rect 56946 8192 57262 8193
rect 56946 8128 56952 8192
rect 57016 8128 57032 8192
rect 57096 8128 57112 8192
rect 57176 8128 57192 8192
rect 57256 8128 57262 8192
rect 59200 8168 60000 8198
rect 56946 8127 57262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 17606 7583 17922 7584
rect 22606 7648 22922 7649
rect 22606 7584 22612 7648
rect 22676 7584 22692 7648
rect 22756 7584 22772 7648
rect 22836 7584 22852 7648
rect 22916 7584 22922 7648
rect 22606 7583 22922 7584
rect 27606 7648 27922 7649
rect 27606 7584 27612 7648
rect 27676 7584 27692 7648
rect 27756 7584 27772 7648
rect 27836 7584 27852 7648
rect 27916 7584 27922 7648
rect 27606 7583 27922 7584
rect 32606 7648 32922 7649
rect 32606 7584 32612 7648
rect 32676 7584 32692 7648
rect 32756 7584 32772 7648
rect 32836 7584 32852 7648
rect 32916 7584 32922 7648
rect 32606 7583 32922 7584
rect 37606 7648 37922 7649
rect 37606 7584 37612 7648
rect 37676 7584 37692 7648
rect 37756 7584 37772 7648
rect 37836 7584 37852 7648
rect 37916 7584 37922 7648
rect 37606 7583 37922 7584
rect 42606 7648 42922 7649
rect 42606 7584 42612 7648
rect 42676 7584 42692 7648
rect 42756 7584 42772 7648
rect 42836 7584 42852 7648
rect 42916 7584 42922 7648
rect 42606 7583 42922 7584
rect 47606 7648 47922 7649
rect 47606 7584 47612 7648
rect 47676 7584 47692 7648
rect 47756 7584 47772 7648
rect 47836 7584 47852 7648
rect 47916 7584 47922 7648
rect 47606 7583 47922 7584
rect 52606 7648 52922 7649
rect 52606 7584 52612 7648
rect 52676 7584 52692 7648
rect 52756 7584 52772 7648
rect 52836 7584 52852 7648
rect 52916 7584 52922 7648
rect 52606 7583 52922 7584
rect 57606 7648 57922 7649
rect 57606 7584 57612 7648
rect 57676 7584 57692 7648
rect 57756 7584 57772 7648
rect 57836 7584 57852 7648
rect 57916 7584 57922 7648
rect 57606 7583 57922 7584
rect 58525 7442 58591 7445
rect 59200 7442 60000 7472
rect 58525 7440 60000 7442
rect 58525 7384 58530 7440
rect 58586 7384 60000 7440
rect 58525 7382 60000 7384
rect 58525 7379 58591 7382
rect 59200 7352 60000 7382
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 21946 7104 22262 7105
rect 21946 7040 21952 7104
rect 22016 7040 22032 7104
rect 22096 7040 22112 7104
rect 22176 7040 22192 7104
rect 22256 7040 22262 7104
rect 21946 7039 22262 7040
rect 26946 7104 27262 7105
rect 26946 7040 26952 7104
rect 27016 7040 27032 7104
rect 27096 7040 27112 7104
rect 27176 7040 27192 7104
rect 27256 7040 27262 7104
rect 26946 7039 27262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 36946 7104 37262 7105
rect 36946 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37262 7104
rect 36946 7039 37262 7040
rect 41946 7104 42262 7105
rect 41946 7040 41952 7104
rect 42016 7040 42032 7104
rect 42096 7040 42112 7104
rect 42176 7040 42192 7104
rect 42256 7040 42262 7104
rect 41946 7039 42262 7040
rect 46946 7104 47262 7105
rect 46946 7040 46952 7104
rect 47016 7040 47032 7104
rect 47096 7040 47112 7104
rect 47176 7040 47192 7104
rect 47256 7040 47262 7104
rect 46946 7039 47262 7040
rect 51946 7104 52262 7105
rect 51946 7040 51952 7104
rect 52016 7040 52032 7104
rect 52096 7040 52112 7104
rect 52176 7040 52192 7104
rect 52256 7040 52262 7104
rect 51946 7039 52262 7040
rect 56946 7104 57262 7105
rect 56946 7040 56952 7104
rect 57016 7040 57032 7104
rect 57096 7040 57112 7104
rect 57176 7040 57192 7104
rect 57256 7040 57262 7104
rect 56946 7039 57262 7040
rect 58525 6626 58591 6629
rect 59200 6626 60000 6656
rect 58525 6624 60000 6626
rect 58525 6568 58530 6624
rect 58586 6568 60000 6624
rect 58525 6566 60000 6568
rect 58525 6563 58591 6566
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 17606 6495 17922 6496
rect 22606 6560 22922 6561
rect 22606 6496 22612 6560
rect 22676 6496 22692 6560
rect 22756 6496 22772 6560
rect 22836 6496 22852 6560
rect 22916 6496 22922 6560
rect 22606 6495 22922 6496
rect 27606 6560 27922 6561
rect 27606 6496 27612 6560
rect 27676 6496 27692 6560
rect 27756 6496 27772 6560
rect 27836 6496 27852 6560
rect 27916 6496 27922 6560
rect 27606 6495 27922 6496
rect 32606 6560 32922 6561
rect 32606 6496 32612 6560
rect 32676 6496 32692 6560
rect 32756 6496 32772 6560
rect 32836 6496 32852 6560
rect 32916 6496 32922 6560
rect 32606 6495 32922 6496
rect 37606 6560 37922 6561
rect 37606 6496 37612 6560
rect 37676 6496 37692 6560
rect 37756 6496 37772 6560
rect 37836 6496 37852 6560
rect 37916 6496 37922 6560
rect 37606 6495 37922 6496
rect 42606 6560 42922 6561
rect 42606 6496 42612 6560
rect 42676 6496 42692 6560
rect 42756 6496 42772 6560
rect 42836 6496 42852 6560
rect 42916 6496 42922 6560
rect 42606 6495 42922 6496
rect 47606 6560 47922 6561
rect 47606 6496 47612 6560
rect 47676 6496 47692 6560
rect 47756 6496 47772 6560
rect 47836 6496 47852 6560
rect 47916 6496 47922 6560
rect 47606 6495 47922 6496
rect 52606 6560 52922 6561
rect 52606 6496 52612 6560
rect 52676 6496 52692 6560
rect 52756 6496 52772 6560
rect 52836 6496 52852 6560
rect 52916 6496 52922 6560
rect 52606 6495 52922 6496
rect 57606 6560 57922 6561
rect 57606 6496 57612 6560
rect 57676 6496 57692 6560
rect 57756 6496 57772 6560
rect 57836 6496 57852 6560
rect 57916 6496 57922 6560
rect 59200 6536 60000 6566
rect 57606 6495 57922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 21946 6016 22262 6017
rect 21946 5952 21952 6016
rect 22016 5952 22032 6016
rect 22096 5952 22112 6016
rect 22176 5952 22192 6016
rect 22256 5952 22262 6016
rect 21946 5951 22262 5952
rect 26946 6016 27262 6017
rect 26946 5952 26952 6016
rect 27016 5952 27032 6016
rect 27096 5952 27112 6016
rect 27176 5952 27192 6016
rect 27256 5952 27262 6016
rect 26946 5951 27262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 36946 6016 37262 6017
rect 36946 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37262 6016
rect 36946 5951 37262 5952
rect 41946 6016 42262 6017
rect 41946 5952 41952 6016
rect 42016 5952 42032 6016
rect 42096 5952 42112 6016
rect 42176 5952 42192 6016
rect 42256 5952 42262 6016
rect 41946 5951 42262 5952
rect 46946 6016 47262 6017
rect 46946 5952 46952 6016
rect 47016 5952 47032 6016
rect 47096 5952 47112 6016
rect 47176 5952 47192 6016
rect 47256 5952 47262 6016
rect 46946 5951 47262 5952
rect 51946 6016 52262 6017
rect 51946 5952 51952 6016
rect 52016 5952 52032 6016
rect 52096 5952 52112 6016
rect 52176 5952 52192 6016
rect 52256 5952 52262 6016
rect 51946 5951 52262 5952
rect 56946 6016 57262 6017
rect 56946 5952 56952 6016
rect 57016 5952 57032 6016
rect 57096 5952 57112 6016
rect 57176 5952 57192 6016
rect 57256 5952 57262 6016
rect 56946 5951 57262 5952
rect 58525 5810 58591 5813
rect 59200 5810 60000 5840
rect 58525 5808 60000 5810
rect 58525 5752 58530 5808
rect 58586 5752 60000 5808
rect 58525 5750 60000 5752
rect 58525 5747 58591 5750
rect 59200 5720 60000 5750
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 17606 5407 17922 5408
rect 22606 5472 22922 5473
rect 22606 5408 22612 5472
rect 22676 5408 22692 5472
rect 22756 5408 22772 5472
rect 22836 5408 22852 5472
rect 22916 5408 22922 5472
rect 22606 5407 22922 5408
rect 27606 5472 27922 5473
rect 27606 5408 27612 5472
rect 27676 5408 27692 5472
rect 27756 5408 27772 5472
rect 27836 5408 27852 5472
rect 27916 5408 27922 5472
rect 27606 5407 27922 5408
rect 32606 5472 32922 5473
rect 32606 5408 32612 5472
rect 32676 5408 32692 5472
rect 32756 5408 32772 5472
rect 32836 5408 32852 5472
rect 32916 5408 32922 5472
rect 32606 5407 32922 5408
rect 37606 5472 37922 5473
rect 37606 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37922 5472
rect 37606 5407 37922 5408
rect 42606 5472 42922 5473
rect 42606 5408 42612 5472
rect 42676 5408 42692 5472
rect 42756 5408 42772 5472
rect 42836 5408 42852 5472
rect 42916 5408 42922 5472
rect 42606 5407 42922 5408
rect 47606 5472 47922 5473
rect 47606 5408 47612 5472
rect 47676 5408 47692 5472
rect 47756 5408 47772 5472
rect 47836 5408 47852 5472
rect 47916 5408 47922 5472
rect 47606 5407 47922 5408
rect 52606 5472 52922 5473
rect 52606 5408 52612 5472
rect 52676 5408 52692 5472
rect 52756 5408 52772 5472
rect 52836 5408 52852 5472
rect 52916 5408 52922 5472
rect 52606 5407 52922 5408
rect 57606 5472 57922 5473
rect 57606 5408 57612 5472
rect 57676 5408 57692 5472
rect 57756 5408 57772 5472
rect 57836 5408 57852 5472
rect 57916 5408 57922 5472
rect 57606 5407 57922 5408
rect 58525 4994 58591 4997
rect 59200 4994 60000 5024
rect 58525 4992 60000 4994
rect 58525 4936 58530 4992
rect 58586 4936 60000 4992
rect 58525 4934 60000 4936
rect 58525 4931 58591 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 21946 4928 22262 4929
rect 21946 4864 21952 4928
rect 22016 4864 22032 4928
rect 22096 4864 22112 4928
rect 22176 4864 22192 4928
rect 22256 4864 22262 4928
rect 21946 4863 22262 4864
rect 26946 4928 27262 4929
rect 26946 4864 26952 4928
rect 27016 4864 27032 4928
rect 27096 4864 27112 4928
rect 27176 4864 27192 4928
rect 27256 4864 27262 4928
rect 26946 4863 27262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 36946 4928 37262 4929
rect 36946 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37262 4928
rect 36946 4863 37262 4864
rect 41946 4928 42262 4929
rect 41946 4864 41952 4928
rect 42016 4864 42032 4928
rect 42096 4864 42112 4928
rect 42176 4864 42192 4928
rect 42256 4864 42262 4928
rect 41946 4863 42262 4864
rect 46946 4928 47262 4929
rect 46946 4864 46952 4928
rect 47016 4864 47032 4928
rect 47096 4864 47112 4928
rect 47176 4864 47192 4928
rect 47256 4864 47262 4928
rect 46946 4863 47262 4864
rect 51946 4928 52262 4929
rect 51946 4864 51952 4928
rect 52016 4864 52032 4928
rect 52096 4864 52112 4928
rect 52176 4864 52192 4928
rect 52256 4864 52262 4928
rect 51946 4863 52262 4864
rect 56946 4928 57262 4929
rect 56946 4864 56952 4928
rect 57016 4864 57032 4928
rect 57096 4864 57112 4928
rect 57176 4864 57192 4928
rect 57256 4864 57262 4928
rect 59200 4904 60000 4934
rect 56946 4863 57262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 17606 4319 17922 4320
rect 22606 4384 22922 4385
rect 22606 4320 22612 4384
rect 22676 4320 22692 4384
rect 22756 4320 22772 4384
rect 22836 4320 22852 4384
rect 22916 4320 22922 4384
rect 22606 4319 22922 4320
rect 27606 4384 27922 4385
rect 27606 4320 27612 4384
rect 27676 4320 27692 4384
rect 27756 4320 27772 4384
rect 27836 4320 27852 4384
rect 27916 4320 27922 4384
rect 27606 4319 27922 4320
rect 32606 4384 32922 4385
rect 32606 4320 32612 4384
rect 32676 4320 32692 4384
rect 32756 4320 32772 4384
rect 32836 4320 32852 4384
rect 32916 4320 32922 4384
rect 32606 4319 32922 4320
rect 37606 4384 37922 4385
rect 37606 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37922 4384
rect 37606 4319 37922 4320
rect 42606 4384 42922 4385
rect 42606 4320 42612 4384
rect 42676 4320 42692 4384
rect 42756 4320 42772 4384
rect 42836 4320 42852 4384
rect 42916 4320 42922 4384
rect 42606 4319 42922 4320
rect 47606 4384 47922 4385
rect 47606 4320 47612 4384
rect 47676 4320 47692 4384
rect 47756 4320 47772 4384
rect 47836 4320 47852 4384
rect 47916 4320 47922 4384
rect 47606 4319 47922 4320
rect 52606 4384 52922 4385
rect 52606 4320 52612 4384
rect 52676 4320 52692 4384
rect 52756 4320 52772 4384
rect 52836 4320 52852 4384
rect 52916 4320 52922 4384
rect 52606 4319 52922 4320
rect 57606 4384 57922 4385
rect 57606 4320 57612 4384
rect 57676 4320 57692 4384
rect 57756 4320 57772 4384
rect 57836 4320 57852 4384
rect 57916 4320 57922 4384
rect 57606 4319 57922 4320
rect 58525 4178 58591 4181
rect 59200 4178 60000 4208
rect 58525 4176 60000 4178
rect 58525 4120 58530 4176
rect 58586 4120 60000 4176
rect 58525 4118 60000 4120
rect 58525 4115 58591 4118
rect 59200 4088 60000 4118
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 16946 3775 17262 3776
rect 21946 3840 22262 3841
rect 21946 3776 21952 3840
rect 22016 3776 22032 3840
rect 22096 3776 22112 3840
rect 22176 3776 22192 3840
rect 22256 3776 22262 3840
rect 21946 3775 22262 3776
rect 26946 3840 27262 3841
rect 26946 3776 26952 3840
rect 27016 3776 27032 3840
rect 27096 3776 27112 3840
rect 27176 3776 27192 3840
rect 27256 3776 27262 3840
rect 26946 3775 27262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 36946 3840 37262 3841
rect 36946 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37262 3840
rect 36946 3775 37262 3776
rect 41946 3840 42262 3841
rect 41946 3776 41952 3840
rect 42016 3776 42032 3840
rect 42096 3776 42112 3840
rect 42176 3776 42192 3840
rect 42256 3776 42262 3840
rect 41946 3775 42262 3776
rect 46946 3840 47262 3841
rect 46946 3776 46952 3840
rect 47016 3776 47032 3840
rect 47096 3776 47112 3840
rect 47176 3776 47192 3840
rect 47256 3776 47262 3840
rect 46946 3775 47262 3776
rect 51946 3840 52262 3841
rect 51946 3776 51952 3840
rect 52016 3776 52032 3840
rect 52096 3776 52112 3840
rect 52176 3776 52192 3840
rect 52256 3776 52262 3840
rect 51946 3775 52262 3776
rect 56946 3840 57262 3841
rect 56946 3776 56952 3840
rect 57016 3776 57032 3840
rect 57096 3776 57112 3840
rect 57176 3776 57192 3840
rect 57256 3776 57262 3840
rect 56946 3775 57262 3776
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 17606 3231 17922 3232
rect 22606 3296 22922 3297
rect 22606 3232 22612 3296
rect 22676 3232 22692 3296
rect 22756 3232 22772 3296
rect 22836 3232 22852 3296
rect 22916 3232 22922 3296
rect 22606 3231 22922 3232
rect 27606 3296 27922 3297
rect 27606 3232 27612 3296
rect 27676 3232 27692 3296
rect 27756 3232 27772 3296
rect 27836 3232 27852 3296
rect 27916 3232 27922 3296
rect 27606 3231 27922 3232
rect 32606 3296 32922 3297
rect 32606 3232 32612 3296
rect 32676 3232 32692 3296
rect 32756 3232 32772 3296
rect 32836 3232 32852 3296
rect 32916 3232 32922 3296
rect 32606 3231 32922 3232
rect 37606 3296 37922 3297
rect 37606 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37922 3296
rect 37606 3231 37922 3232
rect 42606 3296 42922 3297
rect 42606 3232 42612 3296
rect 42676 3232 42692 3296
rect 42756 3232 42772 3296
rect 42836 3232 42852 3296
rect 42916 3232 42922 3296
rect 42606 3231 42922 3232
rect 47606 3296 47922 3297
rect 47606 3232 47612 3296
rect 47676 3232 47692 3296
rect 47756 3232 47772 3296
rect 47836 3232 47852 3296
rect 47916 3232 47922 3296
rect 47606 3231 47922 3232
rect 52606 3296 52922 3297
rect 52606 3232 52612 3296
rect 52676 3232 52692 3296
rect 52756 3232 52772 3296
rect 52836 3232 52852 3296
rect 52916 3232 52922 3296
rect 52606 3231 52922 3232
rect 57606 3296 57922 3297
rect 57606 3232 57612 3296
rect 57676 3232 57692 3296
rect 57756 3232 57772 3296
rect 57836 3232 57852 3296
rect 57916 3232 57922 3296
rect 57606 3231 57922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 16946 2687 17262 2688
rect 21946 2752 22262 2753
rect 21946 2688 21952 2752
rect 22016 2688 22032 2752
rect 22096 2688 22112 2752
rect 22176 2688 22192 2752
rect 22256 2688 22262 2752
rect 21946 2687 22262 2688
rect 26946 2752 27262 2753
rect 26946 2688 26952 2752
rect 27016 2688 27032 2752
rect 27096 2688 27112 2752
rect 27176 2688 27192 2752
rect 27256 2688 27262 2752
rect 26946 2687 27262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 36946 2752 37262 2753
rect 36946 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37262 2752
rect 36946 2687 37262 2688
rect 41946 2752 42262 2753
rect 41946 2688 41952 2752
rect 42016 2688 42032 2752
rect 42096 2688 42112 2752
rect 42176 2688 42192 2752
rect 42256 2688 42262 2752
rect 41946 2687 42262 2688
rect 46946 2752 47262 2753
rect 46946 2688 46952 2752
rect 47016 2688 47032 2752
rect 47096 2688 47112 2752
rect 47176 2688 47192 2752
rect 47256 2688 47262 2752
rect 46946 2687 47262 2688
rect 51946 2752 52262 2753
rect 51946 2688 51952 2752
rect 52016 2688 52032 2752
rect 52096 2688 52112 2752
rect 52176 2688 52192 2752
rect 52256 2688 52262 2752
rect 51946 2687 52262 2688
rect 56946 2752 57262 2753
rect 56946 2688 56952 2752
rect 57016 2688 57032 2752
rect 57096 2688 57112 2752
rect 57176 2688 57192 2752
rect 57256 2688 57262 2752
rect 56946 2687 57262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 17606 2143 17922 2144
rect 22606 2208 22922 2209
rect 22606 2144 22612 2208
rect 22676 2144 22692 2208
rect 22756 2144 22772 2208
rect 22836 2144 22852 2208
rect 22916 2144 22922 2208
rect 22606 2143 22922 2144
rect 27606 2208 27922 2209
rect 27606 2144 27612 2208
rect 27676 2144 27692 2208
rect 27756 2144 27772 2208
rect 27836 2144 27852 2208
rect 27916 2144 27922 2208
rect 27606 2143 27922 2144
rect 32606 2208 32922 2209
rect 32606 2144 32612 2208
rect 32676 2144 32692 2208
rect 32756 2144 32772 2208
rect 32836 2144 32852 2208
rect 32916 2144 32922 2208
rect 32606 2143 32922 2144
rect 37606 2208 37922 2209
rect 37606 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37922 2208
rect 37606 2143 37922 2144
rect 42606 2208 42922 2209
rect 42606 2144 42612 2208
rect 42676 2144 42692 2208
rect 42756 2144 42772 2208
rect 42836 2144 42852 2208
rect 42916 2144 42922 2208
rect 42606 2143 42922 2144
rect 47606 2208 47922 2209
rect 47606 2144 47612 2208
rect 47676 2144 47692 2208
rect 47756 2144 47772 2208
rect 47836 2144 47852 2208
rect 47916 2144 47922 2208
rect 47606 2143 47922 2144
rect 52606 2208 52922 2209
rect 52606 2144 52612 2208
rect 52676 2144 52692 2208
rect 52756 2144 52772 2208
rect 52836 2144 52852 2208
rect 52916 2144 52922 2208
rect 52606 2143 52922 2144
rect 57606 2208 57922 2209
rect 57606 2144 57612 2208
rect 57676 2144 57692 2208
rect 57756 2144 57772 2208
rect 57836 2144 57852 2208
rect 57916 2144 57922 2208
rect 57606 2143 57922 2144
<< via3 >>
rect 2612 57692 2676 57696
rect 2612 57636 2616 57692
rect 2616 57636 2672 57692
rect 2672 57636 2676 57692
rect 2612 57632 2676 57636
rect 2692 57692 2756 57696
rect 2692 57636 2696 57692
rect 2696 57636 2752 57692
rect 2752 57636 2756 57692
rect 2692 57632 2756 57636
rect 2772 57692 2836 57696
rect 2772 57636 2776 57692
rect 2776 57636 2832 57692
rect 2832 57636 2836 57692
rect 2772 57632 2836 57636
rect 2852 57692 2916 57696
rect 2852 57636 2856 57692
rect 2856 57636 2912 57692
rect 2912 57636 2916 57692
rect 2852 57632 2916 57636
rect 7612 57692 7676 57696
rect 7612 57636 7616 57692
rect 7616 57636 7672 57692
rect 7672 57636 7676 57692
rect 7612 57632 7676 57636
rect 7692 57692 7756 57696
rect 7692 57636 7696 57692
rect 7696 57636 7752 57692
rect 7752 57636 7756 57692
rect 7692 57632 7756 57636
rect 7772 57692 7836 57696
rect 7772 57636 7776 57692
rect 7776 57636 7832 57692
rect 7832 57636 7836 57692
rect 7772 57632 7836 57636
rect 7852 57692 7916 57696
rect 7852 57636 7856 57692
rect 7856 57636 7912 57692
rect 7912 57636 7916 57692
rect 7852 57632 7916 57636
rect 12612 57692 12676 57696
rect 12612 57636 12616 57692
rect 12616 57636 12672 57692
rect 12672 57636 12676 57692
rect 12612 57632 12676 57636
rect 12692 57692 12756 57696
rect 12692 57636 12696 57692
rect 12696 57636 12752 57692
rect 12752 57636 12756 57692
rect 12692 57632 12756 57636
rect 12772 57692 12836 57696
rect 12772 57636 12776 57692
rect 12776 57636 12832 57692
rect 12832 57636 12836 57692
rect 12772 57632 12836 57636
rect 12852 57692 12916 57696
rect 12852 57636 12856 57692
rect 12856 57636 12912 57692
rect 12912 57636 12916 57692
rect 12852 57632 12916 57636
rect 17612 57692 17676 57696
rect 17612 57636 17616 57692
rect 17616 57636 17672 57692
rect 17672 57636 17676 57692
rect 17612 57632 17676 57636
rect 17692 57692 17756 57696
rect 17692 57636 17696 57692
rect 17696 57636 17752 57692
rect 17752 57636 17756 57692
rect 17692 57632 17756 57636
rect 17772 57692 17836 57696
rect 17772 57636 17776 57692
rect 17776 57636 17832 57692
rect 17832 57636 17836 57692
rect 17772 57632 17836 57636
rect 17852 57692 17916 57696
rect 17852 57636 17856 57692
rect 17856 57636 17912 57692
rect 17912 57636 17916 57692
rect 17852 57632 17916 57636
rect 22612 57692 22676 57696
rect 22612 57636 22616 57692
rect 22616 57636 22672 57692
rect 22672 57636 22676 57692
rect 22612 57632 22676 57636
rect 22692 57692 22756 57696
rect 22692 57636 22696 57692
rect 22696 57636 22752 57692
rect 22752 57636 22756 57692
rect 22692 57632 22756 57636
rect 22772 57692 22836 57696
rect 22772 57636 22776 57692
rect 22776 57636 22832 57692
rect 22832 57636 22836 57692
rect 22772 57632 22836 57636
rect 22852 57692 22916 57696
rect 22852 57636 22856 57692
rect 22856 57636 22912 57692
rect 22912 57636 22916 57692
rect 22852 57632 22916 57636
rect 27612 57692 27676 57696
rect 27612 57636 27616 57692
rect 27616 57636 27672 57692
rect 27672 57636 27676 57692
rect 27612 57632 27676 57636
rect 27692 57692 27756 57696
rect 27692 57636 27696 57692
rect 27696 57636 27752 57692
rect 27752 57636 27756 57692
rect 27692 57632 27756 57636
rect 27772 57692 27836 57696
rect 27772 57636 27776 57692
rect 27776 57636 27832 57692
rect 27832 57636 27836 57692
rect 27772 57632 27836 57636
rect 27852 57692 27916 57696
rect 27852 57636 27856 57692
rect 27856 57636 27912 57692
rect 27912 57636 27916 57692
rect 27852 57632 27916 57636
rect 32612 57692 32676 57696
rect 32612 57636 32616 57692
rect 32616 57636 32672 57692
rect 32672 57636 32676 57692
rect 32612 57632 32676 57636
rect 32692 57692 32756 57696
rect 32692 57636 32696 57692
rect 32696 57636 32752 57692
rect 32752 57636 32756 57692
rect 32692 57632 32756 57636
rect 32772 57692 32836 57696
rect 32772 57636 32776 57692
rect 32776 57636 32832 57692
rect 32832 57636 32836 57692
rect 32772 57632 32836 57636
rect 32852 57692 32916 57696
rect 32852 57636 32856 57692
rect 32856 57636 32912 57692
rect 32912 57636 32916 57692
rect 32852 57632 32916 57636
rect 37612 57692 37676 57696
rect 37612 57636 37616 57692
rect 37616 57636 37672 57692
rect 37672 57636 37676 57692
rect 37612 57632 37676 57636
rect 37692 57692 37756 57696
rect 37692 57636 37696 57692
rect 37696 57636 37752 57692
rect 37752 57636 37756 57692
rect 37692 57632 37756 57636
rect 37772 57692 37836 57696
rect 37772 57636 37776 57692
rect 37776 57636 37832 57692
rect 37832 57636 37836 57692
rect 37772 57632 37836 57636
rect 37852 57692 37916 57696
rect 37852 57636 37856 57692
rect 37856 57636 37912 57692
rect 37912 57636 37916 57692
rect 37852 57632 37916 57636
rect 42612 57692 42676 57696
rect 42612 57636 42616 57692
rect 42616 57636 42672 57692
rect 42672 57636 42676 57692
rect 42612 57632 42676 57636
rect 42692 57692 42756 57696
rect 42692 57636 42696 57692
rect 42696 57636 42752 57692
rect 42752 57636 42756 57692
rect 42692 57632 42756 57636
rect 42772 57692 42836 57696
rect 42772 57636 42776 57692
rect 42776 57636 42832 57692
rect 42832 57636 42836 57692
rect 42772 57632 42836 57636
rect 42852 57692 42916 57696
rect 42852 57636 42856 57692
rect 42856 57636 42912 57692
rect 42912 57636 42916 57692
rect 42852 57632 42916 57636
rect 47612 57692 47676 57696
rect 47612 57636 47616 57692
rect 47616 57636 47672 57692
rect 47672 57636 47676 57692
rect 47612 57632 47676 57636
rect 47692 57692 47756 57696
rect 47692 57636 47696 57692
rect 47696 57636 47752 57692
rect 47752 57636 47756 57692
rect 47692 57632 47756 57636
rect 47772 57692 47836 57696
rect 47772 57636 47776 57692
rect 47776 57636 47832 57692
rect 47832 57636 47836 57692
rect 47772 57632 47836 57636
rect 47852 57692 47916 57696
rect 47852 57636 47856 57692
rect 47856 57636 47912 57692
rect 47912 57636 47916 57692
rect 47852 57632 47916 57636
rect 52612 57692 52676 57696
rect 52612 57636 52616 57692
rect 52616 57636 52672 57692
rect 52672 57636 52676 57692
rect 52612 57632 52676 57636
rect 52692 57692 52756 57696
rect 52692 57636 52696 57692
rect 52696 57636 52752 57692
rect 52752 57636 52756 57692
rect 52692 57632 52756 57636
rect 52772 57692 52836 57696
rect 52772 57636 52776 57692
rect 52776 57636 52832 57692
rect 52832 57636 52836 57692
rect 52772 57632 52836 57636
rect 52852 57692 52916 57696
rect 52852 57636 52856 57692
rect 52856 57636 52912 57692
rect 52912 57636 52916 57692
rect 52852 57632 52916 57636
rect 57612 57692 57676 57696
rect 57612 57636 57616 57692
rect 57616 57636 57672 57692
rect 57672 57636 57676 57692
rect 57612 57632 57676 57636
rect 57692 57692 57756 57696
rect 57692 57636 57696 57692
rect 57696 57636 57752 57692
rect 57752 57636 57756 57692
rect 57692 57632 57756 57636
rect 57772 57692 57836 57696
rect 57772 57636 57776 57692
rect 57776 57636 57832 57692
rect 57832 57636 57836 57692
rect 57772 57632 57836 57636
rect 57852 57692 57916 57696
rect 57852 57636 57856 57692
rect 57856 57636 57912 57692
rect 57912 57636 57916 57692
rect 57852 57632 57916 57636
rect 1952 57148 2016 57152
rect 1952 57092 1956 57148
rect 1956 57092 2012 57148
rect 2012 57092 2016 57148
rect 1952 57088 2016 57092
rect 2032 57148 2096 57152
rect 2032 57092 2036 57148
rect 2036 57092 2092 57148
rect 2092 57092 2096 57148
rect 2032 57088 2096 57092
rect 2112 57148 2176 57152
rect 2112 57092 2116 57148
rect 2116 57092 2172 57148
rect 2172 57092 2176 57148
rect 2112 57088 2176 57092
rect 2192 57148 2256 57152
rect 2192 57092 2196 57148
rect 2196 57092 2252 57148
rect 2252 57092 2256 57148
rect 2192 57088 2256 57092
rect 6952 57148 7016 57152
rect 6952 57092 6956 57148
rect 6956 57092 7012 57148
rect 7012 57092 7016 57148
rect 6952 57088 7016 57092
rect 7032 57148 7096 57152
rect 7032 57092 7036 57148
rect 7036 57092 7092 57148
rect 7092 57092 7096 57148
rect 7032 57088 7096 57092
rect 7112 57148 7176 57152
rect 7112 57092 7116 57148
rect 7116 57092 7172 57148
rect 7172 57092 7176 57148
rect 7112 57088 7176 57092
rect 7192 57148 7256 57152
rect 7192 57092 7196 57148
rect 7196 57092 7252 57148
rect 7252 57092 7256 57148
rect 7192 57088 7256 57092
rect 11952 57148 12016 57152
rect 11952 57092 11956 57148
rect 11956 57092 12012 57148
rect 12012 57092 12016 57148
rect 11952 57088 12016 57092
rect 12032 57148 12096 57152
rect 12032 57092 12036 57148
rect 12036 57092 12092 57148
rect 12092 57092 12096 57148
rect 12032 57088 12096 57092
rect 12112 57148 12176 57152
rect 12112 57092 12116 57148
rect 12116 57092 12172 57148
rect 12172 57092 12176 57148
rect 12112 57088 12176 57092
rect 12192 57148 12256 57152
rect 12192 57092 12196 57148
rect 12196 57092 12252 57148
rect 12252 57092 12256 57148
rect 12192 57088 12256 57092
rect 16952 57148 17016 57152
rect 16952 57092 16956 57148
rect 16956 57092 17012 57148
rect 17012 57092 17016 57148
rect 16952 57088 17016 57092
rect 17032 57148 17096 57152
rect 17032 57092 17036 57148
rect 17036 57092 17092 57148
rect 17092 57092 17096 57148
rect 17032 57088 17096 57092
rect 17112 57148 17176 57152
rect 17112 57092 17116 57148
rect 17116 57092 17172 57148
rect 17172 57092 17176 57148
rect 17112 57088 17176 57092
rect 17192 57148 17256 57152
rect 17192 57092 17196 57148
rect 17196 57092 17252 57148
rect 17252 57092 17256 57148
rect 17192 57088 17256 57092
rect 21952 57148 22016 57152
rect 21952 57092 21956 57148
rect 21956 57092 22012 57148
rect 22012 57092 22016 57148
rect 21952 57088 22016 57092
rect 22032 57148 22096 57152
rect 22032 57092 22036 57148
rect 22036 57092 22092 57148
rect 22092 57092 22096 57148
rect 22032 57088 22096 57092
rect 22112 57148 22176 57152
rect 22112 57092 22116 57148
rect 22116 57092 22172 57148
rect 22172 57092 22176 57148
rect 22112 57088 22176 57092
rect 22192 57148 22256 57152
rect 22192 57092 22196 57148
rect 22196 57092 22252 57148
rect 22252 57092 22256 57148
rect 22192 57088 22256 57092
rect 26952 57148 27016 57152
rect 26952 57092 26956 57148
rect 26956 57092 27012 57148
rect 27012 57092 27016 57148
rect 26952 57088 27016 57092
rect 27032 57148 27096 57152
rect 27032 57092 27036 57148
rect 27036 57092 27092 57148
rect 27092 57092 27096 57148
rect 27032 57088 27096 57092
rect 27112 57148 27176 57152
rect 27112 57092 27116 57148
rect 27116 57092 27172 57148
rect 27172 57092 27176 57148
rect 27112 57088 27176 57092
rect 27192 57148 27256 57152
rect 27192 57092 27196 57148
rect 27196 57092 27252 57148
rect 27252 57092 27256 57148
rect 27192 57088 27256 57092
rect 31952 57148 32016 57152
rect 31952 57092 31956 57148
rect 31956 57092 32012 57148
rect 32012 57092 32016 57148
rect 31952 57088 32016 57092
rect 32032 57148 32096 57152
rect 32032 57092 32036 57148
rect 32036 57092 32092 57148
rect 32092 57092 32096 57148
rect 32032 57088 32096 57092
rect 32112 57148 32176 57152
rect 32112 57092 32116 57148
rect 32116 57092 32172 57148
rect 32172 57092 32176 57148
rect 32112 57088 32176 57092
rect 32192 57148 32256 57152
rect 32192 57092 32196 57148
rect 32196 57092 32252 57148
rect 32252 57092 32256 57148
rect 32192 57088 32256 57092
rect 36952 57148 37016 57152
rect 36952 57092 36956 57148
rect 36956 57092 37012 57148
rect 37012 57092 37016 57148
rect 36952 57088 37016 57092
rect 37032 57148 37096 57152
rect 37032 57092 37036 57148
rect 37036 57092 37092 57148
rect 37092 57092 37096 57148
rect 37032 57088 37096 57092
rect 37112 57148 37176 57152
rect 37112 57092 37116 57148
rect 37116 57092 37172 57148
rect 37172 57092 37176 57148
rect 37112 57088 37176 57092
rect 37192 57148 37256 57152
rect 37192 57092 37196 57148
rect 37196 57092 37252 57148
rect 37252 57092 37256 57148
rect 37192 57088 37256 57092
rect 41952 57148 42016 57152
rect 41952 57092 41956 57148
rect 41956 57092 42012 57148
rect 42012 57092 42016 57148
rect 41952 57088 42016 57092
rect 42032 57148 42096 57152
rect 42032 57092 42036 57148
rect 42036 57092 42092 57148
rect 42092 57092 42096 57148
rect 42032 57088 42096 57092
rect 42112 57148 42176 57152
rect 42112 57092 42116 57148
rect 42116 57092 42172 57148
rect 42172 57092 42176 57148
rect 42112 57088 42176 57092
rect 42192 57148 42256 57152
rect 42192 57092 42196 57148
rect 42196 57092 42252 57148
rect 42252 57092 42256 57148
rect 42192 57088 42256 57092
rect 46952 57148 47016 57152
rect 46952 57092 46956 57148
rect 46956 57092 47012 57148
rect 47012 57092 47016 57148
rect 46952 57088 47016 57092
rect 47032 57148 47096 57152
rect 47032 57092 47036 57148
rect 47036 57092 47092 57148
rect 47092 57092 47096 57148
rect 47032 57088 47096 57092
rect 47112 57148 47176 57152
rect 47112 57092 47116 57148
rect 47116 57092 47172 57148
rect 47172 57092 47176 57148
rect 47112 57088 47176 57092
rect 47192 57148 47256 57152
rect 47192 57092 47196 57148
rect 47196 57092 47252 57148
rect 47252 57092 47256 57148
rect 47192 57088 47256 57092
rect 51952 57148 52016 57152
rect 51952 57092 51956 57148
rect 51956 57092 52012 57148
rect 52012 57092 52016 57148
rect 51952 57088 52016 57092
rect 52032 57148 52096 57152
rect 52032 57092 52036 57148
rect 52036 57092 52092 57148
rect 52092 57092 52096 57148
rect 52032 57088 52096 57092
rect 52112 57148 52176 57152
rect 52112 57092 52116 57148
rect 52116 57092 52172 57148
rect 52172 57092 52176 57148
rect 52112 57088 52176 57092
rect 52192 57148 52256 57152
rect 52192 57092 52196 57148
rect 52196 57092 52252 57148
rect 52252 57092 52256 57148
rect 52192 57088 52256 57092
rect 56952 57148 57016 57152
rect 56952 57092 56956 57148
rect 56956 57092 57012 57148
rect 57012 57092 57016 57148
rect 56952 57088 57016 57092
rect 57032 57148 57096 57152
rect 57032 57092 57036 57148
rect 57036 57092 57092 57148
rect 57092 57092 57096 57148
rect 57032 57088 57096 57092
rect 57112 57148 57176 57152
rect 57112 57092 57116 57148
rect 57116 57092 57172 57148
rect 57172 57092 57176 57148
rect 57112 57088 57176 57092
rect 57192 57148 57256 57152
rect 57192 57092 57196 57148
rect 57196 57092 57252 57148
rect 57252 57092 57256 57148
rect 57192 57088 57256 57092
rect 2612 56604 2676 56608
rect 2612 56548 2616 56604
rect 2616 56548 2672 56604
rect 2672 56548 2676 56604
rect 2612 56544 2676 56548
rect 2692 56604 2756 56608
rect 2692 56548 2696 56604
rect 2696 56548 2752 56604
rect 2752 56548 2756 56604
rect 2692 56544 2756 56548
rect 2772 56604 2836 56608
rect 2772 56548 2776 56604
rect 2776 56548 2832 56604
rect 2832 56548 2836 56604
rect 2772 56544 2836 56548
rect 2852 56604 2916 56608
rect 2852 56548 2856 56604
rect 2856 56548 2912 56604
rect 2912 56548 2916 56604
rect 2852 56544 2916 56548
rect 7612 56604 7676 56608
rect 7612 56548 7616 56604
rect 7616 56548 7672 56604
rect 7672 56548 7676 56604
rect 7612 56544 7676 56548
rect 7692 56604 7756 56608
rect 7692 56548 7696 56604
rect 7696 56548 7752 56604
rect 7752 56548 7756 56604
rect 7692 56544 7756 56548
rect 7772 56604 7836 56608
rect 7772 56548 7776 56604
rect 7776 56548 7832 56604
rect 7832 56548 7836 56604
rect 7772 56544 7836 56548
rect 7852 56604 7916 56608
rect 7852 56548 7856 56604
rect 7856 56548 7912 56604
rect 7912 56548 7916 56604
rect 7852 56544 7916 56548
rect 12612 56604 12676 56608
rect 12612 56548 12616 56604
rect 12616 56548 12672 56604
rect 12672 56548 12676 56604
rect 12612 56544 12676 56548
rect 12692 56604 12756 56608
rect 12692 56548 12696 56604
rect 12696 56548 12752 56604
rect 12752 56548 12756 56604
rect 12692 56544 12756 56548
rect 12772 56604 12836 56608
rect 12772 56548 12776 56604
rect 12776 56548 12832 56604
rect 12832 56548 12836 56604
rect 12772 56544 12836 56548
rect 12852 56604 12916 56608
rect 12852 56548 12856 56604
rect 12856 56548 12912 56604
rect 12912 56548 12916 56604
rect 12852 56544 12916 56548
rect 17612 56604 17676 56608
rect 17612 56548 17616 56604
rect 17616 56548 17672 56604
rect 17672 56548 17676 56604
rect 17612 56544 17676 56548
rect 17692 56604 17756 56608
rect 17692 56548 17696 56604
rect 17696 56548 17752 56604
rect 17752 56548 17756 56604
rect 17692 56544 17756 56548
rect 17772 56604 17836 56608
rect 17772 56548 17776 56604
rect 17776 56548 17832 56604
rect 17832 56548 17836 56604
rect 17772 56544 17836 56548
rect 17852 56604 17916 56608
rect 17852 56548 17856 56604
rect 17856 56548 17912 56604
rect 17912 56548 17916 56604
rect 17852 56544 17916 56548
rect 22612 56604 22676 56608
rect 22612 56548 22616 56604
rect 22616 56548 22672 56604
rect 22672 56548 22676 56604
rect 22612 56544 22676 56548
rect 22692 56604 22756 56608
rect 22692 56548 22696 56604
rect 22696 56548 22752 56604
rect 22752 56548 22756 56604
rect 22692 56544 22756 56548
rect 22772 56604 22836 56608
rect 22772 56548 22776 56604
rect 22776 56548 22832 56604
rect 22832 56548 22836 56604
rect 22772 56544 22836 56548
rect 22852 56604 22916 56608
rect 22852 56548 22856 56604
rect 22856 56548 22912 56604
rect 22912 56548 22916 56604
rect 22852 56544 22916 56548
rect 27612 56604 27676 56608
rect 27612 56548 27616 56604
rect 27616 56548 27672 56604
rect 27672 56548 27676 56604
rect 27612 56544 27676 56548
rect 27692 56604 27756 56608
rect 27692 56548 27696 56604
rect 27696 56548 27752 56604
rect 27752 56548 27756 56604
rect 27692 56544 27756 56548
rect 27772 56604 27836 56608
rect 27772 56548 27776 56604
rect 27776 56548 27832 56604
rect 27832 56548 27836 56604
rect 27772 56544 27836 56548
rect 27852 56604 27916 56608
rect 27852 56548 27856 56604
rect 27856 56548 27912 56604
rect 27912 56548 27916 56604
rect 27852 56544 27916 56548
rect 32612 56604 32676 56608
rect 32612 56548 32616 56604
rect 32616 56548 32672 56604
rect 32672 56548 32676 56604
rect 32612 56544 32676 56548
rect 32692 56604 32756 56608
rect 32692 56548 32696 56604
rect 32696 56548 32752 56604
rect 32752 56548 32756 56604
rect 32692 56544 32756 56548
rect 32772 56604 32836 56608
rect 32772 56548 32776 56604
rect 32776 56548 32832 56604
rect 32832 56548 32836 56604
rect 32772 56544 32836 56548
rect 32852 56604 32916 56608
rect 32852 56548 32856 56604
rect 32856 56548 32912 56604
rect 32912 56548 32916 56604
rect 32852 56544 32916 56548
rect 37612 56604 37676 56608
rect 37612 56548 37616 56604
rect 37616 56548 37672 56604
rect 37672 56548 37676 56604
rect 37612 56544 37676 56548
rect 37692 56604 37756 56608
rect 37692 56548 37696 56604
rect 37696 56548 37752 56604
rect 37752 56548 37756 56604
rect 37692 56544 37756 56548
rect 37772 56604 37836 56608
rect 37772 56548 37776 56604
rect 37776 56548 37832 56604
rect 37832 56548 37836 56604
rect 37772 56544 37836 56548
rect 37852 56604 37916 56608
rect 37852 56548 37856 56604
rect 37856 56548 37912 56604
rect 37912 56548 37916 56604
rect 37852 56544 37916 56548
rect 42612 56604 42676 56608
rect 42612 56548 42616 56604
rect 42616 56548 42672 56604
rect 42672 56548 42676 56604
rect 42612 56544 42676 56548
rect 42692 56604 42756 56608
rect 42692 56548 42696 56604
rect 42696 56548 42752 56604
rect 42752 56548 42756 56604
rect 42692 56544 42756 56548
rect 42772 56604 42836 56608
rect 42772 56548 42776 56604
rect 42776 56548 42832 56604
rect 42832 56548 42836 56604
rect 42772 56544 42836 56548
rect 42852 56604 42916 56608
rect 42852 56548 42856 56604
rect 42856 56548 42912 56604
rect 42912 56548 42916 56604
rect 42852 56544 42916 56548
rect 47612 56604 47676 56608
rect 47612 56548 47616 56604
rect 47616 56548 47672 56604
rect 47672 56548 47676 56604
rect 47612 56544 47676 56548
rect 47692 56604 47756 56608
rect 47692 56548 47696 56604
rect 47696 56548 47752 56604
rect 47752 56548 47756 56604
rect 47692 56544 47756 56548
rect 47772 56604 47836 56608
rect 47772 56548 47776 56604
rect 47776 56548 47832 56604
rect 47832 56548 47836 56604
rect 47772 56544 47836 56548
rect 47852 56604 47916 56608
rect 47852 56548 47856 56604
rect 47856 56548 47912 56604
rect 47912 56548 47916 56604
rect 47852 56544 47916 56548
rect 52612 56604 52676 56608
rect 52612 56548 52616 56604
rect 52616 56548 52672 56604
rect 52672 56548 52676 56604
rect 52612 56544 52676 56548
rect 52692 56604 52756 56608
rect 52692 56548 52696 56604
rect 52696 56548 52752 56604
rect 52752 56548 52756 56604
rect 52692 56544 52756 56548
rect 52772 56604 52836 56608
rect 52772 56548 52776 56604
rect 52776 56548 52832 56604
rect 52832 56548 52836 56604
rect 52772 56544 52836 56548
rect 52852 56604 52916 56608
rect 52852 56548 52856 56604
rect 52856 56548 52912 56604
rect 52912 56548 52916 56604
rect 52852 56544 52916 56548
rect 57612 56604 57676 56608
rect 57612 56548 57616 56604
rect 57616 56548 57672 56604
rect 57672 56548 57676 56604
rect 57612 56544 57676 56548
rect 57692 56604 57756 56608
rect 57692 56548 57696 56604
rect 57696 56548 57752 56604
rect 57752 56548 57756 56604
rect 57692 56544 57756 56548
rect 57772 56604 57836 56608
rect 57772 56548 57776 56604
rect 57776 56548 57832 56604
rect 57832 56548 57836 56604
rect 57772 56544 57836 56548
rect 57852 56604 57916 56608
rect 57852 56548 57856 56604
rect 57856 56548 57912 56604
rect 57912 56548 57916 56604
rect 57852 56544 57916 56548
rect 1952 56060 2016 56064
rect 1952 56004 1956 56060
rect 1956 56004 2012 56060
rect 2012 56004 2016 56060
rect 1952 56000 2016 56004
rect 2032 56060 2096 56064
rect 2032 56004 2036 56060
rect 2036 56004 2092 56060
rect 2092 56004 2096 56060
rect 2032 56000 2096 56004
rect 2112 56060 2176 56064
rect 2112 56004 2116 56060
rect 2116 56004 2172 56060
rect 2172 56004 2176 56060
rect 2112 56000 2176 56004
rect 2192 56060 2256 56064
rect 2192 56004 2196 56060
rect 2196 56004 2252 56060
rect 2252 56004 2256 56060
rect 2192 56000 2256 56004
rect 6952 56060 7016 56064
rect 6952 56004 6956 56060
rect 6956 56004 7012 56060
rect 7012 56004 7016 56060
rect 6952 56000 7016 56004
rect 7032 56060 7096 56064
rect 7032 56004 7036 56060
rect 7036 56004 7092 56060
rect 7092 56004 7096 56060
rect 7032 56000 7096 56004
rect 7112 56060 7176 56064
rect 7112 56004 7116 56060
rect 7116 56004 7172 56060
rect 7172 56004 7176 56060
rect 7112 56000 7176 56004
rect 7192 56060 7256 56064
rect 7192 56004 7196 56060
rect 7196 56004 7252 56060
rect 7252 56004 7256 56060
rect 7192 56000 7256 56004
rect 11952 56060 12016 56064
rect 11952 56004 11956 56060
rect 11956 56004 12012 56060
rect 12012 56004 12016 56060
rect 11952 56000 12016 56004
rect 12032 56060 12096 56064
rect 12032 56004 12036 56060
rect 12036 56004 12092 56060
rect 12092 56004 12096 56060
rect 12032 56000 12096 56004
rect 12112 56060 12176 56064
rect 12112 56004 12116 56060
rect 12116 56004 12172 56060
rect 12172 56004 12176 56060
rect 12112 56000 12176 56004
rect 12192 56060 12256 56064
rect 12192 56004 12196 56060
rect 12196 56004 12252 56060
rect 12252 56004 12256 56060
rect 12192 56000 12256 56004
rect 16952 56060 17016 56064
rect 16952 56004 16956 56060
rect 16956 56004 17012 56060
rect 17012 56004 17016 56060
rect 16952 56000 17016 56004
rect 17032 56060 17096 56064
rect 17032 56004 17036 56060
rect 17036 56004 17092 56060
rect 17092 56004 17096 56060
rect 17032 56000 17096 56004
rect 17112 56060 17176 56064
rect 17112 56004 17116 56060
rect 17116 56004 17172 56060
rect 17172 56004 17176 56060
rect 17112 56000 17176 56004
rect 17192 56060 17256 56064
rect 17192 56004 17196 56060
rect 17196 56004 17252 56060
rect 17252 56004 17256 56060
rect 17192 56000 17256 56004
rect 21952 56060 22016 56064
rect 21952 56004 21956 56060
rect 21956 56004 22012 56060
rect 22012 56004 22016 56060
rect 21952 56000 22016 56004
rect 22032 56060 22096 56064
rect 22032 56004 22036 56060
rect 22036 56004 22092 56060
rect 22092 56004 22096 56060
rect 22032 56000 22096 56004
rect 22112 56060 22176 56064
rect 22112 56004 22116 56060
rect 22116 56004 22172 56060
rect 22172 56004 22176 56060
rect 22112 56000 22176 56004
rect 22192 56060 22256 56064
rect 22192 56004 22196 56060
rect 22196 56004 22252 56060
rect 22252 56004 22256 56060
rect 22192 56000 22256 56004
rect 26952 56060 27016 56064
rect 26952 56004 26956 56060
rect 26956 56004 27012 56060
rect 27012 56004 27016 56060
rect 26952 56000 27016 56004
rect 27032 56060 27096 56064
rect 27032 56004 27036 56060
rect 27036 56004 27092 56060
rect 27092 56004 27096 56060
rect 27032 56000 27096 56004
rect 27112 56060 27176 56064
rect 27112 56004 27116 56060
rect 27116 56004 27172 56060
rect 27172 56004 27176 56060
rect 27112 56000 27176 56004
rect 27192 56060 27256 56064
rect 27192 56004 27196 56060
rect 27196 56004 27252 56060
rect 27252 56004 27256 56060
rect 27192 56000 27256 56004
rect 31952 56060 32016 56064
rect 31952 56004 31956 56060
rect 31956 56004 32012 56060
rect 32012 56004 32016 56060
rect 31952 56000 32016 56004
rect 32032 56060 32096 56064
rect 32032 56004 32036 56060
rect 32036 56004 32092 56060
rect 32092 56004 32096 56060
rect 32032 56000 32096 56004
rect 32112 56060 32176 56064
rect 32112 56004 32116 56060
rect 32116 56004 32172 56060
rect 32172 56004 32176 56060
rect 32112 56000 32176 56004
rect 32192 56060 32256 56064
rect 32192 56004 32196 56060
rect 32196 56004 32252 56060
rect 32252 56004 32256 56060
rect 32192 56000 32256 56004
rect 36952 56060 37016 56064
rect 36952 56004 36956 56060
rect 36956 56004 37012 56060
rect 37012 56004 37016 56060
rect 36952 56000 37016 56004
rect 37032 56060 37096 56064
rect 37032 56004 37036 56060
rect 37036 56004 37092 56060
rect 37092 56004 37096 56060
rect 37032 56000 37096 56004
rect 37112 56060 37176 56064
rect 37112 56004 37116 56060
rect 37116 56004 37172 56060
rect 37172 56004 37176 56060
rect 37112 56000 37176 56004
rect 37192 56060 37256 56064
rect 37192 56004 37196 56060
rect 37196 56004 37252 56060
rect 37252 56004 37256 56060
rect 37192 56000 37256 56004
rect 41952 56060 42016 56064
rect 41952 56004 41956 56060
rect 41956 56004 42012 56060
rect 42012 56004 42016 56060
rect 41952 56000 42016 56004
rect 42032 56060 42096 56064
rect 42032 56004 42036 56060
rect 42036 56004 42092 56060
rect 42092 56004 42096 56060
rect 42032 56000 42096 56004
rect 42112 56060 42176 56064
rect 42112 56004 42116 56060
rect 42116 56004 42172 56060
rect 42172 56004 42176 56060
rect 42112 56000 42176 56004
rect 42192 56060 42256 56064
rect 42192 56004 42196 56060
rect 42196 56004 42252 56060
rect 42252 56004 42256 56060
rect 42192 56000 42256 56004
rect 46952 56060 47016 56064
rect 46952 56004 46956 56060
rect 46956 56004 47012 56060
rect 47012 56004 47016 56060
rect 46952 56000 47016 56004
rect 47032 56060 47096 56064
rect 47032 56004 47036 56060
rect 47036 56004 47092 56060
rect 47092 56004 47096 56060
rect 47032 56000 47096 56004
rect 47112 56060 47176 56064
rect 47112 56004 47116 56060
rect 47116 56004 47172 56060
rect 47172 56004 47176 56060
rect 47112 56000 47176 56004
rect 47192 56060 47256 56064
rect 47192 56004 47196 56060
rect 47196 56004 47252 56060
rect 47252 56004 47256 56060
rect 47192 56000 47256 56004
rect 51952 56060 52016 56064
rect 51952 56004 51956 56060
rect 51956 56004 52012 56060
rect 52012 56004 52016 56060
rect 51952 56000 52016 56004
rect 52032 56060 52096 56064
rect 52032 56004 52036 56060
rect 52036 56004 52092 56060
rect 52092 56004 52096 56060
rect 52032 56000 52096 56004
rect 52112 56060 52176 56064
rect 52112 56004 52116 56060
rect 52116 56004 52172 56060
rect 52172 56004 52176 56060
rect 52112 56000 52176 56004
rect 52192 56060 52256 56064
rect 52192 56004 52196 56060
rect 52196 56004 52252 56060
rect 52252 56004 52256 56060
rect 52192 56000 52256 56004
rect 56952 56060 57016 56064
rect 56952 56004 56956 56060
rect 56956 56004 57012 56060
rect 57012 56004 57016 56060
rect 56952 56000 57016 56004
rect 57032 56060 57096 56064
rect 57032 56004 57036 56060
rect 57036 56004 57092 56060
rect 57092 56004 57096 56060
rect 57032 56000 57096 56004
rect 57112 56060 57176 56064
rect 57112 56004 57116 56060
rect 57116 56004 57172 56060
rect 57172 56004 57176 56060
rect 57112 56000 57176 56004
rect 57192 56060 57256 56064
rect 57192 56004 57196 56060
rect 57196 56004 57252 56060
rect 57252 56004 57256 56060
rect 57192 56000 57256 56004
rect 2612 55516 2676 55520
rect 2612 55460 2616 55516
rect 2616 55460 2672 55516
rect 2672 55460 2676 55516
rect 2612 55456 2676 55460
rect 2692 55516 2756 55520
rect 2692 55460 2696 55516
rect 2696 55460 2752 55516
rect 2752 55460 2756 55516
rect 2692 55456 2756 55460
rect 2772 55516 2836 55520
rect 2772 55460 2776 55516
rect 2776 55460 2832 55516
rect 2832 55460 2836 55516
rect 2772 55456 2836 55460
rect 2852 55516 2916 55520
rect 2852 55460 2856 55516
rect 2856 55460 2912 55516
rect 2912 55460 2916 55516
rect 2852 55456 2916 55460
rect 7612 55516 7676 55520
rect 7612 55460 7616 55516
rect 7616 55460 7672 55516
rect 7672 55460 7676 55516
rect 7612 55456 7676 55460
rect 7692 55516 7756 55520
rect 7692 55460 7696 55516
rect 7696 55460 7752 55516
rect 7752 55460 7756 55516
rect 7692 55456 7756 55460
rect 7772 55516 7836 55520
rect 7772 55460 7776 55516
rect 7776 55460 7832 55516
rect 7832 55460 7836 55516
rect 7772 55456 7836 55460
rect 7852 55516 7916 55520
rect 7852 55460 7856 55516
rect 7856 55460 7912 55516
rect 7912 55460 7916 55516
rect 7852 55456 7916 55460
rect 12612 55516 12676 55520
rect 12612 55460 12616 55516
rect 12616 55460 12672 55516
rect 12672 55460 12676 55516
rect 12612 55456 12676 55460
rect 12692 55516 12756 55520
rect 12692 55460 12696 55516
rect 12696 55460 12752 55516
rect 12752 55460 12756 55516
rect 12692 55456 12756 55460
rect 12772 55516 12836 55520
rect 12772 55460 12776 55516
rect 12776 55460 12832 55516
rect 12832 55460 12836 55516
rect 12772 55456 12836 55460
rect 12852 55516 12916 55520
rect 12852 55460 12856 55516
rect 12856 55460 12912 55516
rect 12912 55460 12916 55516
rect 12852 55456 12916 55460
rect 17612 55516 17676 55520
rect 17612 55460 17616 55516
rect 17616 55460 17672 55516
rect 17672 55460 17676 55516
rect 17612 55456 17676 55460
rect 17692 55516 17756 55520
rect 17692 55460 17696 55516
rect 17696 55460 17752 55516
rect 17752 55460 17756 55516
rect 17692 55456 17756 55460
rect 17772 55516 17836 55520
rect 17772 55460 17776 55516
rect 17776 55460 17832 55516
rect 17832 55460 17836 55516
rect 17772 55456 17836 55460
rect 17852 55516 17916 55520
rect 17852 55460 17856 55516
rect 17856 55460 17912 55516
rect 17912 55460 17916 55516
rect 17852 55456 17916 55460
rect 22612 55516 22676 55520
rect 22612 55460 22616 55516
rect 22616 55460 22672 55516
rect 22672 55460 22676 55516
rect 22612 55456 22676 55460
rect 22692 55516 22756 55520
rect 22692 55460 22696 55516
rect 22696 55460 22752 55516
rect 22752 55460 22756 55516
rect 22692 55456 22756 55460
rect 22772 55516 22836 55520
rect 22772 55460 22776 55516
rect 22776 55460 22832 55516
rect 22832 55460 22836 55516
rect 22772 55456 22836 55460
rect 22852 55516 22916 55520
rect 22852 55460 22856 55516
rect 22856 55460 22912 55516
rect 22912 55460 22916 55516
rect 22852 55456 22916 55460
rect 27612 55516 27676 55520
rect 27612 55460 27616 55516
rect 27616 55460 27672 55516
rect 27672 55460 27676 55516
rect 27612 55456 27676 55460
rect 27692 55516 27756 55520
rect 27692 55460 27696 55516
rect 27696 55460 27752 55516
rect 27752 55460 27756 55516
rect 27692 55456 27756 55460
rect 27772 55516 27836 55520
rect 27772 55460 27776 55516
rect 27776 55460 27832 55516
rect 27832 55460 27836 55516
rect 27772 55456 27836 55460
rect 27852 55516 27916 55520
rect 27852 55460 27856 55516
rect 27856 55460 27912 55516
rect 27912 55460 27916 55516
rect 27852 55456 27916 55460
rect 32612 55516 32676 55520
rect 32612 55460 32616 55516
rect 32616 55460 32672 55516
rect 32672 55460 32676 55516
rect 32612 55456 32676 55460
rect 32692 55516 32756 55520
rect 32692 55460 32696 55516
rect 32696 55460 32752 55516
rect 32752 55460 32756 55516
rect 32692 55456 32756 55460
rect 32772 55516 32836 55520
rect 32772 55460 32776 55516
rect 32776 55460 32832 55516
rect 32832 55460 32836 55516
rect 32772 55456 32836 55460
rect 32852 55516 32916 55520
rect 32852 55460 32856 55516
rect 32856 55460 32912 55516
rect 32912 55460 32916 55516
rect 32852 55456 32916 55460
rect 37612 55516 37676 55520
rect 37612 55460 37616 55516
rect 37616 55460 37672 55516
rect 37672 55460 37676 55516
rect 37612 55456 37676 55460
rect 37692 55516 37756 55520
rect 37692 55460 37696 55516
rect 37696 55460 37752 55516
rect 37752 55460 37756 55516
rect 37692 55456 37756 55460
rect 37772 55516 37836 55520
rect 37772 55460 37776 55516
rect 37776 55460 37832 55516
rect 37832 55460 37836 55516
rect 37772 55456 37836 55460
rect 37852 55516 37916 55520
rect 37852 55460 37856 55516
rect 37856 55460 37912 55516
rect 37912 55460 37916 55516
rect 37852 55456 37916 55460
rect 42612 55516 42676 55520
rect 42612 55460 42616 55516
rect 42616 55460 42672 55516
rect 42672 55460 42676 55516
rect 42612 55456 42676 55460
rect 42692 55516 42756 55520
rect 42692 55460 42696 55516
rect 42696 55460 42752 55516
rect 42752 55460 42756 55516
rect 42692 55456 42756 55460
rect 42772 55516 42836 55520
rect 42772 55460 42776 55516
rect 42776 55460 42832 55516
rect 42832 55460 42836 55516
rect 42772 55456 42836 55460
rect 42852 55516 42916 55520
rect 42852 55460 42856 55516
rect 42856 55460 42912 55516
rect 42912 55460 42916 55516
rect 42852 55456 42916 55460
rect 47612 55516 47676 55520
rect 47612 55460 47616 55516
rect 47616 55460 47672 55516
rect 47672 55460 47676 55516
rect 47612 55456 47676 55460
rect 47692 55516 47756 55520
rect 47692 55460 47696 55516
rect 47696 55460 47752 55516
rect 47752 55460 47756 55516
rect 47692 55456 47756 55460
rect 47772 55516 47836 55520
rect 47772 55460 47776 55516
rect 47776 55460 47832 55516
rect 47832 55460 47836 55516
rect 47772 55456 47836 55460
rect 47852 55516 47916 55520
rect 47852 55460 47856 55516
rect 47856 55460 47912 55516
rect 47912 55460 47916 55516
rect 47852 55456 47916 55460
rect 52612 55516 52676 55520
rect 52612 55460 52616 55516
rect 52616 55460 52672 55516
rect 52672 55460 52676 55516
rect 52612 55456 52676 55460
rect 52692 55516 52756 55520
rect 52692 55460 52696 55516
rect 52696 55460 52752 55516
rect 52752 55460 52756 55516
rect 52692 55456 52756 55460
rect 52772 55516 52836 55520
rect 52772 55460 52776 55516
rect 52776 55460 52832 55516
rect 52832 55460 52836 55516
rect 52772 55456 52836 55460
rect 52852 55516 52916 55520
rect 52852 55460 52856 55516
rect 52856 55460 52912 55516
rect 52912 55460 52916 55516
rect 52852 55456 52916 55460
rect 57612 55516 57676 55520
rect 57612 55460 57616 55516
rect 57616 55460 57672 55516
rect 57672 55460 57676 55516
rect 57612 55456 57676 55460
rect 57692 55516 57756 55520
rect 57692 55460 57696 55516
rect 57696 55460 57752 55516
rect 57752 55460 57756 55516
rect 57692 55456 57756 55460
rect 57772 55516 57836 55520
rect 57772 55460 57776 55516
rect 57776 55460 57832 55516
rect 57832 55460 57836 55516
rect 57772 55456 57836 55460
rect 57852 55516 57916 55520
rect 57852 55460 57856 55516
rect 57856 55460 57912 55516
rect 57912 55460 57916 55516
rect 57852 55456 57916 55460
rect 1952 54972 2016 54976
rect 1952 54916 1956 54972
rect 1956 54916 2012 54972
rect 2012 54916 2016 54972
rect 1952 54912 2016 54916
rect 2032 54972 2096 54976
rect 2032 54916 2036 54972
rect 2036 54916 2092 54972
rect 2092 54916 2096 54972
rect 2032 54912 2096 54916
rect 2112 54972 2176 54976
rect 2112 54916 2116 54972
rect 2116 54916 2172 54972
rect 2172 54916 2176 54972
rect 2112 54912 2176 54916
rect 2192 54972 2256 54976
rect 2192 54916 2196 54972
rect 2196 54916 2252 54972
rect 2252 54916 2256 54972
rect 2192 54912 2256 54916
rect 6952 54972 7016 54976
rect 6952 54916 6956 54972
rect 6956 54916 7012 54972
rect 7012 54916 7016 54972
rect 6952 54912 7016 54916
rect 7032 54972 7096 54976
rect 7032 54916 7036 54972
rect 7036 54916 7092 54972
rect 7092 54916 7096 54972
rect 7032 54912 7096 54916
rect 7112 54972 7176 54976
rect 7112 54916 7116 54972
rect 7116 54916 7172 54972
rect 7172 54916 7176 54972
rect 7112 54912 7176 54916
rect 7192 54972 7256 54976
rect 7192 54916 7196 54972
rect 7196 54916 7252 54972
rect 7252 54916 7256 54972
rect 7192 54912 7256 54916
rect 11952 54972 12016 54976
rect 11952 54916 11956 54972
rect 11956 54916 12012 54972
rect 12012 54916 12016 54972
rect 11952 54912 12016 54916
rect 12032 54972 12096 54976
rect 12032 54916 12036 54972
rect 12036 54916 12092 54972
rect 12092 54916 12096 54972
rect 12032 54912 12096 54916
rect 12112 54972 12176 54976
rect 12112 54916 12116 54972
rect 12116 54916 12172 54972
rect 12172 54916 12176 54972
rect 12112 54912 12176 54916
rect 12192 54972 12256 54976
rect 12192 54916 12196 54972
rect 12196 54916 12252 54972
rect 12252 54916 12256 54972
rect 12192 54912 12256 54916
rect 16952 54972 17016 54976
rect 16952 54916 16956 54972
rect 16956 54916 17012 54972
rect 17012 54916 17016 54972
rect 16952 54912 17016 54916
rect 17032 54972 17096 54976
rect 17032 54916 17036 54972
rect 17036 54916 17092 54972
rect 17092 54916 17096 54972
rect 17032 54912 17096 54916
rect 17112 54972 17176 54976
rect 17112 54916 17116 54972
rect 17116 54916 17172 54972
rect 17172 54916 17176 54972
rect 17112 54912 17176 54916
rect 17192 54972 17256 54976
rect 17192 54916 17196 54972
rect 17196 54916 17252 54972
rect 17252 54916 17256 54972
rect 17192 54912 17256 54916
rect 21952 54972 22016 54976
rect 21952 54916 21956 54972
rect 21956 54916 22012 54972
rect 22012 54916 22016 54972
rect 21952 54912 22016 54916
rect 22032 54972 22096 54976
rect 22032 54916 22036 54972
rect 22036 54916 22092 54972
rect 22092 54916 22096 54972
rect 22032 54912 22096 54916
rect 22112 54972 22176 54976
rect 22112 54916 22116 54972
rect 22116 54916 22172 54972
rect 22172 54916 22176 54972
rect 22112 54912 22176 54916
rect 22192 54972 22256 54976
rect 22192 54916 22196 54972
rect 22196 54916 22252 54972
rect 22252 54916 22256 54972
rect 22192 54912 22256 54916
rect 26952 54972 27016 54976
rect 26952 54916 26956 54972
rect 26956 54916 27012 54972
rect 27012 54916 27016 54972
rect 26952 54912 27016 54916
rect 27032 54972 27096 54976
rect 27032 54916 27036 54972
rect 27036 54916 27092 54972
rect 27092 54916 27096 54972
rect 27032 54912 27096 54916
rect 27112 54972 27176 54976
rect 27112 54916 27116 54972
rect 27116 54916 27172 54972
rect 27172 54916 27176 54972
rect 27112 54912 27176 54916
rect 27192 54972 27256 54976
rect 27192 54916 27196 54972
rect 27196 54916 27252 54972
rect 27252 54916 27256 54972
rect 27192 54912 27256 54916
rect 31952 54972 32016 54976
rect 31952 54916 31956 54972
rect 31956 54916 32012 54972
rect 32012 54916 32016 54972
rect 31952 54912 32016 54916
rect 32032 54972 32096 54976
rect 32032 54916 32036 54972
rect 32036 54916 32092 54972
rect 32092 54916 32096 54972
rect 32032 54912 32096 54916
rect 32112 54972 32176 54976
rect 32112 54916 32116 54972
rect 32116 54916 32172 54972
rect 32172 54916 32176 54972
rect 32112 54912 32176 54916
rect 32192 54972 32256 54976
rect 32192 54916 32196 54972
rect 32196 54916 32252 54972
rect 32252 54916 32256 54972
rect 32192 54912 32256 54916
rect 36952 54972 37016 54976
rect 36952 54916 36956 54972
rect 36956 54916 37012 54972
rect 37012 54916 37016 54972
rect 36952 54912 37016 54916
rect 37032 54972 37096 54976
rect 37032 54916 37036 54972
rect 37036 54916 37092 54972
rect 37092 54916 37096 54972
rect 37032 54912 37096 54916
rect 37112 54972 37176 54976
rect 37112 54916 37116 54972
rect 37116 54916 37172 54972
rect 37172 54916 37176 54972
rect 37112 54912 37176 54916
rect 37192 54972 37256 54976
rect 37192 54916 37196 54972
rect 37196 54916 37252 54972
rect 37252 54916 37256 54972
rect 37192 54912 37256 54916
rect 41952 54972 42016 54976
rect 41952 54916 41956 54972
rect 41956 54916 42012 54972
rect 42012 54916 42016 54972
rect 41952 54912 42016 54916
rect 42032 54972 42096 54976
rect 42032 54916 42036 54972
rect 42036 54916 42092 54972
rect 42092 54916 42096 54972
rect 42032 54912 42096 54916
rect 42112 54972 42176 54976
rect 42112 54916 42116 54972
rect 42116 54916 42172 54972
rect 42172 54916 42176 54972
rect 42112 54912 42176 54916
rect 42192 54972 42256 54976
rect 42192 54916 42196 54972
rect 42196 54916 42252 54972
rect 42252 54916 42256 54972
rect 42192 54912 42256 54916
rect 46952 54972 47016 54976
rect 46952 54916 46956 54972
rect 46956 54916 47012 54972
rect 47012 54916 47016 54972
rect 46952 54912 47016 54916
rect 47032 54972 47096 54976
rect 47032 54916 47036 54972
rect 47036 54916 47092 54972
rect 47092 54916 47096 54972
rect 47032 54912 47096 54916
rect 47112 54972 47176 54976
rect 47112 54916 47116 54972
rect 47116 54916 47172 54972
rect 47172 54916 47176 54972
rect 47112 54912 47176 54916
rect 47192 54972 47256 54976
rect 47192 54916 47196 54972
rect 47196 54916 47252 54972
rect 47252 54916 47256 54972
rect 47192 54912 47256 54916
rect 51952 54972 52016 54976
rect 51952 54916 51956 54972
rect 51956 54916 52012 54972
rect 52012 54916 52016 54972
rect 51952 54912 52016 54916
rect 52032 54972 52096 54976
rect 52032 54916 52036 54972
rect 52036 54916 52092 54972
rect 52092 54916 52096 54972
rect 52032 54912 52096 54916
rect 52112 54972 52176 54976
rect 52112 54916 52116 54972
rect 52116 54916 52172 54972
rect 52172 54916 52176 54972
rect 52112 54912 52176 54916
rect 52192 54972 52256 54976
rect 52192 54916 52196 54972
rect 52196 54916 52252 54972
rect 52252 54916 52256 54972
rect 52192 54912 52256 54916
rect 56952 54972 57016 54976
rect 56952 54916 56956 54972
rect 56956 54916 57012 54972
rect 57012 54916 57016 54972
rect 56952 54912 57016 54916
rect 57032 54972 57096 54976
rect 57032 54916 57036 54972
rect 57036 54916 57092 54972
rect 57092 54916 57096 54972
rect 57032 54912 57096 54916
rect 57112 54972 57176 54976
rect 57112 54916 57116 54972
rect 57116 54916 57172 54972
rect 57172 54916 57176 54972
rect 57112 54912 57176 54916
rect 57192 54972 57256 54976
rect 57192 54916 57196 54972
rect 57196 54916 57252 54972
rect 57252 54916 57256 54972
rect 57192 54912 57256 54916
rect 2612 54428 2676 54432
rect 2612 54372 2616 54428
rect 2616 54372 2672 54428
rect 2672 54372 2676 54428
rect 2612 54368 2676 54372
rect 2692 54428 2756 54432
rect 2692 54372 2696 54428
rect 2696 54372 2752 54428
rect 2752 54372 2756 54428
rect 2692 54368 2756 54372
rect 2772 54428 2836 54432
rect 2772 54372 2776 54428
rect 2776 54372 2832 54428
rect 2832 54372 2836 54428
rect 2772 54368 2836 54372
rect 2852 54428 2916 54432
rect 2852 54372 2856 54428
rect 2856 54372 2912 54428
rect 2912 54372 2916 54428
rect 2852 54368 2916 54372
rect 7612 54428 7676 54432
rect 7612 54372 7616 54428
rect 7616 54372 7672 54428
rect 7672 54372 7676 54428
rect 7612 54368 7676 54372
rect 7692 54428 7756 54432
rect 7692 54372 7696 54428
rect 7696 54372 7752 54428
rect 7752 54372 7756 54428
rect 7692 54368 7756 54372
rect 7772 54428 7836 54432
rect 7772 54372 7776 54428
rect 7776 54372 7832 54428
rect 7832 54372 7836 54428
rect 7772 54368 7836 54372
rect 7852 54428 7916 54432
rect 7852 54372 7856 54428
rect 7856 54372 7912 54428
rect 7912 54372 7916 54428
rect 7852 54368 7916 54372
rect 12612 54428 12676 54432
rect 12612 54372 12616 54428
rect 12616 54372 12672 54428
rect 12672 54372 12676 54428
rect 12612 54368 12676 54372
rect 12692 54428 12756 54432
rect 12692 54372 12696 54428
rect 12696 54372 12752 54428
rect 12752 54372 12756 54428
rect 12692 54368 12756 54372
rect 12772 54428 12836 54432
rect 12772 54372 12776 54428
rect 12776 54372 12832 54428
rect 12832 54372 12836 54428
rect 12772 54368 12836 54372
rect 12852 54428 12916 54432
rect 12852 54372 12856 54428
rect 12856 54372 12912 54428
rect 12912 54372 12916 54428
rect 12852 54368 12916 54372
rect 17612 54428 17676 54432
rect 17612 54372 17616 54428
rect 17616 54372 17672 54428
rect 17672 54372 17676 54428
rect 17612 54368 17676 54372
rect 17692 54428 17756 54432
rect 17692 54372 17696 54428
rect 17696 54372 17752 54428
rect 17752 54372 17756 54428
rect 17692 54368 17756 54372
rect 17772 54428 17836 54432
rect 17772 54372 17776 54428
rect 17776 54372 17832 54428
rect 17832 54372 17836 54428
rect 17772 54368 17836 54372
rect 17852 54428 17916 54432
rect 17852 54372 17856 54428
rect 17856 54372 17912 54428
rect 17912 54372 17916 54428
rect 17852 54368 17916 54372
rect 22612 54428 22676 54432
rect 22612 54372 22616 54428
rect 22616 54372 22672 54428
rect 22672 54372 22676 54428
rect 22612 54368 22676 54372
rect 22692 54428 22756 54432
rect 22692 54372 22696 54428
rect 22696 54372 22752 54428
rect 22752 54372 22756 54428
rect 22692 54368 22756 54372
rect 22772 54428 22836 54432
rect 22772 54372 22776 54428
rect 22776 54372 22832 54428
rect 22832 54372 22836 54428
rect 22772 54368 22836 54372
rect 22852 54428 22916 54432
rect 22852 54372 22856 54428
rect 22856 54372 22912 54428
rect 22912 54372 22916 54428
rect 22852 54368 22916 54372
rect 27612 54428 27676 54432
rect 27612 54372 27616 54428
rect 27616 54372 27672 54428
rect 27672 54372 27676 54428
rect 27612 54368 27676 54372
rect 27692 54428 27756 54432
rect 27692 54372 27696 54428
rect 27696 54372 27752 54428
rect 27752 54372 27756 54428
rect 27692 54368 27756 54372
rect 27772 54428 27836 54432
rect 27772 54372 27776 54428
rect 27776 54372 27832 54428
rect 27832 54372 27836 54428
rect 27772 54368 27836 54372
rect 27852 54428 27916 54432
rect 27852 54372 27856 54428
rect 27856 54372 27912 54428
rect 27912 54372 27916 54428
rect 27852 54368 27916 54372
rect 32612 54428 32676 54432
rect 32612 54372 32616 54428
rect 32616 54372 32672 54428
rect 32672 54372 32676 54428
rect 32612 54368 32676 54372
rect 32692 54428 32756 54432
rect 32692 54372 32696 54428
rect 32696 54372 32752 54428
rect 32752 54372 32756 54428
rect 32692 54368 32756 54372
rect 32772 54428 32836 54432
rect 32772 54372 32776 54428
rect 32776 54372 32832 54428
rect 32832 54372 32836 54428
rect 32772 54368 32836 54372
rect 32852 54428 32916 54432
rect 32852 54372 32856 54428
rect 32856 54372 32912 54428
rect 32912 54372 32916 54428
rect 32852 54368 32916 54372
rect 37612 54428 37676 54432
rect 37612 54372 37616 54428
rect 37616 54372 37672 54428
rect 37672 54372 37676 54428
rect 37612 54368 37676 54372
rect 37692 54428 37756 54432
rect 37692 54372 37696 54428
rect 37696 54372 37752 54428
rect 37752 54372 37756 54428
rect 37692 54368 37756 54372
rect 37772 54428 37836 54432
rect 37772 54372 37776 54428
rect 37776 54372 37832 54428
rect 37832 54372 37836 54428
rect 37772 54368 37836 54372
rect 37852 54428 37916 54432
rect 37852 54372 37856 54428
rect 37856 54372 37912 54428
rect 37912 54372 37916 54428
rect 37852 54368 37916 54372
rect 42612 54428 42676 54432
rect 42612 54372 42616 54428
rect 42616 54372 42672 54428
rect 42672 54372 42676 54428
rect 42612 54368 42676 54372
rect 42692 54428 42756 54432
rect 42692 54372 42696 54428
rect 42696 54372 42752 54428
rect 42752 54372 42756 54428
rect 42692 54368 42756 54372
rect 42772 54428 42836 54432
rect 42772 54372 42776 54428
rect 42776 54372 42832 54428
rect 42832 54372 42836 54428
rect 42772 54368 42836 54372
rect 42852 54428 42916 54432
rect 42852 54372 42856 54428
rect 42856 54372 42912 54428
rect 42912 54372 42916 54428
rect 42852 54368 42916 54372
rect 47612 54428 47676 54432
rect 47612 54372 47616 54428
rect 47616 54372 47672 54428
rect 47672 54372 47676 54428
rect 47612 54368 47676 54372
rect 47692 54428 47756 54432
rect 47692 54372 47696 54428
rect 47696 54372 47752 54428
rect 47752 54372 47756 54428
rect 47692 54368 47756 54372
rect 47772 54428 47836 54432
rect 47772 54372 47776 54428
rect 47776 54372 47832 54428
rect 47832 54372 47836 54428
rect 47772 54368 47836 54372
rect 47852 54428 47916 54432
rect 47852 54372 47856 54428
rect 47856 54372 47912 54428
rect 47912 54372 47916 54428
rect 47852 54368 47916 54372
rect 52612 54428 52676 54432
rect 52612 54372 52616 54428
rect 52616 54372 52672 54428
rect 52672 54372 52676 54428
rect 52612 54368 52676 54372
rect 52692 54428 52756 54432
rect 52692 54372 52696 54428
rect 52696 54372 52752 54428
rect 52752 54372 52756 54428
rect 52692 54368 52756 54372
rect 52772 54428 52836 54432
rect 52772 54372 52776 54428
rect 52776 54372 52832 54428
rect 52832 54372 52836 54428
rect 52772 54368 52836 54372
rect 52852 54428 52916 54432
rect 52852 54372 52856 54428
rect 52856 54372 52912 54428
rect 52912 54372 52916 54428
rect 52852 54368 52916 54372
rect 57612 54428 57676 54432
rect 57612 54372 57616 54428
rect 57616 54372 57672 54428
rect 57672 54372 57676 54428
rect 57612 54368 57676 54372
rect 57692 54428 57756 54432
rect 57692 54372 57696 54428
rect 57696 54372 57752 54428
rect 57752 54372 57756 54428
rect 57692 54368 57756 54372
rect 57772 54428 57836 54432
rect 57772 54372 57776 54428
rect 57776 54372 57832 54428
rect 57832 54372 57836 54428
rect 57772 54368 57836 54372
rect 57852 54428 57916 54432
rect 57852 54372 57856 54428
rect 57856 54372 57912 54428
rect 57912 54372 57916 54428
rect 57852 54368 57916 54372
rect 1952 53884 2016 53888
rect 1952 53828 1956 53884
rect 1956 53828 2012 53884
rect 2012 53828 2016 53884
rect 1952 53824 2016 53828
rect 2032 53884 2096 53888
rect 2032 53828 2036 53884
rect 2036 53828 2092 53884
rect 2092 53828 2096 53884
rect 2032 53824 2096 53828
rect 2112 53884 2176 53888
rect 2112 53828 2116 53884
rect 2116 53828 2172 53884
rect 2172 53828 2176 53884
rect 2112 53824 2176 53828
rect 2192 53884 2256 53888
rect 2192 53828 2196 53884
rect 2196 53828 2252 53884
rect 2252 53828 2256 53884
rect 2192 53824 2256 53828
rect 6952 53884 7016 53888
rect 6952 53828 6956 53884
rect 6956 53828 7012 53884
rect 7012 53828 7016 53884
rect 6952 53824 7016 53828
rect 7032 53884 7096 53888
rect 7032 53828 7036 53884
rect 7036 53828 7092 53884
rect 7092 53828 7096 53884
rect 7032 53824 7096 53828
rect 7112 53884 7176 53888
rect 7112 53828 7116 53884
rect 7116 53828 7172 53884
rect 7172 53828 7176 53884
rect 7112 53824 7176 53828
rect 7192 53884 7256 53888
rect 7192 53828 7196 53884
rect 7196 53828 7252 53884
rect 7252 53828 7256 53884
rect 7192 53824 7256 53828
rect 11952 53884 12016 53888
rect 11952 53828 11956 53884
rect 11956 53828 12012 53884
rect 12012 53828 12016 53884
rect 11952 53824 12016 53828
rect 12032 53884 12096 53888
rect 12032 53828 12036 53884
rect 12036 53828 12092 53884
rect 12092 53828 12096 53884
rect 12032 53824 12096 53828
rect 12112 53884 12176 53888
rect 12112 53828 12116 53884
rect 12116 53828 12172 53884
rect 12172 53828 12176 53884
rect 12112 53824 12176 53828
rect 12192 53884 12256 53888
rect 12192 53828 12196 53884
rect 12196 53828 12252 53884
rect 12252 53828 12256 53884
rect 12192 53824 12256 53828
rect 16952 53884 17016 53888
rect 16952 53828 16956 53884
rect 16956 53828 17012 53884
rect 17012 53828 17016 53884
rect 16952 53824 17016 53828
rect 17032 53884 17096 53888
rect 17032 53828 17036 53884
rect 17036 53828 17092 53884
rect 17092 53828 17096 53884
rect 17032 53824 17096 53828
rect 17112 53884 17176 53888
rect 17112 53828 17116 53884
rect 17116 53828 17172 53884
rect 17172 53828 17176 53884
rect 17112 53824 17176 53828
rect 17192 53884 17256 53888
rect 17192 53828 17196 53884
rect 17196 53828 17252 53884
rect 17252 53828 17256 53884
rect 17192 53824 17256 53828
rect 21952 53884 22016 53888
rect 21952 53828 21956 53884
rect 21956 53828 22012 53884
rect 22012 53828 22016 53884
rect 21952 53824 22016 53828
rect 22032 53884 22096 53888
rect 22032 53828 22036 53884
rect 22036 53828 22092 53884
rect 22092 53828 22096 53884
rect 22032 53824 22096 53828
rect 22112 53884 22176 53888
rect 22112 53828 22116 53884
rect 22116 53828 22172 53884
rect 22172 53828 22176 53884
rect 22112 53824 22176 53828
rect 22192 53884 22256 53888
rect 22192 53828 22196 53884
rect 22196 53828 22252 53884
rect 22252 53828 22256 53884
rect 22192 53824 22256 53828
rect 26952 53884 27016 53888
rect 26952 53828 26956 53884
rect 26956 53828 27012 53884
rect 27012 53828 27016 53884
rect 26952 53824 27016 53828
rect 27032 53884 27096 53888
rect 27032 53828 27036 53884
rect 27036 53828 27092 53884
rect 27092 53828 27096 53884
rect 27032 53824 27096 53828
rect 27112 53884 27176 53888
rect 27112 53828 27116 53884
rect 27116 53828 27172 53884
rect 27172 53828 27176 53884
rect 27112 53824 27176 53828
rect 27192 53884 27256 53888
rect 27192 53828 27196 53884
rect 27196 53828 27252 53884
rect 27252 53828 27256 53884
rect 27192 53824 27256 53828
rect 31952 53884 32016 53888
rect 31952 53828 31956 53884
rect 31956 53828 32012 53884
rect 32012 53828 32016 53884
rect 31952 53824 32016 53828
rect 32032 53884 32096 53888
rect 32032 53828 32036 53884
rect 32036 53828 32092 53884
rect 32092 53828 32096 53884
rect 32032 53824 32096 53828
rect 32112 53884 32176 53888
rect 32112 53828 32116 53884
rect 32116 53828 32172 53884
rect 32172 53828 32176 53884
rect 32112 53824 32176 53828
rect 32192 53884 32256 53888
rect 32192 53828 32196 53884
rect 32196 53828 32252 53884
rect 32252 53828 32256 53884
rect 32192 53824 32256 53828
rect 36952 53884 37016 53888
rect 36952 53828 36956 53884
rect 36956 53828 37012 53884
rect 37012 53828 37016 53884
rect 36952 53824 37016 53828
rect 37032 53884 37096 53888
rect 37032 53828 37036 53884
rect 37036 53828 37092 53884
rect 37092 53828 37096 53884
rect 37032 53824 37096 53828
rect 37112 53884 37176 53888
rect 37112 53828 37116 53884
rect 37116 53828 37172 53884
rect 37172 53828 37176 53884
rect 37112 53824 37176 53828
rect 37192 53884 37256 53888
rect 37192 53828 37196 53884
rect 37196 53828 37252 53884
rect 37252 53828 37256 53884
rect 37192 53824 37256 53828
rect 41952 53884 42016 53888
rect 41952 53828 41956 53884
rect 41956 53828 42012 53884
rect 42012 53828 42016 53884
rect 41952 53824 42016 53828
rect 42032 53884 42096 53888
rect 42032 53828 42036 53884
rect 42036 53828 42092 53884
rect 42092 53828 42096 53884
rect 42032 53824 42096 53828
rect 42112 53884 42176 53888
rect 42112 53828 42116 53884
rect 42116 53828 42172 53884
rect 42172 53828 42176 53884
rect 42112 53824 42176 53828
rect 42192 53884 42256 53888
rect 42192 53828 42196 53884
rect 42196 53828 42252 53884
rect 42252 53828 42256 53884
rect 42192 53824 42256 53828
rect 46952 53884 47016 53888
rect 46952 53828 46956 53884
rect 46956 53828 47012 53884
rect 47012 53828 47016 53884
rect 46952 53824 47016 53828
rect 47032 53884 47096 53888
rect 47032 53828 47036 53884
rect 47036 53828 47092 53884
rect 47092 53828 47096 53884
rect 47032 53824 47096 53828
rect 47112 53884 47176 53888
rect 47112 53828 47116 53884
rect 47116 53828 47172 53884
rect 47172 53828 47176 53884
rect 47112 53824 47176 53828
rect 47192 53884 47256 53888
rect 47192 53828 47196 53884
rect 47196 53828 47252 53884
rect 47252 53828 47256 53884
rect 47192 53824 47256 53828
rect 51952 53884 52016 53888
rect 51952 53828 51956 53884
rect 51956 53828 52012 53884
rect 52012 53828 52016 53884
rect 51952 53824 52016 53828
rect 52032 53884 52096 53888
rect 52032 53828 52036 53884
rect 52036 53828 52092 53884
rect 52092 53828 52096 53884
rect 52032 53824 52096 53828
rect 52112 53884 52176 53888
rect 52112 53828 52116 53884
rect 52116 53828 52172 53884
rect 52172 53828 52176 53884
rect 52112 53824 52176 53828
rect 52192 53884 52256 53888
rect 52192 53828 52196 53884
rect 52196 53828 52252 53884
rect 52252 53828 52256 53884
rect 52192 53824 52256 53828
rect 56952 53884 57016 53888
rect 56952 53828 56956 53884
rect 56956 53828 57012 53884
rect 57012 53828 57016 53884
rect 56952 53824 57016 53828
rect 57032 53884 57096 53888
rect 57032 53828 57036 53884
rect 57036 53828 57092 53884
rect 57092 53828 57096 53884
rect 57032 53824 57096 53828
rect 57112 53884 57176 53888
rect 57112 53828 57116 53884
rect 57116 53828 57172 53884
rect 57172 53828 57176 53884
rect 57112 53824 57176 53828
rect 57192 53884 57256 53888
rect 57192 53828 57196 53884
rect 57196 53828 57252 53884
rect 57252 53828 57256 53884
rect 57192 53824 57256 53828
rect 2612 53340 2676 53344
rect 2612 53284 2616 53340
rect 2616 53284 2672 53340
rect 2672 53284 2676 53340
rect 2612 53280 2676 53284
rect 2692 53340 2756 53344
rect 2692 53284 2696 53340
rect 2696 53284 2752 53340
rect 2752 53284 2756 53340
rect 2692 53280 2756 53284
rect 2772 53340 2836 53344
rect 2772 53284 2776 53340
rect 2776 53284 2832 53340
rect 2832 53284 2836 53340
rect 2772 53280 2836 53284
rect 2852 53340 2916 53344
rect 2852 53284 2856 53340
rect 2856 53284 2912 53340
rect 2912 53284 2916 53340
rect 2852 53280 2916 53284
rect 7612 53340 7676 53344
rect 7612 53284 7616 53340
rect 7616 53284 7672 53340
rect 7672 53284 7676 53340
rect 7612 53280 7676 53284
rect 7692 53340 7756 53344
rect 7692 53284 7696 53340
rect 7696 53284 7752 53340
rect 7752 53284 7756 53340
rect 7692 53280 7756 53284
rect 7772 53340 7836 53344
rect 7772 53284 7776 53340
rect 7776 53284 7832 53340
rect 7832 53284 7836 53340
rect 7772 53280 7836 53284
rect 7852 53340 7916 53344
rect 7852 53284 7856 53340
rect 7856 53284 7912 53340
rect 7912 53284 7916 53340
rect 7852 53280 7916 53284
rect 12612 53340 12676 53344
rect 12612 53284 12616 53340
rect 12616 53284 12672 53340
rect 12672 53284 12676 53340
rect 12612 53280 12676 53284
rect 12692 53340 12756 53344
rect 12692 53284 12696 53340
rect 12696 53284 12752 53340
rect 12752 53284 12756 53340
rect 12692 53280 12756 53284
rect 12772 53340 12836 53344
rect 12772 53284 12776 53340
rect 12776 53284 12832 53340
rect 12832 53284 12836 53340
rect 12772 53280 12836 53284
rect 12852 53340 12916 53344
rect 12852 53284 12856 53340
rect 12856 53284 12912 53340
rect 12912 53284 12916 53340
rect 12852 53280 12916 53284
rect 17612 53340 17676 53344
rect 17612 53284 17616 53340
rect 17616 53284 17672 53340
rect 17672 53284 17676 53340
rect 17612 53280 17676 53284
rect 17692 53340 17756 53344
rect 17692 53284 17696 53340
rect 17696 53284 17752 53340
rect 17752 53284 17756 53340
rect 17692 53280 17756 53284
rect 17772 53340 17836 53344
rect 17772 53284 17776 53340
rect 17776 53284 17832 53340
rect 17832 53284 17836 53340
rect 17772 53280 17836 53284
rect 17852 53340 17916 53344
rect 17852 53284 17856 53340
rect 17856 53284 17912 53340
rect 17912 53284 17916 53340
rect 17852 53280 17916 53284
rect 22612 53340 22676 53344
rect 22612 53284 22616 53340
rect 22616 53284 22672 53340
rect 22672 53284 22676 53340
rect 22612 53280 22676 53284
rect 22692 53340 22756 53344
rect 22692 53284 22696 53340
rect 22696 53284 22752 53340
rect 22752 53284 22756 53340
rect 22692 53280 22756 53284
rect 22772 53340 22836 53344
rect 22772 53284 22776 53340
rect 22776 53284 22832 53340
rect 22832 53284 22836 53340
rect 22772 53280 22836 53284
rect 22852 53340 22916 53344
rect 22852 53284 22856 53340
rect 22856 53284 22912 53340
rect 22912 53284 22916 53340
rect 22852 53280 22916 53284
rect 27612 53340 27676 53344
rect 27612 53284 27616 53340
rect 27616 53284 27672 53340
rect 27672 53284 27676 53340
rect 27612 53280 27676 53284
rect 27692 53340 27756 53344
rect 27692 53284 27696 53340
rect 27696 53284 27752 53340
rect 27752 53284 27756 53340
rect 27692 53280 27756 53284
rect 27772 53340 27836 53344
rect 27772 53284 27776 53340
rect 27776 53284 27832 53340
rect 27832 53284 27836 53340
rect 27772 53280 27836 53284
rect 27852 53340 27916 53344
rect 27852 53284 27856 53340
rect 27856 53284 27912 53340
rect 27912 53284 27916 53340
rect 27852 53280 27916 53284
rect 32612 53340 32676 53344
rect 32612 53284 32616 53340
rect 32616 53284 32672 53340
rect 32672 53284 32676 53340
rect 32612 53280 32676 53284
rect 32692 53340 32756 53344
rect 32692 53284 32696 53340
rect 32696 53284 32752 53340
rect 32752 53284 32756 53340
rect 32692 53280 32756 53284
rect 32772 53340 32836 53344
rect 32772 53284 32776 53340
rect 32776 53284 32832 53340
rect 32832 53284 32836 53340
rect 32772 53280 32836 53284
rect 32852 53340 32916 53344
rect 32852 53284 32856 53340
rect 32856 53284 32912 53340
rect 32912 53284 32916 53340
rect 32852 53280 32916 53284
rect 37612 53340 37676 53344
rect 37612 53284 37616 53340
rect 37616 53284 37672 53340
rect 37672 53284 37676 53340
rect 37612 53280 37676 53284
rect 37692 53340 37756 53344
rect 37692 53284 37696 53340
rect 37696 53284 37752 53340
rect 37752 53284 37756 53340
rect 37692 53280 37756 53284
rect 37772 53340 37836 53344
rect 37772 53284 37776 53340
rect 37776 53284 37832 53340
rect 37832 53284 37836 53340
rect 37772 53280 37836 53284
rect 37852 53340 37916 53344
rect 37852 53284 37856 53340
rect 37856 53284 37912 53340
rect 37912 53284 37916 53340
rect 37852 53280 37916 53284
rect 42612 53340 42676 53344
rect 42612 53284 42616 53340
rect 42616 53284 42672 53340
rect 42672 53284 42676 53340
rect 42612 53280 42676 53284
rect 42692 53340 42756 53344
rect 42692 53284 42696 53340
rect 42696 53284 42752 53340
rect 42752 53284 42756 53340
rect 42692 53280 42756 53284
rect 42772 53340 42836 53344
rect 42772 53284 42776 53340
rect 42776 53284 42832 53340
rect 42832 53284 42836 53340
rect 42772 53280 42836 53284
rect 42852 53340 42916 53344
rect 42852 53284 42856 53340
rect 42856 53284 42912 53340
rect 42912 53284 42916 53340
rect 42852 53280 42916 53284
rect 47612 53340 47676 53344
rect 47612 53284 47616 53340
rect 47616 53284 47672 53340
rect 47672 53284 47676 53340
rect 47612 53280 47676 53284
rect 47692 53340 47756 53344
rect 47692 53284 47696 53340
rect 47696 53284 47752 53340
rect 47752 53284 47756 53340
rect 47692 53280 47756 53284
rect 47772 53340 47836 53344
rect 47772 53284 47776 53340
rect 47776 53284 47832 53340
rect 47832 53284 47836 53340
rect 47772 53280 47836 53284
rect 47852 53340 47916 53344
rect 47852 53284 47856 53340
rect 47856 53284 47912 53340
rect 47912 53284 47916 53340
rect 47852 53280 47916 53284
rect 52612 53340 52676 53344
rect 52612 53284 52616 53340
rect 52616 53284 52672 53340
rect 52672 53284 52676 53340
rect 52612 53280 52676 53284
rect 52692 53340 52756 53344
rect 52692 53284 52696 53340
rect 52696 53284 52752 53340
rect 52752 53284 52756 53340
rect 52692 53280 52756 53284
rect 52772 53340 52836 53344
rect 52772 53284 52776 53340
rect 52776 53284 52832 53340
rect 52832 53284 52836 53340
rect 52772 53280 52836 53284
rect 52852 53340 52916 53344
rect 52852 53284 52856 53340
rect 52856 53284 52912 53340
rect 52912 53284 52916 53340
rect 52852 53280 52916 53284
rect 57612 53340 57676 53344
rect 57612 53284 57616 53340
rect 57616 53284 57672 53340
rect 57672 53284 57676 53340
rect 57612 53280 57676 53284
rect 57692 53340 57756 53344
rect 57692 53284 57696 53340
rect 57696 53284 57752 53340
rect 57752 53284 57756 53340
rect 57692 53280 57756 53284
rect 57772 53340 57836 53344
rect 57772 53284 57776 53340
rect 57776 53284 57832 53340
rect 57832 53284 57836 53340
rect 57772 53280 57836 53284
rect 57852 53340 57916 53344
rect 57852 53284 57856 53340
rect 57856 53284 57912 53340
rect 57912 53284 57916 53340
rect 57852 53280 57916 53284
rect 1952 52796 2016 52800
rect 1952 52740 1956 52796
rect 1956 52740 2012 52796
rect 2012 52740 2016 52796
rect 1952 52736 2016 52740
rect 2032 52796 2096 52800
rect 2032 52740 2036 52796
rect 2036 52740 2092 52796
rect 2092 52740 2096 52796
rect 2032 52736 2096 52740
rect 2112 52796 2176 52800
rect 2112 52740 2116 52796
rect 2116 52740 2172 52796
rect 2172 52740 2176 52796
rect 2112 52736 2176 52740
rect 2192 52796 2256 52800
rect 2192 52740 2196 52796
rect 2196 52740 2252 52796
rect 2252 52740 2256 52796
rect 2192 52736 2256 52740
rect 6952 52796 7016 52800
rect 6952 52740 6956 52796
rect 6956 52740 7012 52796
rect 7012 52740 7016 52796
rect 6952 52736 7016 52740
rect 7032 52796 7096 52800
rect 7032 52740 7036 52796
rect 7036 52740 7092 52796
rect 7092 52740 7096 52796
rect 7032 52736 7096 52740
rect 7112 52796 7176 52800
rect 7112 52740 7116 52796
rect 7116 52740 7172 52796
rect 7172 52740 7176 52796
rect 7112 52736 7176 52740
rect 7192 52796 7256 52800
rect 7192 52740 7196 52796
rect 7196 52740 7252 52796
rect 7252 52740 7256 52796
rect 7192 52736 7256 52740
rect 11952 52796 12016 52800
rect 11952 52740 11956 52796
rect 11956 52740 12012 52796
rect 12012 52740 12016 52796
rect 11952 52736 12016 52740
rect 12032 52796 12096 52800
rect 12032 52740 12036 52796
rect 12036 52740 12092 52796
rect 12092 52740 12096 52796
rect 12032 52736 12096 52740
rect 12112 52796 12176 52800
rect 12112 52740 12116 52796
rect 12116 52740 12172 52796
rect 12172 52740 12176 52796
rect 12112 52736 12176 52740
rect 12192 52796 12256 52800
rect 12192 52740 12196 52796
rect 12196 52740 12252 52796
rect 12252 52740 12256 52796
rect 12192 52736 12256 52740
rect 16952 52796 17016 52800
rect 16952 52740 16956 52796
rect 16956 52740 17012 52796
rect 17012 52740 17016 52796
rect 16952 52736 17016 52740
rect 17032 52796 17096 52800
rect 17032 52740 17036 52796
rect 17036 52740 17092 52796
rect 17092 52740 17096 52796
rect 17032 52736 17096 52740
rect 17112 52796 17176 52800
rect 17112 52740 17116 52796
rect 17116 52740 17172 52796
rect 17172 52740 17176 52796
rect 17112 52736 17176 52740
rect 17192 52796 17256 52800
rect 17192 52740 17196 52796
rect 17196 52740 17252 52796
rect 17252 52740 17256 52796
rect 17192 52736 17256 52740
rect 21952 52796 22016 52800
rect 21952 52740 21956 52796
rect 21956 52740 22012 52796
rect 22012 52740 22016 52796
rect 21952 52736 22016 52740
rect 22032 52796 22096 52800
rect 22032 52740 22036 52796
rect 22036 52740 22092 52796
rect 22092 52740 22096 52796
rect 22032 52736 22096 52740
rect 22112 52796 22176 52800
rect 22112 52740 22116 52796
rect 22116 52740 22172 52796
rect 22172 52740 22176 52796
rect 22112 52736 22176 52740
rect 22192 52796 22256 52800
rect 22192 52740 22196 52796
rect 22196 52740 22252 52796
rect 22252 52740 22256 52796
rect 22192 52736 22256 52740
rect 26952 52796 27016 52800
rect 26952 52740 26956 52796
rect 26956 52740 27012 52796
rect 27012 52740 27016 52796
rect 26952 52736 27016 52740
rect 27032 52796 27096 52800
rect 27032 52740 27036 52796
rect 27036 52740 27092 52796
rect 27092 52740 27096 52796
rect 27032 52736 27096 52740
rect 27112 52796 27176 52800
rect 27112 52740 27116 52796
rect 27116 52740 27172 52796
rect 27172 52740 27176 52796
rect 27112 52736 27176 52740
rect 27192 52796 27256 52800
rect 27192 52740 27196 52796
rect 27196 52740 27252 52796
rect 27252 52740 27256 52796
rect 27192 52736 27256 52740
rect 31952 52796 32016 52800
rect 31952 52740 31956 52796
rect 31956 52740 32012 52796
rect 32012 52740 32016 52796
rect 31952 52736 32016 52740
rect 32032 52796 32096 52800
rect 32032 52740 32036 52796
rect 32036 52740 32092 52796
rect 32092 52740 32096 52796
rect 32032 52736 32096 52740
rect 32112 52796 32176 52800
rect 32112 52740 32116 52796
rect 32116 52740 32172 52796
rect 32172 52740 32176 52796
rect 32112 52736 32176 52740
rect 32192 52796 32256 52800
rect 32192 52740 32196 52796
rect 32196 52740 32252 52796
rect 32252 52740 32256 52796
rect 32192 52736 32256 52740
rect 36952 52796 37016 52800
rect 36952 52740 36956 52796
rect 36956 52740 37012 52796
rect 37012 52740 37016 52796
rect 36952 52736 37016 52740
rect 37032 52796 37096 52800
rect 37032 52740 37036 52796
rect 37036 52740 37092 52796
rect 37092 52740 37096 52796
rect 37032 52736 37096 52740
rect 37112 52796 37176 52800
rect 37112 52740 37116 52796
rect 37116 52740 37172 52796
rect 37172 52740 37176 52796
rect 37112 52736 37176 52740
rect 37192 52796 37256 52800
rect 37192 52740 37196 52796
rect 37196 52740 37252 52796
rect 37252 52740 37256 52796
rect 37192 52736 37256 52740
rect 41952 52796 42016 52800
rect 41952 52740 41956 52796
rect 41956 52740 42012 52796
rect 42012 52740 42016 52796
rect 41952 52736 42016 52740
rect 42032 52796 42096 52800
rect 42032 52740 42036 52796
rect 42036 52740 42092 52796
rect 42092 52740 42096 52796
rect 42032 52736 42096 52740
rect 42112 52796 42176 52800
rect 42112 52740 42116 52796
rect 42116 52740 42172 52796
rect 42172 52740 42176 52796
rect 42112 52736 42176 52740
rect 42192 52796 42256 52800
rect 42192 52740 42196 52796
rect 42196 52740 42252 52796
rect 42252 52740 42256 52796
rect 42192 52736 42256 52740
rect 46952 52796 47016 52800
rect 46952 52740 46956 52796
rect 46956 52740 47012 52796
rect 47012 52740 47016 52796
rect 46952 52736 47016 52740
rect 47032 52796 47096 52800
rect 47032 52740 47036 52796
rect 47036 52740 47092 52796
rect 47092 52740 47096 52796
rect 47032 52736 47096 52740
rect 47112 52796 47176 52800
rect 47112 52740 47116 52796
rect 47116 52740 47172 52796
rect 47172 52740 47176 52796
rect 47112 52736 47176 52740
rect 47192 52796 47256 52800
rect 47192 52740 47196 52796
rect 47196 52740 47252 52796
rect 47252 52740 47256 52796
rect 47192 52736 47256 52740
rect 51952 52796 52016 52800
rect 51952 52740 51956 52796
rect 51956 52740 52012 52796
rect 52012 52740 52016 52796
rect 51952 52736 52016 52740
rect 52032 52796 52096 52800
rect 52032 52740 52036 52796
rect 52036 52740 52092 52796
rect 52092 52740 52096 52796
rect 52032 52736 52096 52740
rect 52112 52796 52176 52800
rect 52112 52740 52116 52796
rect 52116 52740 52172 52796
rect 52172 52740 52176 52796
rect 52112 52736 52176 52740
rect 52192 52796 52256 52800
rect 52192 52740 52196 52796
rect 52196 52740 52252 52796
rect 52252 52740 52256 52796
rect 52192 52736 52256 52740
rect 56952 52796 57016 52800
rect 56952 52740 56956 52796
rect 56956 52740 57012 52796
rect 57012 52740 57016 52796
rect 56952 52736 57016 52740
rect 57032 52796 57096 52800
rect 57032 52740 57036 52796
rect 57036 52740 57092 52796
rect 57092 52740 57096 52796
rect 57032 52736 57096 52740
rect 57112 52796 57176 52800
rect 57112 52740 57116 52796
rect 57116 52740 57172 52796
rect 57172 52740 57176 52796
rect 57112 52736 57176 52740
rect 57192 52796 57256 52800
rect 57192 52740 57196 52796
rect 57196 52740 57252 52796
rect 57252 52740 57256 52796
rect 57192 52736 57256 52740
rect 2612 52252 2676 52256
rect 2612 52196 2616 52252
rect 2616 52196 2672 52252
rect 2672 52196 2676 52252
rect 2612 52192 2676 52196
rect 2692 52252 2756 52256
rect 2692 52196 2696 52252
rect 2696 52196 2752 52252
rect 2752 52196 2756 52252
rect 2692 52192 2756 52196
rect 2772 52252 2836 52256
rect 2772 52196 2776 52252
rect 2776 52196 2832 52252
rect 2832 52196 2836 52252
rect 2772 52192 2836 52196
rect 2852 52252 2916 52256
rect 2852 52196 2856 52252
rect 2856 52196 2912 52252
rect 2912 52196 2916 52252
rect 2852 52192 2916 52196
rect 7612 52252 7676 52256
rect 7612 52196 7616 52252
rect 7616 52196 7672 52252
rect 7672 52196 7676 52252
rect 7612 52192 7676 52196
rect 7692 52252 7756 52256
rect 7692 52196 7696 52252
rect 7696 52196 7752 52252
rect 7752 52196 7756 52252
rect 7692 52192 7756 52196
rect 7772 52252 7836 52256
rect 7772 52196 7776 52252
rect 7776 52196 7832 52252
rect 7832 52196 7836 52252
rect 7772 52192 7836 52196
rect 7852 52252 7916 52256
rect 7852 52196 7856 52252
rect 7856 52196 7912 52252
rect 7912 52196 7916 52252
rect 7852 52192 7916 52196
rect 12612 52252 12676 52256
rect 12612 52196 12616 52252
rect 12616 52196 12672 52252
rect 12672 52196 12676 52252
rect 12612 52192 12676 52196
rect 12692 52252 12756 52256
rect 12692 52196 12696 52252
rect 12696 52196 12752 52252
rect 12752 52196 12756 52252
rect 12692 52192 12756 52196
rect 12772 52252 12836 52256
rect 12772 52196 12776 52252
rect 12776 52196 12832 52252
rect 12832 52196 12836 52252
rect 12772 52192 12836 52196
rect 12852 52252 12916 52256
rect 12852 52196 12856 52252
rect 12856 52196 12912 52252
rect 12912 52196 12916 52252
rect 12852 52192 12916 52196
rect 17612 52252 17676 52256
rect 17612 52196 17616 52252
rect 17616 52196 17672 52252
rect 17672 52196 17676 52252
rect 17612 52192 17676 52196
rect 17692 52252 17756 52256
rect 17692 52196 17696 52252
rect 17696 52196 17752 52252
rect 17752 52196 17756 52252
rect 17692 52192 17756 52196
rect 17772 52252 17836 52256
rect 17772 52196 17776 52252
rect 17776 52196 17832 52252
rect 17832 52196 17836 52252
rect 17772 52192 17836 52196
rect 17852 52252 17916 52256
rect 17852 52196 17856 52252
rect 17856 52196 17912 52252
rect 17912 52196 17916 52252
rect 17852 52192 17916 52196
rect 22612 52252 22676 52256
rect 22612 52196 22616 52252
rect 22616 52196 22672 52252
rect 22672 52196 22676 52252
rect 22612 52192 22676 52196
rect 22692 52252 22756 52256
rect 22692 52196 22696 52252
rect 22696 52196 22752 52252
rect 22752 52196 22756 52252
rect 22692 52192 22756 52196
rect 22772 52252 22836 52256
rect 22772 52196 22776 52252
rect 22776 52196 22832 52252
rect 22832 52196 22836 52252
rect 22772 52192 22836 52196
rect 22852 52252 22916 52256
rect 22852 52196 22856 52252
rect 22856 52196 22912 52252
rect 22912 52196 22916 52252
rect 22852 52192 22916 52196
rect 27612 52252 27676 52256
rect 27612 52196 27616 52252
rect 27616 52196 27672 52252
rect 27672 52196 27676 52252
rect 27612 52192 27676 52196
rect 27692 52252 27756 52256
rect 27692 52196 27696 52252
rect 27696 52196 27752 52252
rect 27752 52196 27756 52252
rect 27692 52192 27756 52196
rect 27772 52252 27836 52256
rect 27772 52196 27776 52252
rect 27776 52196 27832 52252
rect 27832 52196 27836 52252
rect 27772 52192 27836 52196
rect 27852 52252 27916 52256
rect 27852 52196 27856 52252
rect 27856 52196 27912 52252
rect 27912 52196 27916 52252
rect 27852 52192 27916 52196
rect 32612 52252 32676 52256
rect 32612 52196 32616 52252
rect 32616 52196 32672 52252
rect 32672 52196 32676 52252
rect 32612 52192 32676 52196
rect 32692 52252 32756 52256
rect 32692 52196 32696 52252
rect 32696 52196 32752 52252
rect 32752 52196 32756 52252
rect 32692 52192 32756 52196
rect 32772 52252 32836 52256
rect 32772 52196 32776 52252
rect 32776 52196 32832 52252
rect 32832 52196 32836 52252
rect 32772 52192 32836 52196
rect 32852 52252 32916 52256
rect 32852 52196 32856 52252
rect 32856 52196 32912 52252
rect 32912 52196 32916 52252
rect 32852 52192 32916 52196
rect 37612 52252 37676 52256
rect 37612 52196 37616 52252
rect 37616 52196 37672 52252
rect 37672 52196 37676 52252
rect 37612 52192 37676 52196
rect 37692 52252 37756 52256
rect 37692 52196 37696 52252
rect 37696 52196 37752 52252
rect 37752 52196 37756 52252
rect 37692 52192 37756 52196
rect 37772 52252 37836 52256
rect 37772 52196 37776 52252
rect 37776 52196 37832 52252
rect 37832 52196 37836 52252
rect 37772 52192 37836 52196
rect 37852 52252 37916 52256
rect 37852 52196 37856 52252
rect 37856 52196 37912 52252
rect 37912 52196 37916 52252
rect 37852 52192 37916 52196
rect 42612 52252 42676 52256
rect 42612 52196 42616 52252
rect 42616 52196 42672 52252
rect 42672 52196 42676 52252
rect 42612 52192 42676 52196
rect 42692 52252 42756 52256
rect 42692 52196 42696 52252
rect 42696 52196 42752 52252
rect 42752 52196 42756 52252
rect 42692 52192 42756 52196
rect 42772 52252 42836 52256
rect 42772 52196 42776 52252
rect 42776 52196 42832 52252
rect 42832 52196 42836 52252
rect 42772 52192 42836 52196
rect 42852 52252 42916 52256
rect 42852 52196 42856 52252
rect 42856 52196 42912 52252
rect 42912 52196 42916 52252
rect 42852 52192 42916 52196
rect 47612 52252 47676 52256
rect 47612 52196 47616 52252
rect 47616 52196 47672 52252
rect 47672 52196 47676 52252
rect 47612 52192 47676 52196
rect 47692 52252 47756 52256
rect 47692 52196 47696 52252
rect 47696 52196 47752 52252
rect 47752 52196 47756 52252
rect 47692 52192 47756 52196
rect 47772 52252 47836 52256
rect 47772 52196 47776 52252
rect 47776 52196 47832 52252
rect 47832 52196 47836 52252
rect 47772 52192 47836 52196
rect 47852 52252 47916 52256
rect 47852 52196 47856 52252
rect 47856 52196 47912 52252
rect 47912 52196 47916 52252
rect 47852 52192 47916 52196
rect 52612 52252 52676 52256
rect 52612 52196 52616 52252
rect 52616 52196 52672 52252
rect 52672 52196 52676 52252
rect 52612 52192 52676 52196
rect 52692 52252 52756 52256
rect 52692 52196 52696 52252
rect 52696 52196 52752 52252
rect 52752 52196 52756 52252
rect 52692 52192 52756 52196
rect 52772 52252 52836 52256
rect 52772 52196 52776 52252
rect 52776 52196 52832 52252
rect 52832 52196 52836 52252
rect 52772 52192 52836 52196
rect 52852 52252 52916 52256
rect 52852 52196 52856 52252
rect 52856 52196 52912 52252
rect 52912 52196 52916 52252
rect 52852 52192 52916 52196
rect 57612 52252 57676 52256
rect 57612 52196 57616 52252
rect 57616 52196 57672 52252
rect 57672 52196 57676 52252
rect 57612 52192 57676 52196
rect 57692 52252 57756 52256
rect 57692 52196 57696 52252
rect 57696 52196 57752 52252
rect 57752 52196 57756 52252
rect 57692 52192 57756 52196
rect 57772 52252 57836 52256
rect 57772 52196 57776 52252
rect 57776 52196 57832 52252
rect 57832 52196 57836 52252
rect 57772 52192 57836 52196
rect 57852 52252 57916 52256
rect 57852 52196 57856 52252
rect 57856 52196 57912 52252
rect 57912 52196 57916 52252
rect 57852 52192 57916 52196
rect 1952 51708 2016 51712
rect 1952 51652 1956 51708
rect 1956 51652 2012 51708
rect 2012 51652 2016 51708
rect 1952 51648 2016 51652
rect 2032 51708 2096 51712
rect 2032 51652 2036 51708
rect 2036 51652 2092 51708
rect 2092 51652 2096 51708
rect 2032 51648 2096 51652
rect 2112 51708 2176 51712
rect 2112 51652 2116 51708
rect 2116 51652 2172 51708
rect 2172 51652 2176 51708
rect 2112 51648 2176 51652
rect 2192 51708 2256 51712
rect 2192 51652 2196 51708
rect 2196 51652 2252 51708
rect 2252 51652 2256 51708
rect 2192 51648 2256 51652
rect 6952 51708 7016 51712
rect 6952 51652 6956 51708
rect 6956 51652 7012 51708
rect 7012 51652 7016 51708
rect 6952 51648 7016 51652
rect 7032 51708 7096 51712
rect 7032 51652 7036 51708
rect 7036 51652 7092 51708
rect 7092 51652 7096 51708
rect 7032 51648 7096 51652
rect 7112 51708 7176 51712
rect 7112 51652 7116 51708
rect 7116 51652 7172 51708
rect 7172 51652 7176 51708
rect 7112 51648 7176 51652
rect 7192 51708 7256 51712
rect 7192 51652 7196 51708
rect 7196 51652 7252 51708
rect 7252 51652 7256 51708
rect 7192 51648 7256 51652
rect 11952 51708 12016 51712
rect 11952 51652 11956 51708
rect 11956 51652 12012 51708
rect 12012 51652 12016 51708
rect 11952 51648 12016 51652
rect 12032 51708 12096 51712
rect 12032 51652 12036 51708
rect 12036 51652 12092 51708
rect 12092 51652 12096 51708
rect 12032 51648 12096 51652
rect 12112 51708 12176 51712
rect 12112 51652 12116 51708
rect 12116 51652 12172 51708
rect 12172 51652 12176 51708
rect 12112 51648 12176 51652
rect 12192 51708 12256 51712
rect 12192 51652 12196 51708
rect 12196 51652 12252 51708
rect 12252 51652 12256 51708
rect 12192 51648 12256 51652
rect 16952 51708 17016 51712
rect 16952 51652 16956 51708
rect 16956 51652 17012 51708
rect 17012 51652 17016 51708
rect 16952 51648 17016 51652
rect 17032 51708 17096 51712
rect 17032 51652 17036 51708
rect 17036 51652 17092 51708
rect 17092 51652 17096 51708
rect 17032 51648 17096 51652
rect 17112 51708 17176 51712
rect 17112 51652 17116 51708
rect 17116 51652 17172 51708
rect 17172 51652 17176 51708
rect 17112 51648 17176 51652
rect 17192 51708 17256 51712
rect 17192 51652 17196 51708
rect 17196 51652 17252 51708
rect 17252 51652 17256 51708
rect 17192 51648 17256 51652
rect 21952 51708 22016 51712
rect 21952 51652 21956 51708
rect 21956 51652 22012 51708
rect 22012 51652 22016 51708
rect 21952 51648 22016 51652
rect 22032 51708 22096 51712
rect 22032 51652 22036 51708
rect 22036 51652 22092 51708
rect 22092 51652 22096 51708
rect 22032 51648 22096 51652
rect 22112 51708 22176 51712
rect 22112 51652 22116 51708
rect 22116 51652 22172 51708
rect 22172 51652 22176 51708
rect 22112 51648 22176 51652
rect 22192 51708 22256 51712
rect 22192 51652 22196 51708
rect 22196 51652 22252 51708
rect 22252 51652 22256 51708
rect 22192 51648 22256 51652
rect 26952 51708 27016 51712
rect 26952 51652 26956 51708
rect 26956 51652 27012 51708
rect 27012 51652 27016 51708
rect 26952 51648 27016 51652
rect 27032 51708 27096 51712
rect 27032 51652 27036 51708
rect 27036 51652 27092 51708
rect 27092 51652 27096 51708
rect 27032 51648 27096 51652
rect 27112 51708 27176 51712
rect 27112 51652 27116 51708
rect 27116 51652 27172 51708
rect 27172 51652 27176 51708
rect 27112 51648 27176 51652
rect 27192 51708 27256 51712
rect 27192 51652 27196 51708
rect 27196 51652 27252 51708
rect 27252 51652 27256 51708
rect 27192 51648 27256 51652
rect 31952 51708 32016 51712
rect 31952 51652 31956 51708
rect 31956 51652 32012 51708
rect 32012 51652 32016 51708
rect 31952 51648 32016 51652
rect 32032 51708 32096 51712
rect 32032 51652 32036 51708
rect 32036 51652 32092 51708
rect 32092 51652 32096 51708
rect 32032 51648 32096 51652
rect 32112 51708 32176 51712
rect 32112 51652 32116 51708
rect 32116 51652 32172 51708
rect 32172 51652 32176 51708
rect 32112 51648 32176 51652
rect 32192 51708 32256 51712
rect 32192 51652 32196 51708
rect 32196 51652 32252 51708
rect 32252 51652 32256 51708
rect 32192 51648 32256 51652
rect 36952 51708 37016 51712
rect 36952 51652 36956 51708
rect 36956 51652 37012 51708
rect 37012 51652 37016 51708
rect 36952 51648 37016 51652
rect 37032 51708 37096 51712
rect 37032 51652 37036 51708
rect 37036 51652 37092 51708
rect 37092 51652 37096 51708
rect 37032 51648 37096 51652
rect 37112 51708 37176 51712
rect 37112 51652 37116 51708
rect 37116 51652 37172 51708
rect 37172 51652 37176 51708
rect 37112 51648 37176 51652
rect 37192 51708 37256 51712
rect 37192 51652 37196 51708
rect 37196 51652 37252 51708
rect 37252 51652 37256 51708
rect 37192 51648 37256 51652
rect 41952 51708 42016 51712
rect 41952 51652 41956 51708
rect 41956 51652 42012 51708
rect 42012 51652 42016 51708
rect 41952 51648 42016 51652
rect 42032 51708 42096 51712
rect 42032 51652 42036 51708
rect 42036 51652 42092 51708
rect 42092 51652 42096 51708
rect 42032 51648 42096 51652
rect 42112 51708 42176 51712
rect 42112 51652 42116 51708
rect 42116 51652 42172 51708
rect 42172 51652 42176 51708
rect 42112 51648 42176 51652
rect 42192 51708 42256 51712
rect 42192 51652 42196 51708
rect 42196 51652 42252 51708
rect 42252 51652 42256 51708
rect 42192 51648 42256 51652
rect 46952 51708 47016 51712
rect 46952 51652 46956 51708
rect 46956 51652 47012 51708
rect 47012 51652 47016 51708
rect 46952 51648 47016 51652
rect 47032 51708 47096 51712
rect 47032 51652 47036 51708
rect 47036 51652 47092 51708
rect 47092 51652 47096 51708
rect 47032 51648 47096 51652
rect 47112 51708 47176 51712
rect 47112 51652 47116 51708
rect 47116 51652 47172 51708
rect 47172 51652 47176 51708
rect 47112 51648 47176 51652
rect 47192 51708 47256 51712
rect 47192 51652 47196 51708
rect 47196 51652 47252 51708
rect 47252 51652 47256 51708
rect 47192 51648 47256 51652
rect 51952 51708 52016 51712
rect 51952 51652 51956 51708
rect 51956 51652 52012 51708
rect 52012 51652 52016 51708
rect 51952 51648 52016 51652
rect 52032 51708 52096 51712
rect 52032 51652 52036 51708
rect 52036 51652 52092 51708
rect 52092 51652 52096 51708
rect 52032 51648 52096 51652
rect 52112 51708 52176 51712
rect 52112 51652 52116 51708
rect 52116 51652 52172 51708
rect 52172 51652 52176 51708
rect 52112 51648 52176 51652
rect 52192 51708 52256 51712
rect 52192 51652 52196 51708
rect 52196 51652 52252 51708
rect 52252 51652 52256 51708
rect 52192 51648 52256 51652
rect 56952 51708 57016 51712
rect 56952 51652 56956 51708
rect 56956 51652 57012 51708
rect 57012 51652 57016 51708
rect 56952 51648 57016 51652
rect 57032 51708 57096 51712
rect 57032 51652 57036 51708
rect 57036 51652 57092 51708
rect 57092 51652 57096 51708
rect 57032 51648 57096 51652
rect 57112 51708 57176 51712
rect 57112 51652 57116 51708
rect 57116 51652 57172 51708
rect 57172 51652 57176 51708
rect 57112 51648 57176 51652
rect 57192 51708 57256 51712
rect 57192 51652 57196 51708
rect 57196 51652 57252 51708
rect 57252 51652 57256 51708
rect 57192 51648 57256 51652
rect 2612 51164 2676 51168
rect 2612 51108 2616 51164
rect 2616 51108 2672 51164
rect 2672 51108 2676 51164
rect 2612 51104 2676 51108
rect 2692 51164 2756 51168
rect 2692 51108 2696 51164
rect 2696 51108 2752 51164
rect 2752 51108 2756 51164
rect 2692 51104 2756 51108
rect 2772 51164 2836 51168
rect 2772 51108 2776 51164
rect 2776 51108 2832 51164
rect 2832 51108 2836 51164
rect 2772 51104 2836 51108
rect 2852 51164 2916 51168
rect 2852 51108 2856 51164
rect 2856 51108 2912 51164
rect 2912 51108 2916 51164
rect 2852 51104 2916 51108
rect 7612 51164 7676 51168
rect 7612 51108 7616 51164
rect 7616 51108 7672 51164
rect 7672 51108 7676 51164
rect 7612 51104 7676 51108
rect 7692 51164 7756 51168
rect 7692 51108 7696 51164
rect 7696 51108 7752 51164
rect 7752 51108 7756 51164
rect 7692 51104 7756 51108
rect 7772 51164 7836 51168
rect 7772 51108 7776 51164
rect 7776 51108 7832 51164
rect 7832 51108 7836 51164
rect 7772 51104 7836 51108
rect 7852 51164 7916 51168
rect 7852 51108 7856 51164
rect 7856 51108 7912 51164
rect 7912 51108 7916 51164
rect 7852 51104 7916 51108
rect 12612 51164 12676 51168
rect 12612 51108 12616 51164
rect 12616 51108 12672 51164
rect 12672 51108 12676 51164
rect 12612 51104 12676 51108
rect 12692 51164 12756 51168
rect 12692 51108 12696 51164
rect 12696 51108 12752 51164
rect 12752 51108 12756 51164
rect 12692 51104 12756 51108
rect 12772 51164 12836 51168
rect 12772 51108 12776 51164
rect 12776 51108 12832 51164
rect 12832 51108 12836 51164
rect 12772 51104 12836 51108
rect 12852 51164 12916 51168
rect 12852 51108 12856 51164
rect 12856 51108 12912 51164
rect 12912 51108 12916 51164
rect 12852 51104 12916 51108
rect 17612 51164 17676 51168
rect 17612 51108 17616 51164
rect 17616 51108 17672 51164
rect 17672 51108 17676 51164
rect 17612 51104 17676 51108
rect 17692 51164 17756 51168
rect 17692 51108 17696 51164
rect 17696 51108 17752 51164
rect 17752 51108 17756 51164
rect 17692 51104 17756 51108
rect 17772 51164 17836 51168
rect 17772 51108 17776 51164
rect 17776 51108 17832 51164
rect 17832 51108 17836 51164
rect 17772 51104 17836 51108
rect 17852 51164 17916 51168
rect 17852 51108 17856 51164
rect 17856 51108 17912 51164
rect 17912 51108 17916 51164
rect 17852 51104 17916 51108
rect 22612 51164 22676 51168
rect 22612 51108 22616 51164
rect 22616 51108 22672 51164
rect 22672 51108 22676 51164
rect 22612 51104 22676 51108
rect 22692 51164 22756 51168
rect 22692 51108 22696 51164
rect 22696 51108 22752 51164
rect 22752 51108 22756 51164
rect 22692 51104 22756 51108
rect 22772 51164 22836 51168
rect 22772 51108 22776 51164
rect 22776 51108 22832 51164
rect 22832 51108 22836 51164
rect 22772 51104 22836 51108
rect 22852 51164 22916 51168
rect 22852 51108 22856 51164
rect 22856 51108 22912 51164
rect 22912 51108 22916 51164
rect 22852 51104 22916 51108
rect 27612 51164 27676 51168
rect 27612 51108 27616 51164
rect 27616 51108 27672 51164
rect 27672 51108 27676 51164
rect 27612 51104 27676 51108
rect 27692 51164 27756 51168
rect 27692 51108 27696 51164
rect 27696 51108 27752 51164
rect 27752 51108 27756 51164
rect 27692 51104 27756 51108
rect 27772 51164 27836 51168
rect 27772 51108 27776 51164
rect 27776 51108 27832 51164
rect 27832 51108 27836 51164
rect 27772 51104 27836 51108
rect 27852 51164 27916 51168
rect 27852 51108 27856 51164
rect 27856 51108 27912 51164
rect 27912 51108 27916 51164
rect 27852 51104 27916 51108
rect 32612 51164 32676 51168
rect 32612 51108 32616 51164
rect 32616 51108 32672 51164
rect 32672 51108 32676 51164
rect 32612 51104 32676 51108
rect 32692 51164 32756 51168
rect 32692 51108 32696 51164
rect 32696 51108 32752 51164
rect 32752 51108 32756 51164
rect 32692 51104 32756 51108
rect 32772 51164 32836 51168
rect 32772 51108 32776 51164
rect 32776 51108 32832 51164
rect 32832 51108 32836 51164
rect 32772 51104 32836 51108
rect 32852 51164 32916 51168
rect 32852 51108 32856 51164
rect 32856 51108 32912 51164
rect 32912 51108 32916 51164
rect 32852 51104 32916 51108
rect 37612 51164 37676 51168
rect 37612 51108 37616 51164
rect 37616 51108 37672 51164
rect 37672 51108 37676 51164
rect 37612 51104 37676 51108
rect 37692 51164 37756 51168
rect 37692 51108 37696 51164
rect 37696 51108 37752 51164
rect 37752 51108 37756 51164
rect 37692 51104 37756 51108
rect 37772 51164 37836 51168
rect 37772 51108 37776 51164
rect 37776 51108 37832 51164
rect 37832 51108 37836 51164
rect 37772 51104 37836 51108
rect 37852 51164 37916 51168
rect 37852 51108 37856 51164
rect 37856 51108 37912 51164
rect 37912 51108 37916 51164
rect 37852 51104 37916 51108
rect 42612 51164 42676 51168
rect 42612 51108 42616 51164
rect 42616 51108 42672 51164
rect 42672 51108 42676 51164
rect 42612 51104 42676 51108
rect 42692 51164 42756 51168
rect 42692 51108 42696 51164
rect 42696 51108 42752 51164
rect 42752 51108 42756 51164
rect 42692 51104 42756 51108
rect 42772 51164 42836 51168
rect 42772 51108 42776 51164
rect 42776 51108 42832 51164
rect 42832 51108 42836 51164
rect 42772 51104 42836 51108
rect 42852 51164 42916 51168
rect 42852 51108 42856 51164
rect 42856 51108 42912 51164
rect 42912 51108 42916 51164
rect 42852 51104 42916 51108
rect 47612 51164 47676 51168
rect 47612 51108 47616 51164
rect 47616 51108 47672 51164
rect 47672 51108 47676 51164
rect 47612 51104 47676 51108
rect 47692 51164 47756 51168
rect 47692 51108 47696 51164
rect 47696 51108 47752 51164
rect 47752 51108 47756 51164
rect 47692 51104 47756 51108
rect 47772 51164 47836 51168
rect 47772 51108 47776 51164
rect 47776 51108 47832 51164
rect 47832 51108 47836 51164
rect 47772 51104 47836 51108
rect 47852 51164 47916 51168
rect 47852 51108 47856 51164
rect 47856 51108 47912 51164
rect 47912 51108 47916 51164
rect 47852 51104 47916 51108
rect 52612 51164 52676 51168
rect 52612 51108 52616 51164
rect 52616 51108 52672 51164
rect 52672 51108 52676 51164
rect 52612 51104 52676 51108
rect 52692 51164 52756 51168
rect 52692 51108 52696 51164
rect 52696 51108 52752 51164
rect 52752 51108 52756 51164
rect 52692 51104 52756 51108
rect 52772 51164 52836 51168
rect 52772 51108 52776 51164
rect 52776 51108 52832 51164
rect 52832 51108 52836 51164
rect 52772 51104 52836 51108
rect 52852 51164 52916 51168
rect 52852 51108 52856 51164
rect 52856 51108 52912 51164
rect 52912 51108 52916 51164
rect 52852 51104 52916 51108
rect 57612 51164 57676 51168
rect 57612 51108 57616 51164
rect 57616 51108 57672 51164
rect 57672 51108 57676 51164
rect 57612 51104 57676 51108
rect 57692 51164 57756 51168
rect 57692 51108 57696 51164
rect 57696 51108 57752 51164
rect 57752 51108 57756 51164
rect 57692 51104 57756 51108
rect 57772 51164 57836 51168
rect 57772 51108 57776 51164
rect 57776 51108 57832 51164
rect 57832 51108 57836 51164
rect 57772 51104 57836 51108
rect 57852 51164 57916 51168
rect 57852 51108 57856 51164
rect 57856 51108 57912 51164
rect 57912 51108 57916 51164
rect 57852 51104 57916 51108
rect 1952 50620 2016 50624
rect 1952 50564 1956 50620
rect 1956 50564 2012 50620
rect 2012 50564 2016 50620
rect 1952 50560 2016 50564
rect 2032 50620 2096 50624
rect 2032 50564 2036 50620
rect 2036 50564 2092 50620
rect 2092 50564 2096 50620
rect 2032 50560 2096 50564
rect 2112 50620 2176 50624
rect 2112 50564 2116 50620
rect 2116 50564 2172 50620
rect 2172 50564 2176 50620
rect 2112 50560 2176 50564
rect 2192 50620 2256 50624
rect 2192 50564 2196 50620
rect 2196 50564 2252 50620
rect 2252 50564 2256 50620
rect 2192 50560 2256 50564
rect 6952 50620 7016 50624
rect 6952 50564 6956 50620
rect 6956 50564 7012 50620
rect 7012 50564 7016 50620
rect 6952 50560 7016 50564
rect 7032 50620 7096 50624
rect 7032 50564 7036 50620
rect 7036 50564 7092 50620
rect 7092 50564 7096 50620
rect 7032 50560 7096 50564
rect 7112 50620 7176 50624
rect 7112 50564 7116 50620
rect 7116 50564 7172 50620
rect 7172 50564 7176 50620
rect 7112 50560 7176 50564
rect 7192 50620 7256 50624
rect 7192 50564 7196 50620
rect 7196 50564 7252 50620
rect 7252 50564 7256 50620
rect 7192 50560 7256 50564
rect 11952 50620 12016 50624
rect 11952 50564 11956 50620
rect 11956 50564 12012 50620
rect 12012 50564 12016 50620
rect 11952 50560 12016 50564
rect 12032 50620 12096 50624
rect 12032 50564 12036 50620
rect 12036 50564 12092 50620
rect 12092 50564 12096 50620
rect 12032 50560 12096 50564
rect 12112 50620 12176 50624
rect 12112 50564 12116 50620
rect 12116 50564 12172 50620
rect 12172 50564 12176 50620
rect 12112 50560 12176 50564
rect 12192 50620 12256 50624
rect 12192 50564 12196 50620
rect 12196 50564 12252 50620
rect 12252 50564 12256 50620
rect 12192 50560 12256 50564
rect 16952 50620 17016 50624
rect 16952 50564 16956 50620
rect 16956 50564 17012 50620
rect 17012 50564 17016 50620
rect 16952 50560 17016 50564
rect 17032 50620 17096 50624
rect 17032 50564 17036 50620
rect 17036 50564 17092 50620
rect 17092 50564 17096 50620
rect 17032 50560 17096 50564
rect 17112 50620 17176 50624
rect 17112 50564 17116 50620
rect 17116 50564 17172 50620
rect 17172 50564 17176 50620
rect 17112 50560 17176 50564
rect 17192 50620 17256 50624
rect 17192 50564 17196 50620
rect 17196 50564 17252 50620
rect 17252 50564 17256 50620
rect 17192 50560 17256 50564
rect 21952 50620 22016 50624
rect 21952 50564 21956 50620
rect 21956 50564 22012 50620
rect 22012 50564 22016 50620
rect 21952 50560 22016 50564
rect 22032 50620 22096 50624
rect 22032 50564 22036 50620
rect 22036 50564 22092 50620
rect 22092 50564 22096 50620
rect 22032 50560 22096 50564
rect 22112 50620 22176 50624
rect 22112 50564 22116 50620
rect 22116 50564 22172 50620
rect 22172 50564 22176 50620
rect 22112 50560 22176 50564
rect 22192 50620 22256 50624
rect 22192 50564 22196 50620
rect 22196 50564 22252 50620
rect 22252 50564 22256 50620
rect 22192 50560 22256 50564
rect 26952 50620 27016 50624
rect 26952 50564 26956 50620
rect 26956 50564 27012 50620
rect 27012 50564 27016 50620
rect 26952 50560 27016 50564
rect 27032 50620 27096 50624
rect 27032 50564 27036 50620
rect 27036 50564 27092 50620
rect 27092 50564 27096 50620
rect 27032 50560 27096 50564
rect 27112 50620 27176 50624
rect 27112 50564 27116 50620
rect 27116 50564 27172 50620
rect 27172 50564 27176 50620
rect 27112 50560 27176 50564
rect 27192 50620 27256 50624
rect 27192 50564 27196 50620
rect 27196 50564 27252 50620
rect 27252 50564 27256 50620
rect 27192 50560 27256 50564
rect 31952 50620 32016 50624
rect 31952 50564 31956 50620
rect 31956 50564 32012 50620
rect 32012 50564 32016 50620
rect 31952 50560 32016 50564
rect 32032 50620 32096 50624
rect 32032 50564 32036 50620
rect 32036 50564 32092 50620
rect 32092 50564 32096 50620
rect 32032 50560 32096 50564
rect 32112 50620 32176 50624
rect 32112 50564 32116 50620
rect 32116 50564 32172 50620
rect 32172 50564 32176 50620
rect 32112 50560 32176 50564
rect 32192 50620 32256 50624
rect 32192 50564 32196 50620
rect 32196 50564 32252 50620
rect 32252 50564 32256 50620
rect 32192 50560 32256 50564
rect 36952 50620 37016 50624
rect 36952 50564 36956 50620
rect 36956 50564 37012 50620
rect 37012 50564 37016 50620
rect 36952 50560 37016 50564
rect 37032 50620 37096 50624
rect 37032 50564 37036 50620
rect 37036 50564 37092 50620
rect 37092 50564 37096 50620
rect 37032 50560 37096 50564
rect 37112 50620 37176 50624
rect 37112 50564 37116 50620
rect 37116 50564 37172 50620
rect 37172 50564 37176 50620
rect 37112 50560 37176 50564
rect 37192 50620 37256 50624
rect 37192 50564 37196 50620
rect 37196 50564 37252 50620
rect 37252 50564 37256 50620
rect 37192 50560 37256 50564
rect 41952 50620 42016 50624
rect 41952 50564 41956 50620
rect 41956 50564 42012 50620
rect 42012 50564 42016 50620
rect 41952 50560 42016 50564
rect 42032 50620 42096 50624
rect 42032 50564 42036 50620
rect 42036 50564 42092 50620
rect 42092 50564 42096 50620
rect 42032 50560 42096 50564
rect 42112 50620 42176 50624
rect 42112 50564 42116 50620
rect 42116 50564 42172 50620
rect 42172 50564 42176 50620
rect 42112 50560 42176 50564
rect 42192 50620 42256 50624
rect 42192 50564 42196 50620
rect 42196 50564 42252 50620
rect 42252 50564 42256 50620
rect 42192 50560 42256 50564
rect 46952 50620 47016 50624
rect 46952 50564 46956 50620
rect 46956 50564 47012 50620
rect 47012 50564 47016 50620
rect 46952 50560 47016 50564
rect 47032 50620 47096 50624
rect 47032 50564 47036 50620
rect 47036 50564 47092 50620
rect 47092 50564 47096 50620
rect 47032 50560 47096 50564
rect 47112 50620 47176 50624
rect 47112 50564 47116 50620
rect 47116 50564 47172 50620
rect 47172 50564 47176 50620
rect 47112 50560 47176 50564
rect 47192 50620 47256 50624
rect 47192 50564 47196 50620
rect 47196 50564 47252 50620
rect 47252 50564 47256 50620
rect 47192 50560 47256 50564
rect 51952 50620 52016 50624
rect 51952 50564 51956 50620
rect 51956 50564 52012 50620
rect 52012 50564 52016 50620
rect 51952 50560 52016 50564
rect 52032 50620 52096 50624
rect 52032 50564 52036 50620
rect 52036 50564 52092 50620
rect 52092 50564 52096 50620
rect 52032 50560 52096 50564
rect 52112 50620 52176 50624
rect 52112 50564 52116 50620
rect 52116 50564 52172 50620
rect 52172 50564 52176 50620
rect 52112 50560 52176 50564
rect 52192 50620 52256 50624
rect 52192 50564 52196 50620
rect 52196 50564 52252 50620
rect 52252 50564 52256 50620
rect 52192 50560 52256 50564
rect 56952 50620 57016 50624
rect 56952 50564 56956 50620
rect 56956 50564 57012 50620
rect 57012 50564 57016 50620
rect 56952 50560 57016 50564
rect 57032 50620 57096 50624
rect 57032 50564 57036 50620
rect 57036 50564 57092 50620
rect 57092 50564 57096 50620
rect 57032 50560 57096 50564
rect 57112 50620 57176 50624
rect 57112 50564 57116 50620
rect 57116 50564 57172 50620
rect 57172 50564 57176 50620
rect 57112 50560 57176 50564
rect 57192 50620 57256 50624
rect 57192 50564 57196 50620
rect 57196 50564 57252 50620
rect 57252 50564 57256 50620
rect 57192 50560 57256 50564
rect 2612 50076 2676 50080
rect 2612 50020 2616 50076
rect 2616 50020 2672 50076
rect 2672 50020 2676 50076
rect 2612 50016 2676 50020
rect 2692 50076 2756 50080
rect 2692 50020 2696 50076
rect 2696 50020 2752 50076
rect 2752 50020 2756 50076
rect 2692 50016 2756 50020
rect 2772 50076 2836 50080
rect 2772 50020 2776 50076
rect 2776 50020 2832 50076
rect 2832 50020 2836 50076
rect 2772 50016 2836 50020
rect 2852 50076 2916 50080
rect 2852 50020 2856 50076
rect 2856 50020 2912 50076
rect 2912 50020 2916 50076
rect 2852 50016 2916 50020
rect 7612 50076 7676 50080
rect 7612 50020 7616 50076
rect 7616 50020 7672 50076
rect 7672 50020 7676 50076
rect 7612 50016 7676 50020
rect 7692 50076 7756 50080
rect 7692 50020 7696 50076
rect 7696 50020 7752 50076
rect 7752 50020 7756 50076
rect 7692 50016 7756 50020
rect 7772 50076 7836 50080
rect 7772 50020 7776 50076
rect 7776 50020 7832 50076
rect 7832 50020 7836 50076
rect 7772 50016 7836 50020
rect 7852 50076 7916 50080
rect 7852 50020 7856 50076
rect 7856 50020 7912 50076
rect 7912 50020 7916 50076
rect 7852 50016 7916 50020
rect 12612 50076 12676 50080
rect 12612 50020 12616 50076
rect 12616 50020 12672 50076
rect 12672 50020 12676 50076
rect 12612 50016 12676 50020
rect 12692 50076 12756 50080
rect 12692 50020 12696 50076
rect 12696 50020 12752 50076
rect 12752 50020 12756 50076
rect 12692 50016 12756 50020
rect 12772 50076 12836 50080
rect 12772 50020 12776 50076
rect 12776 50020 12832 50076
rect 12832 50020 12836 50076
rect 12772 50016 12836 50020
rect 12852 50076 12916 50080
rect 12852 50020 12856 50076
rect 12856 50020 12912 50076
rect 12912 50020 12916 50076
rect 12852 50016 12916 50020
rect 17612 50076 17676 50080
rect 17612 50020 17616 50076
rect 17616 50020 17672 50076
rect 17672 50020 17676 50076
rect 17612 50016 17676 50020
rect 17692 50076 17756 50080
rect 17692 50020 17696 50076
rect 17696 50020 17752 50076
rect 17752 50020 17756 50076
rect 17692 50016 17756 50020
rect 17772 50076 17836 50080
rect 17772 50020 17776 50076
rect 17776 50020 17832 50076
rect 17832 50020 17836 50076
rect 17772 50016 17836 50020
rect 17852 50076 17916 50080
rect 17852 50020 17856 50076
rect 17856 50020 17912 50076
rect 17912 50020 17916 50076
rect 17852 50016 17916 50020
rect 22612 50076 22676 50080
rect 22612 50020 22616 50076
rect 22616 50020 22672 50076
rect 22672 50020 22676 50076
rect 22612 50016 22676 50020
rect 22692 50076 22756 50080
rect 22692 50020 22696 50076
rect 22696 50020 22752 50076
rect 22752 50020 22756 50076
rect 22692 50016 22756 50020
rect 22772 50076 22836 50080
rect 22772 50020 22776 50076
rect 22776 50020 22832 50076
rect 22832 50020 22836 50076
rect 22772 50016 22836 50020
rect 22852 50076 22916 50080
rect 22852 50020 22856 50076
rect 22856 50020 22912 50076
rect 22912 50020 22916 50076
rect 22852 50016 22916 50020
rect 27612 50076 27676 50080
rect 27612 50020 27616 50076
rect 27616 50020 27672 50076
rect 27672 50020 27676 50076
rect 27612 50016 27676 50020
rect 27692 50076 27756 50080
rect 27692 50020 27696 50076
rect 27696 50020 27752 50076
rect 27752 50020 27756 50076
rect 27692 50016 27756 50020
rect 27772 50076 27836 50080
rect 27772 50020 27776 50076
rect 27776 50020 27832 50076
rect 27832 50020 27836 50076
rect 27772 50016 27836 50020
rect 27852 50076 27916 50080
rect 27852 50020 27856 50076
rect 27856 50020 27912 50076
rect 27912 50020 27916 50076
rect 27852 50016 27916 50020
rect 32612 50076 32676 50080
rect 32612 50020 32616 50076
rect 32616 50020 32672 50076
rect 32672 50020 32676 50076
rect 32612 50016 32676 50020
rect 32692 50076 32756 50080
rect 32692 50020 32696 50076
rect 32696 50020 32752 50076
rect 32752 50020 32756 50076
rect 32692 50016 32756 50020
rect 32772 50076 32836 50080
rect 32772 50020 32776 50076
rect 32776 50020 32832 50076
rect 32832 50020 32836 50076
rect 32772 50016 32836 50020
rect 32852 50076 32916 50080
rect 32852 50020 32856 50076
rect 32856 50020 32912 50076
rect 32912 50020 32916 50076
rect 32852 50016 32916 50020
rect 37612 50076 37676 50080
rect 37612 50020 37616 50076
rect 37616 50020 37672 50076
rect 37672 50020 37676 50076
rect 37612 50016 37676 50020
rect 37692 50076 37756 50080
rect 37692 50020 37696 50076
rect 37696 50020 37752 50076
rect 37752 50020 37756 50076
rect 37692 50016 37756 50020
rect 37772 50076 37836 50080
rect 37772 50020 37776 50076
rect 37776 50020 37832 50076
rect 37832 50020 37836 50076
rect 37772 50016 37836 50020
rect 37852 50076 37916 50080
rect 37852 50020 37856 50076
rect 37856 50020 37912 50076
rect 37912 50020 37916 50076
rect 37852 50016 37916 50020
rect 42612 50076 42676 50080
rect 42612 50020 42616 50076
rect 42616 50020 42672 50076
rect 42672 50020 42676 50076
rect 42612 50016 42676 50020
rect 42692 50076 42756 50080
rect 42692 50020 42696 50076
rect 42696 50020 42752 50076
rect 42752 50020 42756 50076
rect 42692 50016 42756 50020
rect 42772 50076 42836 50080
rect 42772 50020 42776 50076
rect 42776 50020 42832 50076
rect 42832 50020 42836 50076
rect 42772 50016 42836 50020
rect 42852 50076 42916 50080
rect 42852 50020 42856 50076
rect 42856 50020 42912 50076
rect 42912 50020 42916 50076
rect 42852 50016 42916 50020
rect 47612 50076 47676 50080
rect 47612 50020 47616 50076
rect 47616 50020 47672 50076
rect 47672 50020 47676 50076
rect 47612 50016 47676 50020
rect 47692 50076 47756 50080
rect 47692 50020 47696 50076
rect 47696 50020 47752 50076
rect 47752 50020 47756 50076
rect 47692 50016 47756 50020
rect 47772 50076 47836 50080
rect 47772 50020 47776 50076
rect 47776 50020 47832 50076
rect 47832 50020 47836 50076
rect 47772 50016 47836 50020
rect 47852 50076 47916 50080
rect 47852 50020 47856 50076
rect 47856 50020 47912 50076
rect 47912 50020 47916 50076
rect 47852 50016 47916 50020
rect 52612 50076 52676 50080
rect 52612 50020 52616 50076
rect 52616 50020 52672 50076
rect 52672 50020 52676 50076
rect 52612 50016 52676 50020
rect 52692 50076 52756 50080
rect 52692 50020 52696 50076
rect 52696 50020 52752 50076
rect 52752 50020 52756 50076
rect 52692 50016 52756 50020
rect 52772 50076 52836 50080
rect 52772 50020 52776 50076
rect 52776 50020 52832 50076
rect 52832 50020 52836 50076
rect 52772 50016 52836 50020
rect 52852 50076 52916 50080
rect 52852 50020 52856 50076
rect 52856 50020 52912 50076
rect 52912 50020 52916 50076
rect 52852 50016 52916 50020
rect 57612 50076 57676 50080
rect 57612 50020 57616 50076
rect 57616 50020 57672 50076
rect 57672 50020 57676 50076
rect 57612 50016 57676 50020
rect 57692 50076 57756 50080
rect 57692 50020 57696 50076
rect 57696 50020 57752 50076
rect 57752 50020 57756 50076
rect 57692 50016 57756 50020
rect 57772 50076 57836 50080
rect 57772 50020 57776 50076
rect 57776 50020 57832 50076
rect 57832 50020 57836 50076
rect 57772 50016 57836 50020
rect 57852 50076 57916 50080
rect 57852 50020 57856 50076
rect 57856 50020 57912 50076
rect 57912 50020 57916 50076
rect 57852 50016 57916 50020
rect 1952 49532 2016 49536
rect 1952 49476 1956 49532
rect 1956 49476 2012 49532
rect 2012 49476 2016 49532
rect 1952 49472 2016 49476
rect 2032 49532 2096 49536
rect 2032 49476 2036 49532
rect 2036 49476 2092 49532
rect 2092 49476 2096 49532
rect 2032 49472 2096 49476
rect 2112 49532 2176 49536
rect 2112 49476 2116 49532
rect 2116 49476 2172 49532
rect 2172 49476 2176 49532
rect 2112 49472 2176 49476
rect 2192 49532 2256 49536
rect 2192 49476 2196 49532
rect 2196 49476 2252 49532
rect 2252 49476 2256 49532
rect 2192 49472 2256 49476
rect 6952 49532 7016 49536
rect 6952 49476 6956 49532
rect 6956 49476 7012 49532
rect 7012 49476 7016 49532
rect 6952 49472 7016 49476
rect 7032 49532 7096 49536
rect 7032 49476 7036 49532
rect 7036 49476 7092 49532
rect 7092 49476 7096 49532
rect 7032 49472 7096 49476
rect 7112 49532 7176 49536
rect 7112 49476 7116 49532
rect 7116 49476 7172 49532
rect 7172 49476 7176 49532
rect 7112 49472 7176 49476
rect 7192 49532 7256 49536
rect 7192 49476 7196 49532
rect 7196 49476 7252 49532
rect 7252 49476 7256 49532
rect 7192 49472 7256 49476
rect 11952 49532 12016 49536
rect 11952 49476 11956 49532
rect 11956 49476 12012 49532
rect 12012 49476 12016 49532
rect 11952 49472 12016 49476
rect 12032 49532 12096 49536
rect 12032 49476 12036 49532
rect 12036 49476 12092 49532
rect 12092 49476 12096 49532
rect 12032 49472 12096 49476
rect 12112 49532 12176 49536
rect 12112 49476 12116 49532
rect 12116 49476 12172 49532
rect 12172 49476 12176 49532
rect 12112 49472 12176 49476
rect 12192 49532 12256 49536
rect 12192 49476 12196 49532
rect 12196 49476 12252 49532
rect 12252 49476 12256 49532
rect 12192 49472 12256 49476
rect 16952 49532 17016 49536
rect 16952 49476 16956 49532
rect 16956 49476 17012 49532
rect 17012 49476 17016 49532
rect 16952 49472 17016 49476
rect 17032 49532 17096 49536
rect 17032 49476 17036 49532
rect 17036 49476 17092 49532
rect 17092 49476 17096 49532
rect 17032 49472 17096 49476
rect 17112 49532 17176 49536
rect 17112 49476 17116 49532
rect 17116 49476 17172 49532
rect 17172 49476 17176 49532
rect 17112 49472 17176 49476
rect 17192 49532 17256 49536
rect 17192 49476 17196 49532
rect 17196 49476 17252 49532
rect 17252 49476 17256 49532
rect 17192 49472 17256 49476
rect 21952 49532 22016 49536
rect 21952 49476 21956 49532
rect 21956 49476 22012 49532
rect 22012 49476 22016 49532
rect 21952 49472 22016 49476
rect 22032 49532 22096 49536
rect 22032 49476 22036 49532
rect 22036 49476 22092 49532
rect 22092 49476 22096 49532
rect 22032 49472 22096 49476
rect 22112 49532 22176 49536
rect 22112 49476 22116 49532
rect 22116 49476 22172 49532
rect 22172 49476 22176 49532
rect 22112 49472 22176 49476
rect 22192 49532 22256 49536
rect 22192 49476 22196 49532
rect 22196 49476 22252 49532
rect 22252 49476 22256 49532
rect 22192 49472 22256 49476
rect 26952 49532 27016 49536
rect 26952 49476 26956 49532
rect 26956 49476 27012 49532
rect 27012 49476 27016 49532
rect 26952 49472 27016 49476
rect 27032 49532 27096 49536
rect 27032 49476 27036 49532
rect 27036 49476 27092 49532
rect 27092 49476 27096 49532
rect 27032 49472 27096 49476
rect 27112 49532 27176 49536
rect 27112 49476 27116 49532
rect 27116 49476 27172 49532
rect 27172 49476 27176 49532
rect 27112 49472 27176 49476
rect 27192 49532 27256 49536
rect 27192 49476 27196 49532
rect 27196 49476 27252 49532
rect 27252 49476 27256 49532
rect 27192 49472 27256 49476
rect 31952 49532 32016 49536
rect 31952 49476 31956 49532
rect 31956 49476 32012 49532
rect 32012 49476 32016 49532
rect 31952 49472 32016 49476
rect 32032 49532 32096 49536
rect 32032 49476 32036 49532
rect 32036 49476 32092 49532
rect 32092 49476 32096 49532
rect 32032 49472 32096 49476
rect 32112 49532 32176 49536
rect 32112 49476 32116 49532
rect 32116 49476 32172 49532
rect 32172 49476 32176 49532
rect 32112 49472 32176 49476
rect 32192 49532 32256 49536
rect 32192 49476 32196 49532
rect 32196 49476 32252 49532
rect 32252 49476 32256 49532
rect 32192 49472 32256 49476
rect 36952 49532 37016 49536
rect 36952 49476 36956 49532
rect 36956 49476 37012 49532
rect 37012 49476 37016 49532
rect 36952 49472 37016 49476
rect 37032 49532 37096 49536
rect 37032 49476 37036 49532
rect 37036 49476 37092 49532
rect 37092 49476 37096 49532
rect 37032 49472 37096 49476
rect 37112 49532 37176 49536
rect 37112 49476 37116 49532
rect 37116 49476 37172 49532
rect 37172 49476 37176 49532
rect 37112 49472 37176 49476
rect 37192 49532 37256 49536
rect 37192 49476 37196 49532
rect 37196 49476 37252 49532
rect 37252 49476 37256 49532
rect 37192 49472 37256 49476
rect 41952 49532 42016 49536
rect 41952 49476 41956 49532
rect 41956 49476 42012 49532
rect 42012 49476 42016 49532
rect 41952 49472 42016 49476
rect 42032 49532 42096 49536
rect 42032 49476 42036 49532
rect 42036 49476 42092 49532
rect 42092 49476 42096 49532
rect 42032 49472 42096 49476
rect 42112 49532 42176 49536
rect 42112 49476 42116 49532
rect 42116 49476 42172 49532
rect 42172 49476 42176 49532
rect 42112 49472 42176 49476
rect 42192 49532 42256 49536
rect 42192 49476 42196 49532
rect 42196 49476 42252 49532
rect 42252 49476 42256 49532
rect 42192 49472 42256 49476
rect 46952 49532 47016 49536
rect 46952 49476 46956 49532
rect 46956 49476 47012 49532
rect 47012 49476 47016 49532
rect 46952 49472 47016 49476
rect 47032 49532 47096 49536
rect 47032 49476 47036 49532
rect 47036 49476 47092 49532
rect 47092 49476 47096 49532
rect 47032 49472 47096 49476
rect 47112 49532 47176 49536
rect 47112 49476 47116 49532
rect 47116 49476 47172 49532
rect 47172 49476 47176 49532
rect 47112 49472 47176 49476
rect 47192 49532 47256 49536
rect 47192 49476 47196 49532
rect 47196 49476 47252 49532
rect 47252 49476 47256 49532
rect 47192 49472 47256 49476
rect 51952 49532 52016 49536
rect 51952 49476 51956 49532
rect 51956 49476 52012 49532
rect 52012 49476 52016 49532
rect 51952 49472 52016 49476
rect 52032 49532 52096 49536
rect 52032 49476 52036 49532
rect 52036 49476 52092 49532
rect 52092 49476 52096 49532
rect 52032 49472 52096 49476
rect 52112 49532 52176 49536
rect 52112 49476 52116 49532
rect 52116 49476 52172 49532
rect 52172 49476 52176 49532
rect 52112 49472 52176 49476
rect 52192 49532 52256 49536
rect 52192 49476 52196 49532
rect 52196 49476 52252 49532
rect 52252 49476 52256 49532
rect 52192 49472 52256 49476
rect 56952 49532 57016 49536
rect 56952 49476 56956 49532
rect 56956 49476 57012 49532
rect 57012 49476 57016 49532
rect 56952 49472 57016 49476
rect 57032 49532 57096 49536
rect 57032 49476 57036 49532
rect 57036 49476 57092 49532
rect 57092 49476 57096 49532
rect 57032 49472 57096 49476
rect 57112 49532 57176 49536
rect 57112 49476 57116 49532
rect 57116 49476 57172 49532
rect 57172 49476 57176 49532
rect 57112 49472 57176 49476
rect 57192 49532 57256 49536
rect 57192 49476 57196 49532
rect 57196 49476 57252 49532
rect 57252 49476 57256 49532
rect 57192 49472 57256 49476
rect 2612 48988 2676 48992
rect 2612 48932 2616 48988
rect 2616 48932 2672 48988
rect 2672 48932 2676 48988
rect 2612 48928 2676 48932
rect 2692 48988 2756 48992
rect 2692 48932 2696 48988
rect 2696 48932 2752 48988
rect 2752 48932 2756 48988
rect 2692 48928 2756 48932
rect 2772 48988 2836 48992
rect 2772 48932 2776 48988
rect 2776 48932 2832 48988
rect 2832 48932 2836 48988
rect 2772 48928 2836 48932
rect 2852 48988 2916 48992
rect 2852 48932 2856 48988
rect 2856 48932 2912 48988
rect 2912 48932 2916 48988
rect 2852 48928 2916 48932
rect 7612 48988 7676 48992
rect 7612 48932 7616 48988
rect 7616 48932 7672 48988
rect 7672 48932 7676 48988
rect 7612 48928 7676 48932
rect 7692 48988 7756 48992
rect 7692 48932 7696 48988
rect 7696 48932 7752 48988
rect 7752 48932 7756 48988
rect 7692 48928 7756 48932
rect 7772 48988 7836 48992
rect 7772 48932 7776 48988
rect 7776 48932 7832 48988
rect 7832 48932 7836 48988
rect 7772 48928 7836 48932
rect 7852 48988 7916 48992
rect 7852 48932 7856 48988
rect 7856 48932 7912 48988
rect 7912 48932 7916 48988
rect 7852 48928 7916 48932
rect 12612 48988 12676 48992
rect 12612 48932 12616 48988
rect 12616 48932 12672 48988
rect 12672 48932 12676 48988
rect 12612 48928 12676 48932
rect 12692 48988 12756 48992
rect 12692 48932 12696 48988
rect 12696 48932 12752 48988
rect 12752 48932 12756 48988
rect 12692 48928 12756 48932
rect 12772 48988 12836 48992
rect 12772 48932 12776 48988
rect 12776 48932 12832 48988
rect 12832 48932 12836 48988
rect 12772 48928 12836 48932
rect 12852 48988 12916 48992
rect 12852 48932 12856 48988
rect 12856 48932 12912 48988
rect 12912 48932 12916 48988
rect 12852 48928 12916 48932
rect 17612 48988 17676 48992
rect 17612 48932 17616 48988
rect 17616 48932 17672 48988
rect 17672 48932 17676 48988
rect 17612 48928 17676 48932
rect 17692 48988 17756 48992
rect 17692 48932 17696 48988
rect 17696 48932 17752 48988
rect 17752 48932 17756 48988
rect 17692 48928 17756 48932
rect 17772 48988 17836 48992
rect 17772 48932 17776 48988
rect 17776 48932 17832 48988
rect 17832 48932 17836 48988
rect 17772 48928 17836 48932
rect 17852 48988 17916 48992
rect 17852 48932 17856 48988
rect 17856 48932 17912 48988
rect 17912 48932 17916 48988
rect 17852 48928 17916 48932
rect 22612 48988 22676 48992
rect 22612 48932 22616 48988
rect 22616 48932 22672 48988
rect 22672 48932 22676 48988
rect 22612 48928 22676 48932
rect 22692 48988 22756 48992
rect 22692 48932 22696 48988
rect 22696 48932 22752 48988
rect 22752 48932 22756 48988
rect 22692 48928 22756 48932
rect 22772 48988 22836 48992
rect 22772 48932 22776 48988
rect 22776 48932 22832 48988
rect 22832 48932 22836 48988
rect 22772 48928 22836 48932
rect 22852 48988 22916 48992
rect 22852 48932 22856 48988
rect 22856 48932 22912 48988
rect 22912 48932 22916 48988
rect 22852 48928 22916 48932
rect 27612 48988 27676 48992
rect 27612 48932 27616 48988
rect 27616 48932 27672 48988
rect 27672 48932 27676 48988
rect 27612 48928 27676 48932
rect 27692 48988 27756 48992
rect 27692 48932 27696 48988
rect 27696 48932 27752 48988
rect 27752 48932 27756 48988
rect 27692 48928 27756 48932
rect 27772 48988 27836 48992
rect 27772 48932 27776 48988
rect 27776 48932 27832 48988
rect 27832 48932 27836 48988
rect 27772 48928 27836 48932
rect 27852 48988 27916 48992
rect 27852 48932 27856 48988
rect 27856 48932 27912 48988
rect 27912 48932 27916 48988
rect 27852 48928 27916 48932
rect 32612 48988 32676 48992
rect 32612 48932 32616 48988
rect 32616 48932 32672 48988
rect 32672 48932 32676 48988
rect 32612 48928 32676 48932
rect 32692 48988 32756 48992
rect 32692 48932 32696 48988
rect 32696 48932 32752 48988
rect 32752 48932 32756 48988
rect 32692 48928 32756 48932
rect 32772 48988 32836 48992
rect 32772 48932 32776 48988
rect 32776 48932 32832 48988
rect 32832 48932 32836 48988
rect 32772 48928 32836 48932
rect 32852 48988 32916 48992
rect 32852 48932 32856 48988
rect 32856 48932 32912 48988
rect 32912 48932 32916 48988
rect 32852 48928 32916 48932
rect 37612 48988 37676 48992
rect 37612 48932 37616 48988
rect 37616 48932 37672 48988
rect 37672 48932 37676 48988
rect 37612 48928 37676 48932
rect 37692 48988 37756 48992
rect 37692 48932 37696 48988
rect 37696 48932 37752 48988
rect 37752 48932 37756 48988
rect 37692 48928 37756 48932
rect 37772 48988 37836 48992
rect 37772 48932 37776 48988
rect 37776 48932 37832 48988
rect 37832 48932 37836 48988
rect 37772 48928 37836 48932
rect 37852 48988 37916 48992
rect 37852 48932 37856 48988
rect 37856 48932 37912 48988
rect 37912 48932 37916 48988
rect 37852 48928 37916 48932
rect 42612 48988 42676 48992
rect 42612 48932 42616 48988
rect 42616 48932 42672 48988
rect 42672 48932 42676 48988
rect 42612 48928 42676 48932
rect 42692 48988 42756 48992
rect 42692 48932 42696 48988
rect 42696 48932 42752 48988
rect 42752 48932 42756 48988
rect 42692 48928 42756 48932
rect 42772 48988 42836 48992
rect 42772 48932 42776 48988
rect 42776 48932 42832 48988
rect 42832 48932 42836 48988
rect 42772 48928 42836 48932
rect 42852 48988 42916 48992
rect 42852 48932 42856 48988
rect 42856 48932 42912 48988
rect 42912 48932 42916 48988
rect 42852 48928 42916 48932
rect 47612 48988 47676 48992
rect 47612 48932 47616 48988
rect 47616 48932 47672 48988
rect 47672 48932 47676 48988
rect 47612 48928 47676 48932
rect 47692 48988 47756 48992
rect 47692 48932 47696 48988
rect 47696 48932 47752 48988
rect 47752 48932 47756 48988
rect 47692 48928 47756 48932
rect 47772 48988 47836 48992
rect 47772 48932 47776 48988
rect 47776 48932 47832 48988
rect 47832 48932 47836 48988
rect 47772 48928 47836 48932
rect 47852 48988 47916 48992
rect 47852 48932 47856 48988
rect 47856 48932 47912 48988
rect 47912 48932 47916 48988
rect 47852 48928 47916 48932
rect 52612 48988 52676 48992
rect 52612 48932 52616 48988
rect 52616 48932 52672 48988
rect 52672 48932 52676 48988
rect 52612 48928 52676 48932
rect 52692 48988 52756 48992
rect 52692 48932 52696 48988
rect 52696 48932 52752 48988
rect 52752 48932 52756 48988
rect 52692 48928 52756 48932
rect 52772 48988 52836 48992
rect 52772 48932 52776 48988
rect 52776 48932 52832 48988
rect 52832 48932 52836 48988
rect 52772 48928 52836 48932
rect 52852 48988 52916 48992
rect 52852 48932 52856 48988
rect 52856 48932 52912 48988
rect 52912 48932 52916 48988
rect 52852 48928 52916 48932
rect 57612 48988 57676 48992
rect 57612 48932 57616 48988
rect 57616 48932 57672 48988
rect 57672 48932 57676 48988
rect 57612 48928 57676 48932
rect 57692 48988 57756 48992
rect 57692 48932 57696 48988
rect 57696 48932 57752 48988
rect 57752 48932 57756 48988
rect 57692 48928 57756 48932
rect 57772 48988 57836 48992
rect 57772 48932 57776 48988
rect 57776 48932 57832 48988
rect 57832 48932 57836 48988
rect 57772 48928 57836 48932
rect 57852 48988 57916 48992
rect 57852 48932 57856 48988
rect 57856 48932 57912 48988
rect 57912 48932 57916 48988
rect 57852 48928 57916 48932
rect 1952 48444 2016 48448
rect 1952 48388 1956 48444
rect 1956 48388 2012 48444
rect 2012 48388 2016 48444
rect 1952 48384 2016 48388
rect 2032 48444 2096 48448
rect 2032 48388 2036 48444
rect 2036 48388 2092 48444
rect 2092 48388 2096 48444
rect 2032 48384 2096 48388
rect 2112 48444 2176 48448
rect 2112 48388 2116 48444
rect 2116 48388 2172 48444
rect 2172 48388 2176 48444
rect 2112 48384 2176 48388
rect 2192 48444 2256 48448
rect 2192 48388 2196 48444
rect 2196 48388 2252 48444
rect 2252 48388 2256 48444
rect 2192 48384 2256 48388
rect 6952 48444 7016 48448
rect 6952 48388 6956 48444
rect 6956 48388 7012 48444
rect 7012 48388 7016 48444
rect 6952 48384 7016 48388
rect 7032 48444 7096 48448
rect 7032 48388 7036 48444
rect 7036 48388 7092 48444
rect 7092 48388 7096 48444
rect 7032 48384 7096 48388
rect 7112 48444 7176 48448
rect 7112 48388 7116 48444
rect 7116 48388 7172 48444
rect 7172 48388 7176 48444
rect 7112 48384 7176 48388
rect 7192 48444 7256 48448
rect 7192 48388 7196 48444
rect 7196 48388 7252 48444
rect 7252 48388 7256 48444
rect 7192 48384 7256 48388
rect 11952 48444 12016 48448
rect 11952 48388 11956 48444
rect 11956 48388 12012 48444
rect 12012 48388 12016 48444
rect 11952 48384 12016 48388
rect 12032 48444 12096 48448
rect 12032 48388 12036 48444
rect 12036 48388 12092 48444
rect 12092 48388 12096 48444
rect 12032 48384 12096 48388
rect 12112 48444 12176 48448
rect 12112 48388 12116 48444
rect 12116 48388 12172 48444
rect 12172 48388 12176 48444
rect 12112 48384 12176 48388
rect 12192 48444 12256 48448
rect 12192 48388 12196 48444
rect 12196 48388 12252 48444
rect 12252 48388 12256 48444
rect 12192 48384 12256 48388
rect 16952 48444 17016 48448
rect 16952 48388 16956 48444
rect 16956 48388 17012 48444
rect 17012 48388 17016 48444
rect 16952 48384 17016 48388
rect 17032 48444 17096 48448
rect 17032 48388 17036 48444
rect 17036 48388 17092 48444
rect 17092 48388 17096 48444
rect 17032 48384 17096 48388
rect 17112 48444 17176 48448
rect 17112 48388 17116 48444
rect 17116 48388 17172 48444
rect 17172 48388 17176 48444
rect 17112 48384 17176 48388
rect 17192 48444 17256 48448
rect 17192 48388 17196 48444
rect 17196 48388 17252 48444
rect 17252 48388 17256 48444
rect 17192 48384 17256 48388
rect 21952 48444 22016 48448
rect 21952 48388 21956 48444
rect 21956 48388 22012 48444
rect 22012 48388 22016 48444
rect 21952 48384 22016 48388
rect 22032 48444 22096 48448
rect 22032 48388 22036 48444
rect 22036 48388 22092 48444
rect 22092 48388 22096 48444
rect 22032 48384 22096 48388
rect 22112 48444 22176 48448
rect 22112 48388 22116 48444
rect 22116 48388 22172 48444
rect 22172 48388 22176 48444
rect 22112 48384 22176 48388
rect 22192 48444 22256 48448
rect 22192 48388 22196 48444
rect 22196 48388 22252 48444
rect 22252 48388 22256 48444
rect 22192 48384 22256 48388
rect 26952 48444 27016 48448
rect 26952 48388 26956 48444
rect 26956 48388 27012 48444
rect 27012 48388 27016 48444
rect 26952 48384 27016 48388
rect 27032 48444 27096 48448
rect 27032 48388 27036 48444
rect 27036 48388 27092 48444
rect 27092 48388 27096 48444
rect 27032 48384 27096 48388
rect 27112 48444 27176 48448
rect 27112 48388 27116 48444
rect 27116 48388 27172 48444
rect 27172 48388 27176 48444
rect 27112 48384 27176 48388
rect 27192 48444 27256 48448
rect 27192 48388 27196 48444
rect 27196 48388 27252 48444
rect 27252 48388 27256 48444
rect 27192 48384 27256 48388
rect 31952 48444 32016 48448
rect 31952 48388 31956 48444
rect 31956 48388 32012 48444
rect 32012 48388 32016 48444
rect 31952 48384 32016 48388
rect 32032 48444 32096 48448
rect 32032 48388 32036 48444
rect 32036 48388 32092 48444
rect 32092 48388 32096 48444
rect 32032 48384 32096 48388
rect 32112 48444 32176 48448
rect 32112 48388 32116 48444
rect 32116 48388 32172 48444
rect 32172 48388 32176 48444
rect 32112 48384 32176 48388
rect 32192 48444 32256 48448
rect 32192 48388 32196 48444
rect 32196 48388 32252 48444
rect 32252 48388 32256 48444
rect 32192 48384 32256 48388
rect 36952 48444 37016 48448
rect 36952 48388 36956 48444
rect 36956 48388 37012 48444
rect 37012 48388 37016 48444
rect 36952 48384 37016 48388
rect 37032 48444 37096 48448
rect 37032 48388 37036 48444
rect 37036 48388 37092 48444
rect 37092 48388 37096 48444
rect 37032 48384 37096 48388
rect 37112 48444 37176 48448
rect 37112 48388 37116 48444
rect 37116 48388 37172 48444
rect 37172 48388 37176 48444
rect 37112 48384 37176 48388
rect 37192 48444 37256 48448
rect 37192 48388 37196 48444
rect 37196 48388 37252 48444
rect 37252 48388 37256 48444
rect 37192 48384 37256 48388
rect 41952 48444 42016 48448
rect 41952 48388 41956 48444
rect 41956 48388 42012 48444
rect 42012 48388 42016 48444
rect 41952 48384 42016 48388
rect 42032 48444 42096 48448
rect 42032 48388 42036 48444
rect 42036 48388 42092 48444
rect 42092 48388 42096 48444
rect 42032 48384 42096 48388
rect 42112 48444 42176 48448
rect 42112 48388 42116 48444
rect 42116 48388 42172 48444
rect 42172 48388 42176 48444
rect 42112 48384 42176 48388
rect 42192 48444 42256 48448
rect 42192 48388 42196 48444
rect 42196 48388 42252 48444
rect 42252 48388 42256 48444
rect 42192 48384 42256 48388
rect 46952 48444 47016 48448
rect 46952 48388 46956 48444
rect 46956 48388 47012 48444
rect 47012 48388 47016 48444
rect 46952 48384 47016 48388
rect 47032 48444 47096 48448
rect 47032 48388 47036 48444
rect 47036 48388 47092 48444
rect 47092 48388 47096 48444
rect 47032 48384 47096 48388
rect 47112 48444 47176 48448
rect 47112 48388 47116 48444
rect 47116 48388 47172 48444
rect 47172 48388 47176 48444
rect 47112 48384 47176 48388
rect 47192 48444 47256 48448
rect 47192 48388 47196 48444
rect 47196 48388 47252 48444
rect 47252 48388 47256 48444
rect 47192 48384 47256 48388
rect 51952 48444 52016 48448
rect 51952 48388 51956 48444
rect 51956 48388 52012 48444
rect 52012 48388 52016 48444
rect 51952 48384 52016 48388
rect 52032 48444 52096 48448
rect 52032 48388 52036 48444
rect 52036 48388 52092 48444
rect 52092 48388 52096 48444
rect 52032 48384 52096 48388
rect 52112 48444 52176 48448
rect 52112 48388 52116 48444
rect 52116 48388 52172 48444
rect 52172 48388 52176 48444
rect 52112 48384 52176 48388
rect 52192 48444 52256 48448
rect 52192 48388 52196 48444
rect 52196 48388 52252 48444
rect 52252 48388 52256 48444
rect 52192 48384 52256 48388
rect 56952 48444 57016 48448
rect 56952 48388 56956 48444
rect 56956 48388 57012 48444
rect 57012 48388 57016 48444
rect 56952 48384 57016 48388
rect 57032 48444 57096 48448
rect 57032 48388 57036 48444
rect 57036 48388 57092 48444
rect 57092 48388 57096 48444
rect 57032 48384 57096 48388
rect 57112 48444 57176 48448
rect 57112 48388 57116 48444
rect 57116 48388 57172 48444
rect 57172 48388 57176 48444
rect 57112 48384 57176 48388
rect 57192 48444 57256 48448
rect 57192 48388 57196 48444
rect 57196 48388 57252 48444
rect 57252 48388 57256 48444
rect 57192 48384 57256 48388
rect 2612 47900 2676 47904
rect 2612 47844 2616 47900
rect 2616 47844 2672 47900
rect 2672 47844 2676 47900
rect 2612 47840 2676 47844
rect 2692 47900 2756 47904
rect 2692 47844 2696 47900
rect 2696 47844 2752 47900
rect 2752 47844 2756 47900
rect 2692 47840 2756 47844
rect 2772 47900 2836 47904
rect 2772 47844 2776 47900
rect 2776 47844 2832 47900
rect 2832 47844 2836 47900
rect 2772 47840 2836 47844
rect 2852 47900 2916 47904
rect 2852 47844 2856 47900
rect 2856 47844 2912 47900
rect 2912 47844 2916 47900
rect 2852 47840 2916 47844
rect 7612 47900 7676 47904
rect 7612 47844 7616 47900
rect 7616 47844 7672 47900
rect 7672 47844 7676 47900
rect 7612 47840 7676 47844
rect 7692 47900 7756 47904
rect 7692 47844 7696 47900
rect 7696 47844 7752 47900
rect 7752 47844 7756 47900
rect 7692 47840 7756 47844
rect 7772 47900 7836 47904
rect 7772 47844 7776 47900
rect 7776 47844 7832 47900
rect 7832 47844 7836 47900
rect 7772 47840 7836 47844
rect 7852 47900 7916 47904
rect 7852 47844 7856 47900
rect 7856 47844 7912 47900
rect 7912 47844 7916 47900
rect 7852 47840 7916 47844
rect 12612 47900 12676 47904
rect 12612 47844 12616 47900
rect 12616 47844 12672 47900
rect 12672 47844 12676 47900
rect 12612 47840 12676 47844
rect 12692 47900 12756 47904
rect 12692 47844 12696 47900
rect 12696 47844 12752 47900
rect 12752 47844 12756 47900
rect 12692 47840 12756 47844
rect 12772 47900 12836 47904
rect 12772 47844 12776 47900
rect 12776 47844 12832 47900
rect 12832 47844 12836 47900
rect 12772 47840 12836 47844
rect 12852 47900 12916 47904
rect 12852 47844 12856 47900
rect 12856 47844 12912 47900
rect 12912 47844 12916 47900
rect 12852 47840 12916 47844
rect 17612 47900 17676 47904
rect 17612 47844 17616 47900
rect 17616 47844 17672 47900
rect 17672 47844 17676 47900
rect 17612 47840 17676 47844
rect 17692 47900 17756 47904
rect 17692 47844 17696 47900
rect 17696 47844 17752 47900
rect 17752 47844 17756 47900
rect 17692 47840 17756 47844
rect 17772 47900 17836 47904
rect 17772 47844 17776 47900
rect 17776 47844 17832 47900
rect 17832 47844 17836 47900
rect 17772 47840 17836 47844
rect 17852 47900 17916 47904
rect 17852 47844 17856 47900
rect 17856 47844 17912 47900
rect 17912 47844 17916 47900
rect 17852 47840 17916 47844
rect 22612 47900 22676 47904
rect 22612 47844 22616 47900
rect 22616 47844 22672 47900
rect 22672 47844 22676 47900
rect 22612 47840 22676 47844
rect 22692 47900 22756 47904
rect 22692 47844 22696 47900
rect 22696 47844 22752 47900
rect 22752 47844 22756 47900
rect 22692 47840 22756 47844
rect 22772 47900 22836 47904
rect 22772 47844 22776 47900
rect 22776 47844 22832 47900
rect 22832 47844 22836 47900
rect 22772 47840 22836 47844
rect 22852 47900 22916 47904
rect 22852 47844 22856 47900
rect 22856 47844 22912 47900
rect 22912 47844 22916 47900
rect 22852 47840 22916 47844
rect 27612 47900 27676 47904
rect 27612 47844 27616 47900
rect 27616 47844 27672 47900
rect 27672 47844 27676 47900
rect 27612 47840 27676 47844
rect 27692 47900 27756 47904
rect 27692 47844 27696 47900
rect 27696 47844 27752 47900
rect 27752 47844 27756 47900
rect 27692 47840 27756 47844
rect 27772 47900 27836 47904
rect 27772 47844 27776 47900
rect 27776 47844 27832 47900
rect 27832 47844 27836 47900
rect 27772 47840 27836 47844
rect 27852 47900 27916 47904
rect 27852 47844 27856 47900
rect 27856 47844 27912 47900
rect 27912 47844 27916 47900
rect 27852 47840 27916 47844
rect 32612 47900 32676 47904
rect 32612 47844 32616 47900
rect 32616 47844 32672 47900
rect 32672 47844 32676 47900
rect 32612 47840 32676 47844
rect 32692 47900 32756 47904
rect 32692 47844 32696 47900
rect 32696 47844 32752 47900
rect 32752 47844 32756 47900
rect 32692 47840 32756 47844
rect 32772 47900 32836 47904
rect 32772 47844 32776 47900
rect 32776 47844 32832 47900
rect 32832 47844 32836 47900
rect 32772 47840 32836 47844
rect 32852 47900 32916 47904
rect 32852 47844 32856 47900
rect 32856 47844 32912 47900
rect 32912 47844 32916 47900
rect 32852 47840 32916 47844
rect 37612 47900 37676 47904
rect 37612 47844 37616 47900
rect 37616 47844 37672 47900
rect 37672 47844 37676 47900
rect 37612 47840 37676 47844
rect 37692 47900 37756 47904
rect 37692 47844 37696 47900
rect 37696 47844 37752 47900
rect 37752 47844 37756 47900
rect 37692 47840 37756 47844
rect 37772 47900 37836 47904
rect 37772 47844 37776 47900
rect 37776 47844 37832 47900
rect 37832 47844 37836 47900
rect 37772 47840 37836 47844
rect 37852 47900 37916 47904
rect 37852 47844 37856 47900
rect 37856 47844 37912 47900
rect 37912 47844 37916 47900
rect 37852 47840 37916 47844
rect 42612 47900 42676 47904
rect 42612 47844 42616 47900
rect 42616 47844 42672 47900
rect 42672 47844 42676 47900
rect 42612 47840 42676 47844
rect 42692 47900 42756 47904
rect 42692 47844 42696 47900
rect 42696 47844 42752 47900
rect 42752 47844 42756 47900
rect 42692 47840 42756 47844
rect 42772 47900 42836 47904
rect 42772 47844 42776 47900
rect 42776 47844 42832 47900
rect 42832 47844 42836 47900
rect 42772 47840 42836 47844
rect 42852 47900 42916 47904
rect 42852 47844 42856 47900
rect 42856 47844 42912 47900
rect 42912 47844 42916 47900
rect 42852 47840 42916 47844
rect 47612 47900 47676 47904
rect 47612 47844 47616 47900
rect 47616 47844 47672 47900
rect 47672 47844 47676 47900
rect 47612 47840 47676 47844
rect 47692 47900 47756 47904
rect 47692 47844 47696 47900
rect 47696 47844 47752 47900
rect 47752 47844 47756 47900
rect 47692 47840 47756 47844
rect 47772 47900 47836 47904
rect 47772 47844 47776 47900
rect 47776 47844 47832 47900
rect 47832 47844 47836 47900
rect 47772 47840 47836 47844
rect 47852 47900 47916 47904
rect 47852 47844 47856 47900
rect 47856 47844 47912 47900
rect 47912 47844 47916 47900
rect 47852 47840 47916 47844
rect 52612 47900 52676 47904
rect 52612 47844 52616 47900
rect 52616 47844 52672 47900
rect 52672 47844 52676 47900
rect 52612 47840 52676 47844
rect 52692 47900 52756 47904
rect 52692 47844 52696 47900
rect 52696 47844 52752 47900
rect 52752 47844 52756 47900
rect 52692 47840 52756 47844
rect 52772 47900 52836 47904
rect 52772 47844 52776 47900
rect 52776 47844 52832 47900
rect 52832 47844 52836 47900
rect 52772 47840 52836 47844
rect 52852 47900 52916 47904
rect 52852 47844 52856 47900
rect 52856 47844 52912 47900
rect 52912 47844 52916 47900
rect 52852 47840 52916 47844
rect 57612 47900 57676 47904
rect 57612 47844 57616 47900
rect 57616 47844 57672 47900
rect 57672 47844 57676 47900
rect 57612 47840 57676 47844
rect 57692 47900 57756 47904
rect 57692 47844 57696 47900
rect 57696 47844 57752 47900
rect 57752 47844 57756 47900
rect 57692 47840 57756 47844
rect 57772 47900 57836 47904
rect 57772 47844 57776 47900
rect 57776 47844 57832 47900
rect 57832 47844 57836 47900
rect 57772 47840 57836 47844
rect 57852 47900 57916 47904
rect 57852 47844 57856 47900
rect 57856 47844 57912 47900
rect 57912 47844 57916 47900
rect 57852 47840 57916 47844
rect 1952 47356 2016 47360
rect 1952 47300 1956 47356
rect 1956 47300 2012 47356
rect 2012 47300 2016 47356
rect 1952 47296 2016 47300
rect 2032 47356 2096 47360
rect 2032 47300 2036 47356
rect 2036 47300 2092 47356
rect 2092 47300 2096 47356
rect 2032 47296 2096 47300
rect 2112 47356 2176 47360
rect 2112 47300 2116 47356
rect 2116 47300 2172 47356
rect 2172 47300 2176 47356
rect 2112 47296 2176 47300
rect 2192 47356 2256 47360
rect 2192 47300 2196 47356
rect 2196 47300 2252 47356
rect 2252 47300 2256 47356
rect 2192 47296 2256 47300
rect 6952 47356 7016 47360
rect 6952 47300 6956 47356
rect 6956 47300 7012 47356
rect 7012 47300 7016 47356
rect 6952 47296 7016 47300
rect 7032 47356 7096 47360
rect 7032 47300 7036 47356
rect 7036 47300 7092 47356
rect 7092 47300 7096 47356
rect 7032 47296 7096 47300
rect 7112 47356 7176 47360
rect 7112 47300 7116 47356
rect 7116 47300 7172 47356
rect 7172 47300 7176 47356
rect 7112 47296 7176 47300
rect 7192 47356 7256 47360
rect 7192 47300 7196 47356
rect 7196 47300 7252 47356
rect 7252 47300 7256 47356
rect 7192 47296 7256 47300
rect 11952 47356 12016 47360
rect 11952 47300 11956 47356
rect 11956 47300 12012 47356
rect 12012 47300 12016 47356
rect 11952 47296 12016 47300
rect 12032 47356 12096 47360
rect 12032 47300 12036 47356
rect 12036 47300 12092 47356
rect 12092 47300 12096 47356
rect 12032 47296 12096 47300
rect 12112 47356 12176 47360
rect 12112 47300 12116 47356
rect 12116 47300 12172 47356
rect 12172 47300 12176 47356
rect 12112 47296 12176 47300
rect 12192 47356 12256 47360
rect 12192 47300 12196 47356
rect 12196 47300 12252 47356
rect 12252 47300 12256 47356
rect 12192 47296 12256 47300
rect 16952 47356 17016 47360
rect 16952 47300 16956 47356
rect 16956 47300 17012 47356
rect 17012 47300 17016 47356
rect 16952 47296 17016 47300
rect 17032 47356 17096 47360
rect 17032 47300 17036 47356
rect 17036 47300 17092 47356
rect 17092 47300 17096 47356
rect 17032 47296 17096 47300
rect 17112 47356 17176 47360
rect 17112 47300 17116 47356
rect 17116 47300 17172 47356
rect 17172 47300 17176 47356
rect 17112 47296 17176 47300
rect 17192 47356 17256 47360
rect 17192 47300 17196 47356
rect 17196 47300 17252 47356
rect 17252 47300 17256 47356
rect 17192 47296 17256 47300
rect 21952 47356 22016 47360
rect 21952 47300 21956 47356
rect 21956 47300 22012 47356
rect 22012 47300 22016 47356
rect 21952 47296 22016 47300
rect 22032 47356 22096 47360
rect 22032 47300 22036 47356
rect 22036 47300 22092 47356
rect 22092 47300 22096 47356
rect 22032 47296 22096 47300
rect 22112 47356 22176 47360
rect 22112 47300 22116 47356
rect 22116 47300 22172 47356
rect 22172 47300 22176 47356
rect 22112 47296 22176 47300
rect 22192 47356 22256 47360
rect 22192 47300 22196 47356
rect 22196 47300 22252 47356
rect 22252 47300 22256 47356
rect 22192 47296 22256 47300
rect 26952 47356 27016 47360
rect 26952 47300 26956 47356
rect 26956 47300 27012 47356
rect 27012 47300 27016 47356
rect 26952 47296 27016 47300
rect 27032 47356 27096 47360
rect 27032 47300 27036 47356
rect 27036 47300 27092 47356
rect 27092 47300 27096 47356
rect 27032 47296 27096 47300
rect 27112 47356 27176 47360
rect 27112 47300 27116 47356
rect 27116 47300 27172 47356
rect 27172 47300 27176 47356
rect 27112 47296 27176 47300
rect 27192 47356 27256 47360
rect 27192 47300 27196 47356
rect 27196 47300 27252 47356
rect 27252 47300 27256 47356
rect 27192 47296 27256 47300
rect 31952 47356 32016 47360
rect 31952 47300 31956 47356
rect 31956 47300 32012 47356
rect 32012 47300 32016 47356
rect 31952 47296 32016 47300
rect 32032 47356 32096 47360
rect 32032 47300 32036 47356
rect 32036 47300 32092 47356
rect 32092 47300 32096 47356
rect 32032 47296 32096 47300
rect 32112 47356 32176 47360
rect 32112 47300 32116 47356
rect 32116 47300 32172 47356
rect 32172 47300 32176 47356
rect 32112 47296 32176 47300
rect 32192 47356 32256 47360
rect 32192 47300 32196 47356
rect 32196 47300 32252 47356
rect 32252 47300 32256 47356
rect 32192 47296 32256 47300
rect 36952 47356 37016 47360
rect 36952 47300 36956 47356
rect 36956 47300 37012 47356
rect 37012 47300 37016 47356
rect 36952 47296 37016 47300
rect 37032 47356 37096 47360
rect 37032 47300 37036 47356
rect 37036 47300 37092 47356
rect 37092 47300 37096 47356
rect 37032 47296 37096 47300
rect 37112 47356 37176 47360
rect 37112 47300 37116 47356
rect 37116 47300 37172 47356
rect 37172 47300 37176 47356
rect 37112 47296 37176 47300
rect 37192 47356 37256 47360
rect 37192 47300 37196 47356
rect 37196 47300 37252 47356
rect 37252 47300 37256 47356
rect 37192 47296 37256 47300
rect 41952 47356 42016 47360
rect 41952 47300 41956 47356
rect 41956 47300 42012 47356
rect 42012 47300 42016 47356
rect 41952 47296 42016 47300
rect 42032 47356 42096 47360
rect 42032 47300 42036 47356
rect 42036 47300 42092 47356
rect 42092 47300 42096 47356
rect 42032 47296 42096 47300
rect 42112 47356 42176 47360
rect 42112 47300 42116 47356
rect 42116 47300 42172 47356
rect 42172 47300 42176 47356
rect 42112 47296 42176 47300
rect 42192 47356 42256 47360
rect 42192 47300 42196 47356
rect 42196 47300 42252 47356
rect 42252 47300 42256 47356
rect 42192 47296 42256 47300
rect 46952 47356 47016 47360
rect 46952 47300 46956 47356
rect 46956 47300 47012 47356
rect 47012 47300 47016 47356
rect 46952 47296 47016 47300
rect 47032 47356 47096 47360
rect 47032 47300 47036 47356
rect 47036 47300 47092 47356
rect 47092 47300 47096 47356
rect 47032 47296 47096 47300
rect 47112 47356 47176 47360
rect 47112 47300 47116 47356
rect 47116 47300 47172 47356
rect 47172 47300 47176 47356
rect 47112 47296 47176 47300
rect 47192 47356 47256 47360
rect 47192 47300 47196 47356
rect 47196 47300 47252 47356
rect 47252 47300 47256 47356
rect 47192 47296 47256 47300
rect 51952 47356 52016 47360
rect 51952 47300 51956 47356
rect 51956 47300 52012 47356
rect 52012 47300 52016 47356
rect 51952 47296 52016 47300
rect 52032 47356 52096 47360
rect 52032 47300 52036 47356
rect 52036 47300 52092 47356
rect 52092 47300 52096 47356
rect 52032 47296 52096 47300
rect 52112 47356 52176 47360
rect 52112 47300 52116 47356
rect 52116 47300 52172 47356
rect 52172 47300 52176 47356
rect 52112 47296 52176 47300
rect 52192 47356 52256 47360
rect 52192 47300 52196 47356
rect 52196 47300 52252 47356
rect 52252 47300 52256 47356
rect 52192 47296 52256 47300
rect 56952 47356 57016 47360
rect 56952 47300 56956 47356
rect 56956 47300 57012 47356
rect 57012 47300 57016 47356
rect 56952 47296 57016 47300
rect 57032 47356 57096 47360
rect 57032 47300 57036 47356
rect 57036 47300 57092 47356
rect 57092 47300 57096 47356
rect 57032 47296 57096 47300
rect 57112 47356 57176 47360
rect 57112 47300 57116 47356
rect 57116 47300 57172 47356
rect 57172 47300 57176 47356
rect 57112 47296 57176 47300
rect 57192 47356 57256 47360
rect 57192 47300 57196 47356
rect 57196 47300 57252 47356
rect 57252 47300 57256 47356
rect 57192 47296 57256 47300
rect 2612 46812 2676 46816
rect 2612 46756 2616 46812
rect 2616 46756 2672 46812
rect 2672 46756 2676 46812
rect 2612 46752 2676 46756
rect 2692 46812 2756 46816
rect 2692 46756 2696 46812
rect 2696 46756 2752 46812
rect 2752 46756 2756 46812
rect 2692 46752 2756 46756
rect 2772 46812 2836 46816
rect 2772 46756 2776 46812
rect 2776 46756 2832 46812
rect 2832 46756 2836 46812
rect 2772 46752 2836 46756
rect 2852 46812 2916 46816
rect 2852 46756 2856 46812
rect 2856 46756 2912 46812
rect 2912 46756 2916 46812
rect 2852 46752 2916 46756
rect 7612 46812 7676 46816
rect 7612 46756 7616 46812
rect 7616 46756 7672 46812
rect 7672 46756 7676 46812
rect 7612 46752 7676 46756
rect 7692 46812 7756 46816
rect 7692 46756 7696 46812
rect 7696 46756 7752 46812
rect 7752 46756 7756 46812
rect 7692 46752 7756 46756
rect 7772 46812 7836 46816
rect 7772 46756 7776 46812
rect 7776 46756 7832 46812
rect 7832 46756 7836 46812
rect 7772 46752 7836 46756
rect 7852 46812 7916 46816
rect 7852 46756 7856 46812
rect 7856 46756 7912 46812
rect 7912 46756 7916 46812
rect 7852 46752 7916 46756
rect 12612 46812 12676 46816
rect 12612 46756 12616 46812
rect 12616 46756 12672 46812
rect 12672 46756 12676 46812
rect 12612 46752 12676 46756
rect 12692 46812 12756 46816
rect 12692 46756 12696 46812
rect 12696 46756 12752 46812
rect 12752 46756 12756 46812
rect 12692 46752 12756 46756
rect 12772 46812 12836 46816
rect 12772 46756 12776 46812
rect 12776 46756 12832 46812
rect 12832 46756 12836 46812
rect 12772 46752 12836 46756
rect 12852 46812 12916 46816
rect 12852 46756 12856 46812
rect 12856 46756 12912 46812
rect 12912 46756 12916 46812
rect 12852 46752 12916 46756
rect 17612 46812 17676 46816
rect 17612 46756 17616 46812
rect 17616 46756 17672 46812
rect 17672 46756 17676 46812
rect 17612 46752 17676 46756
rect 17692 46812 17756 46816
rect 17692 46756 17696 46812
rect 17696 46756 17752 46812
rect 17752 46756 17756 46812
rect 17692 46752 17756 46756
rect 17772 46812 17836 46816
rect 17772 46756 17776 46812
rect 17776 46756 17832 46812
rect 17832 46756 17836 46812
rect 17772 46752 17836 46756
rect 17852 46812 17916 46816
rect 17852 46756 17856 46812
rect 17856 46756 17912 46812
rect 17912 46756 17916 46812
rect 17852 46752 17916 46756
rect 22612 46812 22676 46816
rect 22612 46756 22616 46812
rect 22616 46756 22672 46812
rect 22672 46756 22676 46812
rect 22612 46752 22676 46756
rect 22692 46812 22756 46816
rect 22692 46756 22696 46812
rect 22696 46756 22752 46812
rect 22752 46756 22756 46812
rect 22692 46752 22756 46756
rect 22772 46812 22836 46816
rect 22772 46756 22776 46812
rect 22776 46756 22832 46812
rect 22832 46756 22836 46812
rect 22772 46752 22836 46756
rect 22852 46812 22916 46816
rect 22852 46756 22856 46812
rect 22856 46756 22912 46812
rect 22912 46756 22916 46812
rect 22852 46752 22916 46756
rect 27612 46812 27676 46816
rect 27612 46756 27616 46812
rect 27616 46756 27672 46812
rect 27672 46756 27676 46812
rect 27612 46752 27676 46756
rect 27692 46812 27756 46816
rect 27692 46756 27696 46812
rect 27696 46756 27752 46812
rect 27752 46756 27756 46812
rect 27692 46752 27756 46756
rect 27772 46812 27836 46816
rect 27772 46756 27776 46812
rect 27776 46756 27832 46812
rect 27832 46756 27836 46812
rect 27772 46752 27836 46756
rect 27852 46812 27916 46816
rect 27852 46756 27856 46812
rect 27856 46756 27912 46812
rect 27912 46756 27916 46812
rect 27852 46752 27916 46756
rect 32612 46812 32676 46816
rect 32612 46756 32616 46812
rect 32616 46756 32672 46812
rect 32672 46756 32676 46812
rect 32612 46752 32676 46756
rect 32692 46812 32756 46816
rect 32692 46756 32696 46812
rect 32696 46756 32752 46812
rect 32752 46756 32756 46812
rect 32692 46752 32756 46756
rect 32772 46812 32836 46816
rect 32772 46756 32776 46812
rect 32776 46756 32832 46812
rect 32832 46756 32836 46812
rect 32772 46752 32836 46756
rect 32852 46812 32916 46816
rect 32852 46756 32856 46812
rect 32856 46756 32912 46812
rect 32912 46756 32916 46812
rect 32852 46752 32916 46756
rect 37612 46812 37676 46816
rect 37612 46756 37616 46812
rect 37616 46756 37672 46812
rect 37672 46756 37676 46812
rect 37612 46752 37676 46756
rect 37692 46812 37756 46816
rect 37692 46756 37696 46812
rect 37696 46756 37752 46812
rect 37752 46756 37756 46812
rect 37692 46752 37756 46756
rect 37772 46812 37836 46816
rect 37772 46756 37776 46812
rect 37776 46756 37832 46812
rect 37832 46756 37836 46812
rect 37772 46752 37836 46756
rect 37852 46812 37916 46816
rect 37852 46756 37856 46812
rect 37856 46756 37912 46812
rect 37912 46756 37916 46812
rect 37852 46752 37916 46756
rect 42612 46812 42676 46816
rect 42612 46756 42616 46812
rect 42616 46756 42672 46812
rect 42672 46756 42676 46812
rect 42612 46752 42676 46756
rect 42692 46812 42756 46816
rect 42692 46756 42696 46812
rect 42696 46756 42752 46812
rect 42752 46756 42756 46812
rect 42692 46752 42756 46756
rect 42772 46812 42836 46816
rect 42772 46756 42776 46812
rect 42776 46756 42832 46812
rect 42832 46756 42836 46812
rect 42772 46752 42836 46756
rect 42852 46812 42916 46816
rect 42852 46756 42856 46812
rect 42856 46756 42912 46812
rect 42912 46756 42916 46812
rect 42852 46752 42916 46756
rect 47612 46812 47676 46816
rect 47612 46756 47616 46812
rect 47616 46756 47672 46812
rect 47672 46756 47676 46812
rect 47612 46752 47676 46756
rect 47692 46812 47756 46816
rect 47692 46756 47696 46812
rect 47696 46756 47752 46812
rect 47752 46756 47756 46812
rect 47692 46752 47756 46756
rect 47772 46812 47836 46816
rect 47772 46756 47776 46812
rect 47776 46756 47832 46812
rect 47832 46756 47836 46812
rect 47772 46752 47836 46756
rect 47852 46812 47916 46816
rect 47852 46756 47856 46812
rect 47856 46756 47912 46812
rect 47912 46756 47916 46812
rect 47852 46752 47916 46756
rect 52612 46812 52676 46816
rect 52612 46756 52616 46812
rect 52616 46756 52672 46812
rect 52672 46756 52676 46812
rect 52612 46752 52676 46756
rect 52692 46812 52756 46816
rect 52692 46756 52696 46812
rect 52696 46756 52752 46812
rect 52752 46756 52756 46812
rect 52692 46752 52756 46756
rect 52772 46812 52836 46816
rect 52772 46756 52776 46812
rect 52776 46756 52832 46812
rect 52832 46756 52836 46812
rect 52772 46752 52836 46756
rect 52852 46812 52916 46816
rect 52852 46756 52856 46812
rect 52856 46756 52912 46812
rect 52912 46756 52916 46812
rect 52852 46752 52916 46756
rect 57612 46812 57676 46816
rect 57612 46756 57616 46812
rect 57616 46756 57672 46812
rect 57672 46756 57676 46812
rect 57612 46752 57676 46756
rect 57692 46812 57756 46816
rect 57692 46756 57696 46812
rect 57696 46756 57752 46812
rect 57752 46756 57756 46812
rect 57692 46752 57756 46756
rect 57772 46812 57836 46816
rect 57772 46756 57776 46812
rect 57776 46756 57832 46812
rect 57832 46756 57836 46812
rect 57772 46752 57836 46756
rect 57852 46812 57916 46816
rect 57852 46756 57856 46812
rect 57856 46756 57912 46812
rect 57912 46756 57916 46812
rect 57852 46752 57916 46756
rect 1952 46268 2016 46272
rect 1952 46212 1956 46268
rect 1956 46212 2012 46268
rect 2012 46212 2016 46268
rect 1952 46208 2016 46212
rect 2032 46268 2096 46272
rect 2032 46212 2036 46268
rect 2036 46212 2092 46268
rect 2092 46212 2096 46268
rect 2032 46208 2096 46212
rect 2112 46268 2176 46272
rect 2112 46212 2116 46268
rect 2116 46212 2172 46268
rect 2172 46212 2176 46268
rect 2112 46208 2176 46212
rect 2192 46268 2256 46272
rect 2192 46212 2196 46268
rect 2196 46212 2252 46268
rect 2252 46212 2256 46268
rect 2192 46208 2256 46212
rect 6952 46268 7016 46272
rect 6952 46212 6956 46268
rect 6956 46212 7012 46268
rect 7012 46212 7016 46268
rect 6952 46208 7016 46212
rect 7032 46268 7096 46272
rect 7032 46212 7036 46268
rect 7036 46212 7092 46268
rect 7092 46212 7096 46268
rect 7032 46208 7096 46212
rect 7112 46268 7176 46272
rect 7112 46212 7116 46268
rect 7116 46212 7172 46268
rect 7172 46212 7176 46268
rect 7112 46208 7176 46212
rect 7192 46268 7256 46272
rect 7192 46212 7196 46268
rect 7196 46212 7252 46268
rect 7252 46212 7256 46268
rect 7192 46208 7256 46212
rect 11952 46268 12016 46272
rect 11952 46212 11956 46268
rect 11956 46212 12012 46268
rect 12012 46212 12016 46268
rect 11952 46208 12016 46212
rect 12032 46268 12096 46272
rect 12032 46212 12036 46268
rect 12036 46212 12092 46268
rect 12092 46212 12096 46268
rect 12032 46208 12096 46212
rect 12112 46268 12176 46272
rect 12112 46212 12116 46268
rect 12116 46212 12172 46268
rect 12172 46212 12176 46268
rect 12112 46208 12176 46212
rect 12192 46268 12256 46272
rect 12192 46212 12196 46268
rect 12196 46212 12252 46268
rect 12252 46212 12256 46268
rect 12192 46208 12256 46212
rect 16952 46268 17016 46272
rect 16952 46212 16956 46268
rect 16956 46212 17012 46268
rect 17012 46212 17016 46268
rect 16952 46208 17016 46212
rect 17032 46268 17096 46272
rect 17032 46212 17036 46268
rect 17036 46212 17092 46268
rect 17092 46212 17096 46268
rect 17032 46208 17096 46212
rect 17112 46268 17176 46272
rect 17112 46212 17116 46268
rect 17116 46212 17172 46268
rect 17172 46212 17176 46268
rect 17112 46208 17176 46212
rect 17192 46268 17256 46272
rect 17192 46212 17196 46268
rect 17196 46212 17252 46268
rect 17252 46212 17256 46268
rect 17192 46208 17256 46212
rect 21952 46268 22016 46272
rect 21952 46212 21956 46268
rect 21956 46212 22012 46268
rect 22012 46212 22016 46268
rect 21952 46208 22016 46212
rect 22032 46268 22096 46272
rect 22032 46212 22036 46268
rect 22036 46212 22092 46268
rect 22092 46212 22096 46268
rect 22032 46208 22096 46212
rect 22112 46268 22176 46272
rect 22112 46212 22116 46268
rect 22116 46212 22172 46268
rect 22172 46212 22176 46268
rect 22112 46208 22176 46212
rect 22192 46268 22256 46272
rect 22192 46212 22196 46268
rect 22196 46212 22252 46268
rect 22252 46212 22256 46268
rect 22192 46208 22256 46212
rect 26952 46268 27016 46272
rect 26952 46212 26956 46268
rect 26956 46212 27012 46268
rect 27012 46212 27016 46268
rect 26952 46208 27016 46212
rect 27032 46268 27096 46272
rect 27032 46212 27036 46268
rect 27036 46212 27092 46268
rect 27092 46212 27096 46268
rect 27032 46208 27096 46212
rect 27112 46268 27176 46272
rect 27112 46212 27116 46268
rect 27116 46212 27172 46268
rect 27172 46212 27176 46268
rect 27112 46208 27176 46212
rect 27192 46268 27256 46272
rect 27192 46212 27196 46268
rect 27196 46212 27252 46268
rect 27252 46212 27256 46268
rect 27192 46208 27256 46212
rect 31952 46268 32016 46272
rect 31952 46212 31956 46268
rect 31956 46212 32012 46268
rect 32012 46212 32016 46268
rect 31952 46208 32016 46212
rect 32032 46268 32096 46272
rect 32032 46212 32036 46268
rect 32036 46212 32092 46268
rect 32092 46212 32096 46268
rect 32032 46208 32096 46212
rect 32112 46268 32176 46272
rect 32112 46212 32116 46268
rect 32116 46212 32172 46268
rect 32172 46212 32176 46268
rect 32112 46208 32176 46212
rect 32192 46268 32256 46272
rect 32192 46212 32196 46268
rect 32196 46212 32252 46268
rect 32252 46212 32256 46268
rect 32192 46208 32256 46212
rect 36952 46268 37016 46272
rect 36952 46212 36956 46268
rect 36956 46212 37012 46268
rect 37012 46212 37016 46268
rect 36952 46208 37016 46212
rect 37032 46268 37096 46272
rect 37032 46212 37036 46268
rect 37036 46212 37092 46268
rect 37092 46212 37096 46268
rect 37032 46208 37096 46212
rect 37112 46268 37176 46272
rect 37112 46212 37116 46268
rect 37116 46212 37172 46268
rect 37172 46212 37176 46268
rect 37112 46208 37176 46212
rect 37192 46268 37256 46272
rect 37192 46212 37196 46268
rect 37196 46212 37252 46268
rect 37252 46212 37256 46268
rect 37192 46208 37256 46212
rect 41952 46268 42016 46272
rect 41952 46212 41956 46268
rect 41956 46212 42012 46268
rect 42012 46212 42016 46268
rect 41952 46208 42016 46212
rect 42032 46268 42096 46272
rect 42032 46212 42036 46268
rect 42036 46212 42092 46268
rect 42092 46212 42096 46268
rect 42032 46208 42096 46212
rect 42112 46268 42176 46272
rect 42112 46212 42116 46268
rect 42116 46212 42172 46268
rect 42172 46212 42176 46268
rect 42112 46208 42176 46212
rect 42192 46268 42256 46272
rect 42192 46212 42196 46268
rect 42196 46212 42252 46268
rect 42252 46212 42256 46268
rect 42192 46208 42256 46212
rect 46952 46268 47016 46272
rect 46952 46212 46956 46268
rect 46956 46212 47012 46268
rect 47012 46212 47016 46268
rect 46952 46208 47016 46212
rect 47032 46268 47096 46272
rect 47032 46212 47036 46268
rect 47036 46212 47092 46268
rect 47092 46212 47096 46268
rect 47032 46208 47096 46212
rect 47112 46268 47176 46272
rect 47112 46212 47116 46268
rect 47116 46212 47172 46268
rect 47172 46212 47176 46268
rect 47112 46208 47176 46212
rect 47192 46268 47256 46272
rect 47192 46212 47196 46268
rect 47196 46212 47252 46268
rect 47252 46212 47256 46268
rect 47192 46208 47256 46212
rect 51952 46268 52016 46272
rect 51952 46212 51956 46268
rect 51956 46212 52012 46268
rect 52012 46212 52016 46268
rect 51952 46208 52016 46212
rect 52032 46268 52096 46272
rect 52032 46212 52036 46268
rect 52036 46212 52092 46268
rect 52092 46212 52096 46268
rect 52032 46208 52096 46212
rect 52112 46268 52176 46272
rect 52112 46212 52116 46268
rect 52116 46212 52172 46268
rect 52172 46212 52176 46268
rect 52112 46208 52176 46212
rect 52192 46268 52256 46272
rect 52192 46212 52196 46268
rect 52196 46212 52252 46268
rect 52252 46212 52256 46268
rect 52192 46208 52256 46212
rect 56952 46268 57016 46272
rect 56952 46212 56956 46268
rect 56956 46212 57012 46268
rect 57012 46212 57016 46268
rect 56952 46208 57016 46212
rect 57032 46268 57096 46272
rect 57032 46212 57036 46268
rect 57036 46212 57092 46268
rect 57092 46212 57096 46268
rect 57032 46208 57096 46212
rect 57112 46268 57176 46272
rect 57112 46212 57116 46268
rect 57116 46212 57172 46268
rect 57172 46212 57176 46268
rect 57112 46208 57176 46212
rect 57192 46268 57256 46272
rect 57192 46212 57196 46268
rect 57196 46212 57252 46268
rect 57252 46212 57256 46268
rect 57192 46208 57256 46212
rect 2612 45724 2676 45728
rect 2612 45668 2616 45724
rect 2616 45668 2672 45724
rect 2672 45668 2676 45724
rect 2612 45664 2676 45668
rect 2692 45724 2756 45728
rect 2692 45668 2696 45724
rect 2696 45668 2752 45724
rect 2752 45668 2756 45724
rect 2692 45664 2756 45668
rect 2772 45724 2836 45728
rect 2772 45668 2776 45724
rect 2776 45668 2832 45724
rect 2832 45668 2836 45724
rect 2772 45664 2836 45668
rect 2852 45724 2916 45728
rect 2852 45668 2856 45724
rect 2856 45668 2912 45724
rect 2912 45668 2916 45724
rect 2852 45664 2916 45668
rect 7612 45724 7676 45728
rect 7612 45668 7616 45724
rect 7616 45668 7672 45724
rect 7672 45668 7676 45724
rect 7612 45664 7676 45668
rect 7692 45724 7756 45728
rect 7692 45668 7696 45724
rect 7696 45668 7752 45724
rect 7752 45668 7756 45724
rect 7692 45664 7756 45668
rect 7772 45724 7836 45728
rect 7772 45668 7776 45724
rect 7776 45668 7832 45724
rect 7832 45668 7836 45724
rect 7772 45664 7836 45668
rect 7852 45724 7916 45728
rect 7852 45668 7856 45724
rect 7856 45668 7912 45724
rect 7912 45668 7916 45724
rect 7852 45664 7916 45668
rect 12612 45724 12676 45728
rect 12612 45668 12616 45724
rect 12616 45668 12672 45724
rect 12672 45668 12676 45724
rect 12612 45664 12676 45668
rect 12692 45724 12756 45728
rect 12692 45668 12696 45724
rect 12696 45668 12752 45724
rect 12752 45668 12756 45724
rect 12692 45664 12756 45668
rect 12772 45724 12836 45728
rect 12772 45668 12776 45724
rect 12776 45668 12832 45724
rect 12832 45668 12836 45724
rect 12772 45664 12836 45668
rect 12852 45724 12916 45728
rect 12852 45668 12856 45724
rect 12856 45668 12912 45724
rect 12912 45668 12916 45724
rect 12852 45664 12916 45668
rect 17612 45724 17676 45728
rect 17612 45668 17616 45724
rect 17616 45668 17672 45724
rect 17672 45668 17676 45724
rect 17612 45664 17676 45668
rect 17692 45724 17756 45728
rect 17692 45668 17696 45724
rect 17696 45668 17752 45724
rect 17752 45668 17756 45724
rect 17692 45664 17756 45668
rect 17772 45724 17836 45728
rect 17772 45668 17776 45724
rect 17776 45668 17832 45724
rect 17832 45668 17836 45724
rect 17772 45664 17836 45668
rect 17852 45724 17916 45728
rect 17852 45668 17856 45724
rect 17856 45668 17912 45724
rect 17912 45668 17916 45724
rect 17852 45664 17916 45668
rect 22612 45724 22676 45728
rect 22612 45668 22616 45724
rect 22616 45668 22672 45724
rect 22672 45668 22676 45724
rect 22612 45664 22676 45668
rect 22692 45724 22756 45728
rect 22692 45668 22696 45724
rect 22696 45668 22752 45724
rect 22752 45668 22756 45724
rect 22692 45664 22756 45668
rect 22772 45724 22836 45728
rect 22772 45668 22776 45724
rect 22776 45668 22832 45724
rect 22832 45668 22836 45724
rect 22772 45664 22836 45668
rect 22852 45724 22916 45728
rect 22852 45668 22856 45724
rect 22856 45668 22912 45724
rect 22912 45668 22916 45724
rect 22852 45664 22916 45668
rect 27612 45724 27676 45728
rect 27612 45668 27616 45724
rect 27616 45668 27672 45724
rect 27672 45668 27676 45724
rect 27612 45664 27676 45668
rect 27692 45724 27756 45728
rect 27692 45668 27696 45724
rect 27696 45668 27752 45724
rect 27752 45668 27756 45724
rect 27692 45664 27756 45668
rect 27772 45724 27836 45728
rect 27772 45668 27776 45724
rect 27776 45668 27832 45724
rect 27832 45668 27836 45724
rect 27772 45664 27836 45668
rect 27852 45724 27916 45728
rect 27852 45668 27856 45724
rect 27856 45668 27912 45724
rect 27912 45668 27916 45724
rect 27852 45664 27916 45668
rect 32612 45724 32676 45728
rect 32612 45668 32616 45724
rect 32616 45668 32672 45724
rect 32672 45668 32676 45724
rect 32612 45664 32676 45668
rect 32692 45724 32756 45728
rect 32692 45668 32696 45724
rect 32696 45668 32752 45724
rect 32752 45668 32756 45724
rect 32692 45664 32756 45668
rect 32772 45724 32836 45728
rect 32772 45668 32776 45724
rect 32776 45668 32832 45724
rect 32832 45668 32836 45724
rect 32772 45664 32836 45668
rect 32852 45724 32916 45728
rect 32852 45668 32856 45724
rect 32856 45668 32912 45724
rect 32912 45668 32916 45724
rect 32852 45664 32916 45668
rect 37612 45724 37676 45728
rect 37612 45668 37616 45724
rect 37616 45668 37672 45724
rect 37672 45668 37676 45724
rect 37612 45664 37676 45668
rect 37692 45724 37756 45728
rect 37692 45668 37696 45724
rect 37696 45668 37752 45724
rect 37752 45668 37756 45724
rect 37692 45664 37756 45668
rect 37772 45724 37836 45728
rect 37772 45668 37776 45724
rect 37776 45668 37832 45724
rect 37832 45668 37836 45724
rect 37772 45664 37836 45668
rect 37852 45724 37916 45728
rect 37852 45668 37856 45724
rect 37856 45668 37912 45724
rect 37912 45668 37916 45724
rect 37852 45664 37916 45668
rect 42612 45724 42676 45728
rect 42612 45668 42616 45724
rect 42616 45668 42672 45724
rect 42672 45668 42676 45724
rect 42612 45664 42676 45668
rect 42692 45724 42756 45728
rect 42692 45668 42696 45724
rect 42696 45668 42752 45724
rect 42752 45668 42756 45724
rect 42692 45664 42756 45668
rect 42772 45724 42836 45728
rect 42772 45668 42776 45724
rect 42776 45668 42832 45724
rect 42832 45668 42836 45724
rect 42772 45664 42836 45668
rect 42852 45724 42916 45728
rect 42852 45668 42856 45724
rect 42856 45668 42912 45724
rect 42912 45668 42916 45724
rect 42852 45664 42916 45668
rect 47612 45724 47676 45728
rect 47612 45668 47616 45724
rect 47616 45668 47672 45724
rect 47672 45668 47676 45724
rect 47612 45664 47676 45668
rect 47692 45724 47756 45728
rect 47692 45668 47696 45724
rect 47696 45668 47752 45724
rect 47752 45668 47756 45724
rect 47692 45664 47756 45668
rect 47772 45724 47836 45728
rect 47772 45668 47776 45724
rect 47776 45668 47832 45724
rect 47832 45668 47836 45724
rect 47772 45664 47836 45668
rect 47852 45724 47916 45728
rect 47852 45668 47856 45724
rect 47856 45668 47912 45724
rect 47912 45668 47916 45724
rect 47852 45664 47916 45668
rect 52612 45724 52676 45728
rect 52612 45668 52616 45724
rect 52616 45668 52672 45724
rect 52672 45668 52676 45724
rect 52612 45664 52676 45668
rect 52692 45724 52756 45728
rect 52692 45668 52696 45724
rect 52696 45668 52752 45724
rect 52752 45668 52756 45724
rect 52692 45664 52756 45668
rect 52772 45724 52836 45728
rect 52772 45668 52776 45724
rect 52776 45668 52832 45724
rect 52832 45668 52836 45724
rect 52772 45664 52836 45668
rect 52852 45724 52916 45728
rect 52852 45668 52856 45724
rect 52856 45668 52912 45724
rect 52912 45668 52916 45724
rect 52852 45664 52916 45668
rect 57612 45724 57676 45728
rect 57612 45668 57616 45724
rect 57616 45668 57672 45724
rect 57672 45668 57676 45724
rect 57612 45664 57676 45668
rect 57692 45724 57756 45728
rect 57692 45668 57696 45724
rect 57696 45668 57752 45724
rect 57752 45668 57756 45724
rect 57692 45664 57756 45668
rect 57772 45724 57836 45728
rect 57772 45668 57776 45724
rect 57776 45668 57832 45724
rect 57832 45668 57836 45724
rect 57772 45664 57836 45668
rect 57852 45724 57916 45728
rect 57852 45668 57856 45724
rect 57856 45668 57912 45724
rect 57912 45668 57916 45724
rect 57852 45664 57916 45668
rect 1952 45180 2016 45184
rect 1952 45124 1956 45180
rect 1956 45124 2012 45180
rect 2012 45124 2016 45180
rect 1952 45120 2016 45124
rect 2032 45180 2096 45184
rect 2032 45124 2036 45180
rect 2036 45124 2092 45180
rect 2092 45124 2096 45180
rect 2032 45120 2096 45124
rect 2112 45180 2176 45184
rect 2112 45124 2116 45180
rect 2116 45124 2172 45180
rect 2172 45124 2176 45180
rect 2112 45120 2176 45124
rect 2192 45180 2256 45184
rect 2192 45124 2196 45180
rect 2196 45124 2252 45180
rect 2252 45124 2256 45180
rect 2192 45120 2256 45124
rect 6952 45180 7016 45184
rect 6952 45124 6956 45180
rect 6956 45124 7012 45180
rect 7012 45124 7016 45180
rect 6952 45120 7016 45124
rect 7032 45180 7096 45184
rect 7032 45124 7036 45180
rect 7036 45124 7092 45180
rect 7092 45124 7096 45180
rect 7032 45120 7096 45124
rect 7112 45180 7176 45184
rect 7112 45124 7116 45180
rect 7116 45124 7172 45180
rect 7172 45124 7176 45180
rect 7112 45120 7176 45124
rect 7192 45180 7256 45184
rect 7192 45124 7196 45180
rect 7196 45124 7252 45180
rect 7252 45124 7256 45180
rect 7192 45120 7256 45124
rect 11952 45180 12016 45184
rect 11952 45124 11956 45180
rect 11956 45124 12012 45180
rect 12012 45124 12016 45180
rect 11952 45120 12016 45124
rect 12032 45180 12096 45184
rect 12032 45124 12036 45180
rect 12036 45124 12092 45180
rect 12092 45124 12096 45180
rect 12032 45120 12096 45124
rect 12112 45180 12176 45184
rect 12112 45124 12116 45180
rect 12116 45124 12172 45180
rect 12172 45124 12176 45180
rect 12112 45120 12176 45124
rect 12192 45180 12256 45184
rect 12192 45124 12196 45180
rect 12196 45124 12252 45180
rect 12252 45124 12256 45180
rect 12192 45120 12256 45124
rect 16952 45180 17016 45184
rect 16952 45124 16956 45180
rect 16956 45124 17012 45180
rect 17012 45124 17016 45180
rect 16952 45120 17016 45124
rect 17032 45180 17096 45184
rect 17032 45124 17036 45180
rect 17036 45124 17092 45180
rect 17092 45124 17096 45180
rect 17032 45120 17096 45124
rect 17112 45180 17176 45184
rect 17112 45124 17116 45180
rect 17116 45124 17172 45180
rect 17172 45124 17176 45180
rect 17112 45120 17176 45124
rect 17192 45180 17256 45184
rect 17192 45124 17196 45180
rect 17196 45124 17252 45180
rect 17252 45124 17256 45180
rect 17192 45120 17256 45124
rect 21952 45180 22016 45184
rect 21952 45124 21956 45180
rect 21956 45124 22012 45180
rect 22012 45124 22016 45180
rect 21952 45120 22016 45124
rect 22032 45180 22096 45184
rect 22032 45124 22036 45180
rect 22036 45124 22092 45180
rect 22092 45124 22096 45180
rect 22032 45120 22096 45124
rect 22112 45180 22176 45184
rect 22112 45124 22116 45180
rect 22116 45124 22172 45180
rect 22172 45124 22176 45180
rect 22112 45120 22176 45124
rect 22192 45180 22256 45184
rect 22192 45124 22196 45180
rect 22196 45124 22252 45180
rect 22252 45124 22256 45180
rect 22192 45120 22256 45124
rect 26952 45180 27016 45184
rect 26952 45124 26956 45180
rect 26956 45124 27012 45180
rect 27012 45124 27016 45180
rect 26952 45120 27016 45124
rect 27032 45180 27096 45184
rect 27032 45124 27036 45180
rect 27036 45124 27092 45180
rect 27092 45124 27096 45180
rect 27032 45120 27096 45124
rect 27112 45180 27176 45184
rect 27112 45124 27116 45180
rect 27116 45124 27172 45180
rect 27172 45124 27176 45180
rect 27112 45120 27176 45124
rect 27192 45180 27256 45184
rect 27192 45124 27196 45180
rect 27196 45124 27252 45180
rect 27252 45124 27256 45180
rect 27192 45120 27256 45124
rect 31952 45180 32016 45184
rect 31952 45124 31956 45180
rect 31956 45124 32012 45180
rect 32012 45124 32016 45180
rect 31952 45120 32016 45124
rect 32032 45180 32096 45184
rect 32032 45124 32036 45180
rect 32036 45124 32092 45180
rect 32092 45124 32096 45180
rect 32032 45120 32096 45124
rect 32112 45180 32176 45184
rect 32112 45124 32116 45180
rect 32116 45124 32172 45180
rect 32172 45124 32176 45180
rect 32112 45120 32176 45124
rect 32192 45180 32256 45184
rect 32192 45124 32196 45180
rect 32196 45124 32252 45180
rect 32252 45124 32256 45180
rect 32192 45120 32256 45124
rect 36952 45180 37016 45184
rect 36952 45124 36956 45180
rect 36956 45124 37012 45180
rect 37012 45124 37016 45180
rect 36952 45120 37016 45124
rect 37032 45180 37096 45184
rect 37032 45124 37036 45180
rect 37036 45124 37092 45180
rect 37092 45124 37096 45180
rect 37032 45120 37096 45124
rect 37112 45180 37176 45184
rect 37112 45124 37116 45180
rect 37116 45124 37172 45180
rect 37172 45124 37176 45180
rect 37112 45120 37176 45124
rect 37192 45180 37256 45184
rect 37192 45124 37196 45180
rect 37196 45124 37252 45180
rect 37252 45124 37256 45180
rect 37192 45120 37256 45124
rect 41952 45180 42016 45184
rect 41952 45124 41956 45180
rect 41956 45124 42012 45180
rect 42012 45124 42016 45180
rect 41952 45120 42016 45124
rect 42032 45180 42096 45184
rect 42032 45124 42036 45180
rect 42036 45124 42092 45180
rect 42092 45124 42096 45180
rect 42032 45120 42096 45124
rect 42112 45180 42176 45184
rect 42112 45124 42116 45180
rect 42116 45124 42172 45180
rect 42172 45124 42176 45180
rect 42112 45120 42176 45124
rect 42192 45180 42256 45184
rect 42192 45124 42196 45180
rect 42196 45124 42252 45180
rect 42252 45124 42256 45180
rect 42192 45120 42256 45124
rect 46952 45180 47016 45184
rect 46952 45124 46956 45180
rect 46956 45124 47012 45180
rect 47012 45124 47016 45180
rect 46952 45120 47016 45124
rect 47032 45180 47096 45184
rect 47032 45124 47036 45180
rect 47036 45124 47092 45180
rect 47092 45124 47096 45180
rect 47032 45120 47096 45124
rect 47112 45180 47176 45184
rect 47112 45124 47116 45180
rect 47116 45124 47172 45180
rect 47172 45124 47176 45180
rect 47112 45120 47176 45124
rect 47192 45180 47256 45184
rect 47192 45124 47196 45180
rect 47196 45124 47252 45180
rect 47252 45124 47256 45180
rect 47192 45120 47256 45124
rect 51952 45180 52016 45184
rect 51952 45124 51956 45180
rect 51956 45124 52012 45180
rect 52012 45124 52016 45180
rect 51952 45120 52016 45124
rect 52032 45180 52096 45184
rect 52032 45124 52036 45180
rect 52036 45124 52092 45180
rect 52092 45124 52096 45180
rect 52032 45120 52096 45124
rect 52112 45180 52176 45184
rect 52112 45124 52116 45180
rect 52116 45124 52172 45180
rect 52172 45124 52176 45180
rect 52112 45120 52176 45124
rect 52192 45180 52256 45184
rect 52192 45124 52196 45180
rect 52196 45124 52252 45180
rect 52252 45124 52256 45180
rect 52192 45120 52256 45124
rect 56952 45180 57016 45184
rect 56952 45124 56956 45180
rect 56956 45124 57012 45180
rect 57012 45124 57016 45180
rect 56952 45120 57016 45124
rect 57032 45180 57096 45184
rect 57032 45124 57036 45180
rect 57036 45124 57092 45180
rect 57092 45124 57096 45180
rect 57032 45120 57096 45124
rect 57112 45180 57176 45184
rect 57112 45124 57116 45180
rect 57116 45124 57172 45180
rect 57172 45124 57176 45180
rect 57112 45120 57176 45124
rect 57192 45180 57256 45184
rect 57192 45124 57196 45180
rect 57196 45124 57252 45180
rect 57252 45124 57256 45180
rect 57192 45120 57256 45124
rect 2612 44636 2676 44640
rect 2612 44580 2616 44636
rect 2616 44580 2672 44636
rect 2672 44580 2676 44636
rect 2612 44576 2676 44580
rect 2692 44636 2756 44640
rect 2692 44580 2696 44636
rect 2696 44580 2752 44636
rect 2752 44580 2756 44636
rect 2692 44576 2756 44580
rect 2772 44636 2836 44640
rect 2772 44580 2776 44636
rect 2776 44580 2832 44636
rect 2832 44580 2836 44636
rect 2772 44576 2836 44580
rect 2852 44636 2916 44640
rect 2852 44580 2856 44636
rect 2856 44580 2912 44636
rect 2912 44580 2916 44636
rect 2852 44576 2916 44580
rect 7612 44636 7676 44640
rect 7612 44580 7616 44636
rect 7616 44580 7672 44636
rect 7672 44580 7676 44636
rect 7612 44576 7676 44580
rect 7692 44636 7756 44640
rect 7692 44580 7696 44636
rect 7696 44580 7752 44636
rect 7752 44580 7756 44636
rect 7692 44576 7756 44580
rect 7772 44636 7836 44640
rect 7772 44580 7776 44636
rect 7776 44580 7832 44636
rect 7832 44580 7836 44636
rect 7772 44576 7836 44580
rect 7852 44636 7916 44640
rect 7852 44580 7856 44636
rect 7856 44580 7912 44636
rect 7912 44580 7916 44636
rect 7852 44576 7916 44580
rect 12612 44636 12676 44640
rect 12612 44580 12616 44636
rect 12616 44580 12672 44636
rect 12672 44580 12676 44636
rect 12612 44576 12676 44580
rect 12692 44636 12756 44640
rect 12692 44580 12696 44636
rect 12696 44580 12752 44636
rect 12752 44580 12756 44636
rect 12692 44576 12756 44580
rect 12772 44636 12836 44640
rect 12772 44580 12776 44636
rect 12776 44580 12832 44636
rect 12832 44580 12836 44636
rect 12772 44576 12836 44580
rect 12852 44636 12916 44640
rect 12852 44580 12856 44636
rect 12856 44580 12912 44636
rect 12912 44580 12916 44636
rect 12852 44576 12916 44580
rect 17612 44636 17676 44640
rect 17612 44580 17616 44636
rect 17616 44580 17672 44636
rect 17672 44580 17676 44636
rect 17612 44576 17676 44580
rect 17692 44636 17756 44640
rect 17692 44580 17696 44636
rect 17696 44580 17752 44636
rect 17752 44580 17756 44636
rect 17692 44576 17756 44580
rect 17772 44636 17836 44640
rect 17772 44580 17776 44636
rect 17776 44580 17832 44636
rect 17832 44580 17836 44636
rect 17772 44576 17836 44580
rect 17852 44636 17916 44640
rect 17852 44580 17856 44636
rect 17856 44580 17912 44636
rect 17912 44580 17916 44636
rect 17852 44576 17916 44580
rect 22612 44636 22676 44640
rect 22612 44580 22616 44636
rect 22616 44580 22672 44636
rect 22672 44580 22676 44636
rect 22612 44576 22676 44580
rect 22692 44636 22756 44640
rect 22692 44580 22696 44636
rect 22696 44580 22752 44636
rect 22752 44580 22756 44636
rect 22692 44576 22756 44580
rect 22772 44636 22836 44640
rect 22772 44580 22776 44636
rect 22776 44580 22832 44636
rect 22832 44580 22836 44636
rect 22772 44576 22836 44580
rect 22852 44636 22916 44640
rect 22852 44580 22856 44636
rect 22856 44580 22912 44636
rect 22912 44580 22916 44636
rect 22852 44576 22916 44580
rect 27612 44636 27676 44640
rect 27612 44580 27616 44636
rect 27616 44580 27672 44636
rect 27672 44580 27676 44636
rect 27612 44576 27676 44580
rect 27692 44636 27756 44640
rect 27692 44580 27696 44636
rect 27696 44580 27752 44636
rect 27752 44580 27756 44636
rect 27692 44576 27756 44580
rect 27772 44636 27836 44640
rect 27772 44580 27776 44636
rect 27776 44580 27832 44636
rect 27832 44580 27836 44636
rect 27772 44576 27836 44580
rect 27852 44636 27916 44640
rect 27852 44580 27856 44636
rect 27856 44580 27912 44636
rect 27912 44580 27916 44636
rect 27852 44576 27916 44580
rect 32612 44636 32676 44640
rect 32612 44580 32616 44636
rect 32616 44580 32672 44636
rect 32672 44580 32676 44636
rect 32612 44576 32676 44580
rect 32692 44636 32756 44640
rect 32692 44580 32696 44636
rect 32696 44580 32752 44636
rect 32752 44580 32756 44636
rect 32692 44576 32756 44580
rect 32772 44636 32836 44640
rect 32772 44580 32776 44636
rect 32776 44580 32832 44636
rect 32832 44580 32836 44636
rect 32772 44576 32836 44580
rect 32852 44636 32916 44640
rect 32852 44580 32856 44636
rect 32856 44580 32912 44636
rect 32912 44580 32916 44636
rect 32852 44576 32916 44580
rect 37612 44636 37676 44640
rect 37612 44580 37616 44636
rect 37616 44580 37672 44636
rect 37672 44580 37676 44636
rect 37612 44576 37676 44580
rect 37692 44636 37756 44640
rect 37692 44580 37696 44636
rect 37696 44580 37752 44636
rect 37752 44580 37756 44636
rect 37692 44576 37756 44580
rect 37772 44636 37836 44640
rect 37772 44580 37776 44636
rect 37776 44580 37832 44636
rect 37832 44580 37836 44636
rect 37772 44576 37836 44580
rect 37852 44636 37916 44640
rect 37852 44580 37856 44636
rect 37856 44580 37912 44636
rect 37912 44580 37916 44636
rect 37852 44576 37916 44580
rect 42612 44636 42676 44640
rect 42612 44580 42616 44636
rect 42616 44580 42672 44636
rect 42672 44580 42676 44636
rect 42612 44576 42676 44580
rect 42692 44636 42756 44640
rect 42692 44580 42696 44636
rect 42696 44580 42752 44636
rect 42752 44580 42756 44636
rect 42692 44576 42756 44580
rect 42772 44636 42836 44640
rect 42772 44580 42776 44636
rect 42776 44580 42832 44636
rect 42832 44580 42836 44636
rect 42772 44576 42836 44580
rect 42852 44636 42916 44640
rect 42852 44580 42856 44636
rect 42856 44580 42912 44636
rect 42912 44580 42916 44636
rect 42852 44576 42916 44580
rect 47612 44636 47676 44640
rect 47612 44580 47616 44636
rect 47616 44580 47672 44636
rect 47672 44580 47676 44636
rect 47612 44576 47676 44580
rect 47692 44636 47756 44640
rect 47692 44580 47696 44636
rect 47696 44580 47752 44636
rect 47752 44580 47756 44636
rect 47692 44576 47756 44580
rect 47772 44636 47836 44640
rect 47772 44580 47776 44636
rect 47776 44580 47832 44636
rect 47832 44580 47836 44636
rect 47772 44576 47836 44580
rect 47852 44636 47916 44640
rect 47852 44580 47856 44636
rect 47856 44580 47912 44636
rect 47912 44580 47916 44636
rect 47852 44576 47916 44580
rect 52612 44636 52676 44640
rect 52612 44580 52616 44636
rect 52616 44580 52672 44636
rect 52672 44580 52676 44636
rect 52612 44576 52676 44580
rect 52692 44636 52756 44640
rect 52692 44580 52696 44636
rect 52696 44580 52752 44636
rect 52752 44580 52756 44636
rect 52692 44576 52756 44580
rect 52772 44636 52836 44640
rect 52772 44580 52776 44636
rect 52776 44580 52832 44636
rect 52832 44580 52836 44636
rect 52772 44576 52836 44580
rect 52852 44636 52916 44640
rect 52852 44580 52856 44636
rect 52856 44580 52912 44636
rect 52912 44580 52916 44636
rect 52852 44576 52916 44580
rect 57612 44636 57676 44640
rect 57612 44580 57616 44636
rect 57616 44580 57672 44636
rect 57672 44580 57676 44636
rect 57612 44576 57676 44580
rect 57692 44636 57756 44640
rect 57692 44580 57696 44636
rect 57696 44580 57752 44636
rect 57752 44580 57756 44636
rect 57692 44576 57756 44580
rect 57772 44636 57836 44640
rect 57772 44580 57776 44636
rect 57776 44580 57832 44636
rect 57832 44580 57836 44636
rect 57772 44576 57836 44580
rect 57852 44636 57916 44640
rect 57852 44580 57856 44636
rect 57856 44580 57912 44636
rect 57912 44580 57916 44636
rect 57852 44576 57916 44580
rect 1952 44092 2016 44096
rect 1952 44036 1956 44092
rect 1956 44036 2012 44092
rect 2012 44036 2016 44092
rect 1952 44032 2016 44036
rect 2032 44092 2096 44096
rect 2032 44036 2036 44092
rect 2036 44036 2092 44092
rect 2092 44036 2096 44092
rect 2032 44032 2096 44036
rect 2112 44092 2176 44096
rect 2112 44036 2116 44092
rect 2116 44036 2172 44092
rect 2172 44036 2176 44092
rect 2112 44032 2176 44036
rect 2192 44092 2256 44096
rect 2192 44036 2196 44092
rect 2196 44036 2252 44092
rect 2252 44036 2256 44092
rect 2192 44032 2256 44036
rect 6952 44092 7016 44096
rect 6952 44036 6956 44092
rect 6956 44036 7012 44092
rect 7012 44036 7016 44092
rect 6952 44032 7016 44036
rect 7032 44092 7096 44096
rect 7032 44036 7036 44092
rect 7036 44036 7092 44092
rect 7092 44036 7096 44092
rect 7032 44032 7096 44036
rect 7112 44092 7176 44096
rect 7112 44036 7116 44092
rect 7116 44036 7172 44092
rect 7172 44036 7176 44092
rect 7112 44032 7176 44036
rect 7192 44092 7256 44096
rect 7192 44036 7196 44092
rect 7196 44036 7252 44092
rect 7252 44036 7256 44092
rect 7192 44032 7256 44036
rect 11952 44092 12016 44096
rect 11952 44036 11956 44092
rect 11956 44036 12012 44092
rect 12012 44036 12016 44092
rect 11952 44032 12016 44036
rect 12032 44092 12096 44096
rect 12032 44036 12036 44092
rect 12036 44036 12092 44092
rect 12092 44036 12096 44092
rect 12032 44032 12096 44036
rect 12112 44092 12176 44096
rect 12112 44036 12116 44092
rect 12116 44036 12172 44092
rect 12172 44036 12176 44092
rect 12112 44032 12176 44036
rect 12192 44092 12256 44096
rect 12192 44036 12196 44092
rect 12196 44036 12252 44092
rect 12252 44036 12256 44092
rect 12192 44032 12256 44036
rect 16952 44092 17016 44096
rect 16952 44036 16956 44092
rect 16956 44036 17012 44092
rect 17012 44036 17016 44092
rect 16952 44032 17016 44036
rect 17032 44092 17096 44096
rect 17032 44036 17036 44092
rect 17036 44036 17092 44092
rect 17092 44036 17096 44092
rect 17032 44032 17096 44036
rect 17112 44092 17176 44096
rect 17112 44036 17116 44092
rect 17116 44036 17172 44092
rect 17172 44036 17176 44092
rect 17112 44032 17176 44036
rect 17192 44092 17256 44096
rect 17192 44036 17196 44092
rect 17196 44036 17252 44092
rect 17252 44036 17256 44092
rect 17192 44032 17256 44036
rect 21952 44092 22016 44096
rect 21952 44036 21956 44092
rect 21956 44036 22012 44092
rect 22012 44036 22016 44092
rect 21952 44032 22016 44036
rect 22032 44092 22096 44096
rect 22032 44036 22036 44092
rect 22036 44036 22092 44092
rect 22092 44036 22096 44092
rect 22032 44032 22096 44036
rect 22112 44092 22176 44096
rect 22112 44036 22116 44092
rect 22116 44036 22172 44092
rect 22172 44036 22176 44092
rect 22112 44032 22176 44036
rect 22192 44092 22256 44096
rect 22192 44036 22196 44092
rect 22196 44036 22252 44092
rect 22252 44036 22256 44092
rect 22192 44032 22256 44036
rect 26952 44092 27016 44096
rect 26952 44036 26956 44092
rect 26956 44036 27012 44092
rect 27012 44036 27016 44092
rect 26952 44032 27016 44036
rect 27032 44092 27096 44096
rect 27032 44036 27036 44092
rect 27036 44036 27092 44092
rect 27092 44036 27096 44092
rect 27032 44032 27096 44036
rect 27112 44092 27176 44096
rect 27112 44036 27116 44092
rect 27116 44036 27172 44092
rect 27172 44036 27176 44092
rect 27112 44032 27176 44036
rect 27192 44092 27256 44096
rect 27192 44036 27196 44092
rect 27196 44036 27252 44092
rect 27252 44036 27256 44092
rect 27192 44032 27256 44036
rect 31952 44092 32016 44096
rect 31952 44036 31956 44092
rect 31956 44036 32012 44092
rect 32012 44036 32016 44092
rect 31952 44032 32016 44036
rect 32032 44092 32096 44096
rect 32032 44036 32036 44092
rect 32036 44036 32092 44092
rect 32092 44036 32096 44092
rect 32032 44032 32096 44036
rect 32112 44092 32176 44096
rect 32112 44036 32116 44092
rect 32116 44036 32172 44092
rect 32172 44036 32176 44092
rect 32112 44032 32176 44036
rect 32192 44092 32256 44096
rect 32192 44036 32196 44092
rect 32196 44036 32252 44092
rect 32252 44036 32256 44092
rect 32192 44032 32256 44036
rect 36952 44092 37016 44096
rect 36952 44036 36956 44092
rect 36956 44036 37012 44092
rect 37012 44036 37016 44092
rect 36952 44032 37016 44036
rect 37032 44092 37096 44096
rect 37032 44036 37036 44092
rect 37036 44036 37092 44092
rect 37092 44036 37096 44092
rect 37032 44032 37096 44036
rect 37112 44092 37176 44096
rect 37112 44036 37116 44092
rect 37116 44036 37172 44092
rect 37172 44036 37176 44092
rect 37112 44032 37176 44036
rect 37192 44092 37256 44096
rect 37192 44036 37196 44092
rect 37196 44036 37252 44092
rect 37252 44036 37256 44092
rect 37192 44032 37256 44036
rect 41952 44092 42016 44096
rect 41952 44036 41956 44092
rect 41956 44036 42012 44092
rect 42012 44036 42016 44092
rect 41952 44032 42016 44036
rect 42032 44092 42096 44096
rect 42032 44036 42036 44092
rect 42036 44036 42092 44092
rect 42092 44036 42096 44092
rect 42032 44032 42096 44036
rect 42112 44092 42176 44096
rect 42112 44036 42116 44092
rect 42116 44036 42172 44092
rect 42172 44036 42176 44092
rect 42112 44032 42176 44036
rect 42192 44092 42256 44096
rect 42192 44036 42196 44092
rect 42196 44036 42252 44092
rect 42252 44036 42256 44092
rect 42192 44032 42256 44036
rect 46952 44092 47016 44096
rect 46952 44036 46956 44092
rect 46956 44036 47012 44092
rect 47012 44036 47016 44092
rect 46952 44032 47016 44036
rect 47032 44092 47096 44096
rect 47032 44036 47036 44092
rect 47036 44036 47092 44092
rect 47092 44036 47096 44092
rect 47032 44032 47096 44036
rect 47112 44092 47176 44096
rect 47112 44036 47116 44092
rect 47116 44036 47172 44092
rect 47172 44036 47176 44092
rect 47112 44032 47176 44036
rect 47192 44092 47256 44096
rect 47192 44036 47196 44092
rect 47196 44036 47252 44092
rect 47252 44036 47256 44092
rect 47192 44032 47256 44036
rect 51952 44092 52016 44096
rect 51952 44036 51956 44092
rect 51956 44036 52012 44092
rect 52012 44036 52016 44092
rect 51952 44032 52016 44036
rect 52032 44092 52096 44096
rect 52032 44036 52036 44092
rect 52036 44036 52092 44092
rect 52092 44036 52096 44092
rect 52032 44032 52096 44036
rect 52112 44092 52176 44096
rect 52112 44036 52116 44092
rect 52116 44036 52172 44092
rect 52172 44036 52176 44092
rect 52112 44032 52176 44036
rect 52192 44092 52256 44096
rect 52192 44036 52196 44092
rect 52196 44036 52252 44092
rect 52252 44036 52256 44092
rect 52192 44032 52256 44036
rect 56952 44092 57016 44096
rect 56952 44036 56956 44092
rect 56956 44036 57012 44092
rect 57012 44036 57016 44092
rect 56952 44032 57016 44036
rect 57032 44092 57096 44096
rect 57032 44036 57036 44092
rect 57036 44036 57092 44092
rect 57092 44036 57096 44092
rect 57032 44032 57096 44036
rect 57112 44092 57176 44096
rect 57112 44036 57116 44092
rect 57116 44036 57172 44092
rect 57172 44036 57176 44092
rect 57112 44032 57176 44036
rect 57192 44092 57256 44096
rect 57192 44036 57196 44092
rect 57196 44036 57252 44092
rect 57252 44036 57256 44092
rect 57192 44032 57256 44036
rect 2612 43548 2676 43552
rect 2612 43492 2616 43548
rect 2616 43492 2672 43548
rect 2672 43492 2676 43548
rect 2612 43488 2676 43492
rect 2692 43548 2756 43552
rect 2692 43492 2696 43548
rect 2696 43492 2752 43548
rect 2752 43492 2756 43548
rect 2692 43488 2756 43492
rect 2772 43548 2836 43552
rect 2772 43492 2776 43548
rect 2776 43492 2832 43548
rect 2832 43492 2836 43548
rect 2772 43488 2836 43492
rect 2852 43548 2916 43552
rect 2852 43492 2856 43548
rect 2856 43492 2912 43548
rect 2912 43492 2916 43548
rect 2852 43488 2916 43492
rect 7612 43548 7676 43552
rect 7612 43492 7616 43548
rect 7616 43492 7672 43548
rect 7672 43492 7676 43548
rect 7612 43488 7676 43492
rect 7692 43548 7756 43552
rect 7692 43492 7696 43548
rect 7696 43492 7752 43548
rect 7752 43492 7756 43548
rect 7692 43488 7756 43492
rect 7772 43548 7836 43552
rect 7772 43492 7776 43548
rect 7776 43492 7832 43548
rect 7832 43492 7836 43548
rect 7772 43488 7836 43492
rect 7852 43548 7916 43552
rect 7852 43492 7856 43548
rect 7856 43492 7912 43548
rect 7912 43492 7916 43548
rect 7852 43488 7916 43492
rect 12612 43548 12676 43552
rect 12612 43492 12616 43548
rect 12616 43492 12672 43548
rect 12672 43492 12676 43548
rect 12612 43488 12676 43492
rect 12692 43548 12756 43552
rect 12692 43492 12696 43548
rect 12696 43492 12752 43548
rect 12752 43492 12756 43548
rect 12692 43488 12756 43492
rect 12772 43548 12836 43552
rect 12772 43492 12776 43548
rect 12776 43492 12832 43548
rect 12832 43492 12836 43548
rect 12772 43488 12836 43492
rect 12852 43548 12916 43552
rect 12852 43492 12856 43548
rect 12856 43492 12912 43548
rect 12912 43492 12916 43548
rect 12852 43488 12916 43492
rect 17612 43548 17676 43552
rect 17612 43492 17616 43548
rect 17616 43492 17672 43548
rect 17672 43492 17676 43548
rect 17612 43488 17676 43492
rect 17692 43548 17756 43552
rect 17692 43492 17696 43548
rect 17696 43492 17752 43548
rect 17752 43492 17756 43548
rect 17692 43488 17756 43492
rect 17772 43548 17836 43552
rect 17772 43492 17776 43548
rect 17776 43492 17832 43548
rect 17832 43492 17836 43548
rect 17772 43488 17836 43492
rect 17852 43548 17916 43552
rect 17852 43492 17856 43548
rect 17856 43492 17912 43548
rect 17912 43492 17916 43548
rect 17852 43488 17916 43492
rect 22612 43548 22676 43552
rect 22612 43492 22616 43548
rect 22616 43492 22672 43548
rect 22672 43492 22676 43548
rect 22612 43488 22676 43492
rect 22692 43548 22756 43552
rect 22692 43492 22696 43548
rect 22696 43492 22752 43548
rect 22752 43492 22756 43548
rect 22692 43488 22756 43492
rect 22772 43548 22836 43552
rect 22772 43492 22776 43548
rect 22776 43492 22832 43548
rect 22832 43492 22836 43548
rect 22772 43488 22836 43492
rect 22852 43548 22916 43552
rect 22852 43492 22856 43548
rect 22856 43492 22912 43548
rect 22912 43492 22916 43548
rect 22852 43488 22916 43492
rect 27612 43548 27676 43552
rect 27612 43492 27616 43548
rect 27616 43492 27672 43548
rect 27672 43492 27676 43548
rect 27612 43488 27676 43492
rect 27692 43548 27756 43552
rect 27692 43492 27696 43548
rect 27696 43492 27752 43548
rect 27752 43492 27756 43548
rect 27692 43488 27756 43492
rect 27772 43548 27836 43552
rect 27772 43492 27776 43548
rect 27776 43492 27832 43548
rect 27832 43492 27836 43548
rect 27772 43488 27836 43492
rect 27852 43548 27916 43552
rect 27852 43492 27856 43548
rect 27856 43492 27912 43548
rect 27912 43492 27916 43548
rect 27852 43488 27916 43492
rect 32612 43548 32676 43552
rect 32612 43492 32616 43548
rect 32616 43492 32672 43548
rect 32672 43492 32676 43548
rect 32612 43488 32676 43492
rect 32692 43548 32756 43552
rect 32692 43492 32696 43548
rect 32696 43492 32752 43548
rect 32752 43492 32756 43548
rect 32692 43488 32756 43492
rect 32772 43548 32836 43552
rect 32772 43492 32776 43548
rect 32776 43492 32832 43548
rect 32832 43492 32836 43548
rect 32772 43488 32836 43492
rect 32852 43548 32916 43552
rect 32852 43492 32856 43548
rect 32856 43492 32912 43548
rect 32912 43492 32916 43548
rect 32852 43488 32916 43492
rect 37612 43548 37676 43552
rect 37612 43492 37616 43548
rect 37616 43492 37672 43548
rect 37672 43492 37676 43548
rect 37612 43488 37676 43492
rect 37692 43548 37756 43552
rect 37692 43492 37696 43548
rect 37696 43492 37752 43548
rect 37752 43492 37756 43548
rect 37692 43488 37756 43492
rect 37772 43548 37836 43552
rect 37772 43492 37776 43548
rect 37776 43492 37832 43548
rect 37832 43492 37836 43548
rect 37772 43488 37836 43492
rect 37852 43548 37916 43552
rect 37852 43492 37856 43548
rect 37856 43492 37912 43548
rect 37912 43492 37916 43548
rect 37852 43488 37916 43492
rect 42612 43548 42676 43552
rect 42612 43492 42616 43548
rect 42616 43492 42672 43548
rect 42672 43492 42676 43548
rect 42612 43488 42676 43492
rect 42692 43548 42756 43552
rect 42692 43492 42696 43548
rect 42696 43492 42752 43548
rect 42752 43492 42756 43548
rect 42692 43488 42756 43492
rect 42772 43548 42836 43552
rect 42772 43492 42776 43548
rect 42776 43492 42832 43548
rect 42832 43492 42836 43548
rect 42772 43488 42836 43492
rect 42852 43548 42916 43552
rect 42852 43492 42856 43548
rect 42856 43492 42912 43548
rect 42912 43492 42916 43548
rect 42852 43488 42916 43492
rect 47612 43548 47676 43552
rect 47612 43492 47616 43548
rect 47616 43492 47672 43548
rect 47672 43492 47676 43548
rect 47612 43488 47676 43492
rect 47692 43548 47756 43552
rect 47692 43492 47696 43548
rect 47696 43492 47752 43548
rect 47752 43492 47756 43548
rect 47692 43488 47756 43492
rect 47772 43548 47836 43552
rect 47772 43492 47776 43548
rect 47776 43492 47832 43548
rect 47832 43492 47836 43548
rect 47772 43488 47836 43492
rect 47852 43548 47916 43552
rect 47852 43492 47856 43548
rect 47856 43492 47912 43548
rect 47912 43492 47916 43548
rect 47852 43488 47916 43492
rect 52612 43548 52676 43552
rect 52612 43492 52616 43548
rect 52616 43492 52672 43548
rect 52672 43492 52676 43548
rect 52612 43488 52676 43492
rect 52692 43548 52756 43552
rect 52692 43492 52696 43548
rect 52696 43492 52752 43548
rect 52752 43492 52756 43548
rect 52692 43488 52756 43492
rect 52772 43548 52836 43552
rect 52772 43492 52776 43548
rect 52776 43492 52832 43548
rect 52832 43492 52836 43548
rect 52772 43488 52836 43492
rect 52852 43548 52916 43552
rect 52852 43492 52856 43548
rect 52856 43492 52912 43548
rect 52912 43492 52916 43548
rect 52852 43488 52916 43492
rect 57612 43548 57676 43552
rect 57612 43492 57616 43548
rect 57616 43492 57672 43548
rect 57672 43492 57676 43548
rect 57612 43488 57676 43492
rect 57692 43548 57756 43552
rect 57692 43492 57696 43548
rect 57696 43492 57752 43548
rect 57752 43492 57756 43548
rect 57692 43488 57756 43492
rect 57772 43548 57836 43552
rect 57772 43492 57776 43548
rect 57776 43492 57832 43548
rect 57832 43492 57836 43548
rect 57772 43488 57836 43492
rect 57852 43548 57916 43552
rect 57852 43492 57856 43548
rect 57856 43492 57912 43548
rect 57912 43492 57916 43548
rect 57852 43488 57916 43492
rect 1952 43004 2016 43008
rect 1952 42948 1956 43004
rect 1956 42948 2012 43004
rect 2012 42948 2016 43004
rect 1952 42944 2016 42948
rect 2032 43004 2096 43008
rect 2032 42948 2036 43004
rect 2036 42948 2092 43004
rect 2092 42948 2096 43004
rect 2032 42944 2096 42948
rect 2112 43004 2176 43008
rect 2112 42948 2116 43004
rect 2116 42948 2172 43004
rect 2172 42948 2176 43004
rect 2112 42944 2176 42948
rect 2192 43004 2256 43008
rect 2192 42948 2196 43004
rect 2196 42948 2252 43004
rect 2252 42948 2256 43004
rect 2192 42944 2256 42948
rect 6952 43004 7016 43008
rect 6952 42948 6956 43004
rect 6956 42948 7012 43004
rect 7012 42948 7016 43004
rect 6952 42944 7016 42948
rect 7032 43004 7096 43008
rect 7032 42948 7036 43004
rect 7036 42948 7092 43004
rect 7092 42948 7096 43004
rect 7032 42944 7096 42948
rect 7112 43004 7176 43008
rect 7112 42948 7116 43004
rect 7116 42948 7172 43004
rect 7172 42948 7176 43004
rect 7112 42944 7176 42948
rect 7192 43004 7256 43008
rect 7192 42948 7196 43004
rect 7196 42948 7252 43004
rect 7252 42948 7256 43004
rect 7192 42944 7256 42948
rect 11952 43004 12016 43008
rect 11952 42948 11956 43004
rect 11956 42948 12012 43004
rect 12012 42948 12016 43004
rect 11952 42944 12016 42948
rect 12032 43004 12096 43008
rect 12032 42948 12036 43004
rect 12036 42948 12092 43004
rect 12092 42948 12096 43004
rect 12032 42944 12096 42948
rect 12112 43004 12176 43008
rect 12112 42948 12116 43004
rect 12116 42948 12172 43004
rect 12172 42948 12176 43004
rect 12112 42944 12176 42948
rect 12192 43004 12256 43008
rect 12192 42948 12196 43004
rect 12196 42948 12252 43004
rect 12252 42948 12256 43004
rect 12192 42944 12256 42948
rect 16952 43004 17016 43008
rect 16952 42948 16956 43004
rect 16956 42948 17012 43004
rect 17012 42948 17016 43004
rect 16952 42944 17016 42948
rect 17032 43004 17096 43008
rect 17032 42948 17036 43004
rect 17036 42948 17092 43004
rect 17092 42948 17096 43004
rect 17032 42944 17096 42948
rect 17112 43004 17176 43008
rect 17112 42948 17116 43004
rect 17116 42948 17172 43004
rect 17172 42948 17176 43004
rect 17112 42944 17176 42948
rect 17192 43004 17256 43008
rect 17192 42948 17196 43004
rect 17196 42948 17252 43004
rect 17252 42948 17256 43004
rect 17192 42944 17256 42948
rect 21952 43004 22016 43008
rect 21952 42948 21956 43004
rect 21956 42948 22012 43004
rect 22012 42948 22016 43004
rect 21952 42944 22016 42948
rect 22032 43004 22096 43008
rect 22032 42948 22036 43004
rect 22036 42948 22092 43004
rect 22092 42948 22096 43004
rect 22032 42944 22096 42948
rect 22112 43004 22176 43008
rect 22112 42948 22116 43004
rect 22116 42948 22172 43004
rect 22172 42948 22176 43004
rect 22112 42944 22176 42948
rect 22192 43004 22256 43008
rect 22192 42948 22196 43004
rect 22196 42948 22252 43004
rect 22252 42948 22256 43004
rect 22192 42944 22256 42948
rect 26952 43004 27016 43008
rect 26952 42948 26956 43004
rect 26956 42948 27012 43004
rect 27012 42948 27016 43004
rect 26952 42944 27016 42948
rect 27032 43004 27096 43008
rect 27032 42948 27036 43004
rect 27036 42948 27092 43004
rect 27092 42948 27096 43004
rect 27032 42944 27096 42948
rect 27112 43004 27176 43008
rect 27112 42948 27116 43004
rect 27116 42948 27172 43004
rect 27172 42948 27176 43004
rect 27112 42944 27176 42948
rect 27192 43004 27256 43008
rect 27192 42948 27196 43004
rect 27196 42948 27252 43004
rect 27252 42948 27256 43004
rect 27192 42944 27256 42948
rect 31952 43004 32016 43008
rect 31952 42948 31956 43004
rect 31956 42948 32012 43004
rect 32012 42948 32016 43004
rect 31952 42944 32016 42948
rect 32032 43004 32096 43008
rect 32032 42948 32036 43004
rect 32036 42948 32092 43004
rect 32092 42948 32096 43004
rect 32032 42944 32096 42948
rect 32112 43004 32176 43008
rect 32112 42948 32116 43004
rect 32116 42948 32172 43004
rect 32172 42948 32176 43004
rect 32112 42944 32176 42948
rect 32192 43004 32256 43008
rect 32192 42948 32196 43004
rect 32196 42948 32252 43004
rect 32252 42948 32256 43004
rect 32192 42944 32256 42948
rect 36952 43004 37016 43008
rect 36952 42948 36956 43004
rect 36956 42948 37012 43004
rect 37012 42948 37016 43004
rect 36952 42944 37016 42948
rect 37032 43004 37096 43008
rect 37032 42948 37036 43004
rect 37036 42948 37092 43004
rect 37092 42948 37096 43004
rect 37032 42944 37096 42948
rect 37112 43004 37176 43008
rect 37112 42948 37116 43004
rect 37116 42948 37172 43004
rect 37172 42948 37176 43004
rect 37112 42944 37176 42948
rect 37192 43004 37256 43008
rect 37192 42948 37196 43004
rect 37196 42948 37252 43004
rect 37252 42948 37256 43004
rect 37192 42944 37256 42948
rect 41952 43004 42016 43008
rect 41952 42948 41956 43004
rect 41956 42948 42012 43004
rect 42012 42948 42016 43004
rect 41952 42944 42016 42948
rect 42032 43004 42096 43008
rect 42032 42948 42036 43004
rect 42036 42948 42092 43004
rect 42092 42948 42096 43004
rect 42032 42944 42096 42948
rect 42112 43004 42176 43008
rect 42112 42948 42116 43004
rect 42116 42948 42172 43004
rect 42172 42948 42176 43004
rect 42112 42944 42176 42948
rect 42192 43004 42256 43008
rect 42192 42948 42196 43004
rect 42196 42948 42252 43004
rect 42252 42948 42256 43004
rect 42192 42944 42256 42948
rect 46952 43004 47016 43008
rect 46952 42948 46956 43004
rect 46956 42948 47012 43004
rect 47012 42948 47016 43004
rect 46952 42944 47016 42948
rect 47032 43004 47096 43008
rect 47032 42948 47036 43004
rect 47036 42948 47092 43004
rect 47092 42948 47096 43004
rect 47032 42944 47096 42948
rect 47112 43004 47176 43008
rect 47112 42948 47116 43004
rect 47116 42948 47172 43004
rect 47172 42948 47176 43004
rect 47112 42944 47176 42948
rect 47192 43004 47256 43008
rect 47192 42948 47196 43004
rect 47196 42948 47252 43004
rect 47252 42948 47256 43004
rect 47192 42944 47256 42948
rect 51952 43004 52016 43008
rect 51952 42948 51956 43004
rect 51956 42948 52012 43004
rect 52012 42948 52016 43004
rect 51952 42944 52016 42948
rect 52032 43004 52096 43008
rect 52032 42948 52036 43004
rect 52036 42948 52092 43004
rect 52092 42948 52096 43004
rect 52032 42944 52096 42948
rect 52112 43004 52176 43008
rect 52112 42948 52116 43004
rect 52116 42948 52172 43004
rect 52172 42948 52176 43004
rect 52112 42944 52176 42948
rect 52192 43004 52256 43008
rect 52192 42948 52196 43004
rect 52196 42948 52252 43004
rect 52252 42948 52256 43004
rect 52192 42944 52256 42948
rect 56952 43004 57016 43008
rect 56952 42948 56956 43004
rect 56956 42948 57012 43004
rect 57012 42948 57016 43004
rect 56952 42944 57016 42948
rect 57032 43004 57096 43008
rect 57032 42948 57036 43004
rect 57036 42948 57092 43004
rect 57092 42948 57096 43004
rect 57032 42944 57096 42948
rect 57112 43004 57176 43008
rect 57112 42948 57116 43004
rect 57116 42948 57172 43004
rect 57172 42948 57176 43004
rect 57112 42944 57176 42948
rect 57192 43004 57256 43008
rect 57192 42948 57196 43004
rect 57196 42948 57252 43004
rect 57252 42948 57256 43004
rect 57192 42944 57256 42948
rect 2612 42460 2676 42464
rect 2612 42404 2616 42460
rect 2616 42404 2672 42460
rect 2672 42404 2676 42460
rect 2612 42400 2676 42404
rect 2692 42460 2756 42464
rect 2692 42404 2696 42460
rect 2696 42404 2752 42460
rect 2752 42404 2756 42460
rect 2692 42400 2756 42404
rect 2772 42460 2836 42464
rect 2772 42404 2776 42460
rect 2776 42404 2832 42460
rect 2832 42404 2836 42460
rect 2772 42400 2836 42404
rect 2852 42460 2916 42464
rect 2852 42404 2856 42460
rect 2856 42404 2912 42460
rect 2912 42404 2916 42460
rect 2852 42400 2916 42404
rect 7612 42460 7676 42464
rect 7612 42404 7616 42460
rect 7616 42404 7672 42460
rect 7672 42404 7676 42460
rect 7612 42400 7676 42404
rect 7692 42460 7756 42464
rect 7692 42404 7696 42460
rect 7696 42404 7752 42460
rect 7752 42404 7756 42460
rect 7692 42400 7756 42404
rect 7772 42460 7836 42464
rect 7772 42404 7776 42460
rect 7776 42404 7832 42460
rect 7832 42404 7836 42460
rect 7772 42400 7836 42404
rect 7852 42460 7916 42464
rect 7852 42404 7856 42460
rect 7856 42404 7912 42460
rect 7912 42404 7916 42460
rect 7852 42400 7916 42404
rect 12612 42460 12676 42464
rect 12612 42404 12616 42460
rect 12616 42404 12672 42460
rect 12672 42404 12676 42460
rect 12612 42400 12676 42404
rect 12692 42460 12756 42464
rect 12692 42404 12696 42460
rect 12696 42404 12752 42460
rect 12752 42404 12756 42460
rect 12692 42400 12756 42404
rect 12772 42460 12836 42464
rect 12772 42404 12776 42460
rect 12776 42404 12832 42460
rect 12832 42404 12836 42460
rect 12772 42400 12836 42404
rect 12852 42460 12916 42464
rect 12852 42404 12856 42460
rect 12856 42404 12912 42460
rect 12912 42404 12916 42460
rect 12852 42400 12916 42404
rect 17612 42460 17676 42464
rect 17612 42404 17616 42460
rect 17616 42404 17672 42460
rect 17672 42404 17676 42460
rect 17612 42400 17676 42404
rect 17692 42460 17756 42464
rect 17692 42404 17696 42460
rect 17696 42404 17752 42460
rect 17752 42404 17756 42460
rect 17692 42400 17756 42404
rect 17772 42460 17836 42464
rect 17772 42404 17776 42460
rect 17776 42404 17832 42460
rect 17832 42404 17836 42460
rect 17772 42400 17836 42404
rect 17852 42460 17916 42464
rect 17852 42404 17856 42460
rect 17856 42404 17912 42460
rect 17912 42404 17916 42460
rect 17852 42400 17916 42404
rect 22612 42460 22676 42464
rect 22612 42404 22616 42460
rect 22616 42404 22672 42460
rect 22672 42404 22676 42460
rect 22612 42400 22676 42404
rect 22692 42460 22756 42464
rect 22692 42404 22696 42460
rect 22696 42404 22752 42460
rect 22752 42404 22756 42460
rect 22692 42400 22756 42404
rect 22772 42460 22836 42464
rect 22772 42404 22776 42460
rect 22776 42404 22832 42460
rect 22832 42404 22836 42460
rect 22772 42400 22836 42404
rect 22852 42460 22916 42464
rect 22852 42404 22856 42460
rect 22856 42404 22912 42460
rect 22912 42404 22916 42460
rect 22852 42400 22916 42404
rect 27612 42460 27676 42464
rect 27612 42404 27616 42460
rect 27616 42404 27672 42460
rect 27672 42404 27676 42460
rect 27612 42400 27676 42404
rect 27692 42460 27756 42464
rect 27692 42404 27696 42460
rect 27696 42404 27752 42460
rect 27752 42404 27756 42460
rect 27692 42400 27756 42404
rect 27772 42460 27836 42464
rect 27772 42404 27776 42460
rect 27776 42404 27832 42460
rect 27832 42404 27836 42460
rect 27772 42400 27836 42404
rect 27852 42460 27916 42464
rect 27852 42404 27856 42460
rect 27856 42404 27912 42460
rect 27912 42404 27916 42460
rect 27852 42400 27916 42404
rect 32612 42460 32676 42464
rect 32612 42404 32616 42460
rect 32616 42404 32672 42460
rect 32672 42404 32676 42460
rect 32612 42400 32676 42404
rect 32692 42460 32756 42464
rect 32692 42404 32696 42460
rect 32696 42404 32752 42460
rect 32752 42404 32756 42460
rect 32692 42400 32756 42404
rect 32772 42460 32836 42464
rect 32772 42404 32776 42460
rect 32776 42404 32832 42460
rect 32832 42404 32836 42460
rect 32772 42400 32836 42404
rect 32852 42460 32916 42464
rect 32852 42404 32856 42460
rect 32856 42404 32912 42460
rect 32912 42404 32916 42460
rect 32852 42400 32916 42404
rect 37612 42460 37676 42464
rect 37612 42404 37616 42460
rect 37616 42404 37672 42460
rect 37672 42404 37676 42460
rect 37612 42400 37676 42404
rect 37692 42460 37756 42464
rect 37692 42404 37696 42460
rect 37696 42404 37752 42460
rect 37752 42404 37756 42460
rect 37692 42400 37756 42404
rect 37772 42460 37836 42464
rect 37772 42404 37776 42460
rect 37776 42404 37832 42460
rect 37832 42404 37836 42460
rect 37772 42400 37836 42404
rect 37852 42460 37916 42464
rect 37852 42404 37856 42460
rect 37856 42404 37912 42460
rect 37912 42404 37916 42460
rect 37852 42400 37916 42404
rect 42612 42460 42676 42464
rect 42612 42404 42616 42460
rect 42616 42404 42672 42460
rect 42672 42404 42676 42460
rect 42612 42400 42676 42404
rect 42692 42460 42756 42464
rect 42692 42404 42696 42460
rect 42696 42404 42752 42460
rect 42752 42404 42756 42460
rect 42692 42400 42756 42404
rect 42772 42460 42836 42464
rect 42772 42404 42776 42460
rect 42776 42404 42832 42460
rect 42832 42404 42836 42460
rect 42772 42400 42836 42404
rect 42852 42460 42916 42464
rect 42852 42404 42856 42460
rect 42856 42404 42912 42460
rect 42912 42404 42916 42460
rect 42852 42400 42916 42404
rect 47612 42460 47676 42464
rect 47612 42404 47616 42460
rect 47616 42404 47672 42460
rect 47672 42404 47676 42460
rect 47612 42400 47676 42404
rect 47692 42460 47756 42464
rect 47692 42404 47696 42460
rect 47696 42404 47752 42460
rect 47752 42404 47756 42460
rect 47692 42400 47756 42404
rect 47772 42460 47836 42464
rect 47772 42404 47776 42460
rect 47776 42404 47832 42460
rect 47832 42404 47836 42460
rect 47772 42400 47836 42404
rect 47852 42460 47916 42464
rect 47852 42404 47856 42460
rect 47856 42404 47912 42460
rect 47912 42404 47916 42460
rect 47852 42400 47916 42404
rect 52612 42460 52676 42464
rect 52612 42404 52616 42460
rect 52616 42404 52672 42460
rect 52672 42404 52676 42460
rect 52612 42400 52676 42404
rect 52692 42460 52756 42464
rect 52692 42404 52696 42460
rect 52696 42404 52752 42460
rect 52752 42404 52756 42460
rect 52692 42400 52756 42404
rect 52772 42460 52836 42464
rect 52772 42404 52776 42460
rect 52776 42404 52832 42460
rect 52832 42404 52836 42460
rect 52772 42400 52836 42404
rect 52852 42460 52916 42464
rect 52852 42404 52856 42460
rect 52856 42404 52912 42460
rect 52912 42404 52916 42460
rect 52852 42400 52916 42404
rect 57612 42460 57676 42464
rect 57612 42404 57616 42460
rect 57616 42404 57672 42460
rect 57672 42404 57676 42460
rect 57612 42400 57676 42404
rect 57692 42460 57756 42464
rect 57692 42404 57696 42460
rect 57696 42404 57752 42460
rect 57752 42404 57756 42460
rect 57692 42400 57756 42404
rect 57772 42460 57836 42464
rect 57772 42404 57776 42460
rect 57776 42404 57832 42460
rect 57832 42404 57836 42460
rect 57772 42400 57836 42404
rect 57852 42460 57916 42464
rect 57852 42404 57856 42460
rect 57856 42404 57912 42460
rect 57912 42404 57916 42460
rect 57852 42400 57916 42404
rect 1952 41916 2016 41920
rect 1952 41860 1956 41916
rect 1956 41860 2012 41916
rect 2012 41860 2016 41916
rect 1952 41856 2016 41860
rect 2032 41916 2096 41920
rect 2032 41860 2036 41916
rect 2036 41860 2092 41916
rect 2092 41860 2096 41916
rect 2032 41856 2096 41860
rect 2112 41916 2176 41920
rect 2112 41860 2116 41916
rect 2116 41860 2172 41916
rect 2172 41860 2176 41916
rect 2112 41856 2176 41860
rect 2192 41916 2256 41920
rect 2192 41860 2196 41916
rect 2196 41860 2252 41916
rect 2252 41860 2256 41916
rect 2192 41856 2256 41860
rect 6952 41916 7016 41920
rect 6952 41860 6956 41916
rect 6956 41860 7012 41916
rect 7012 41860 7016 41916
rect 6952 41856 7016 41860
rect 7032 41916 7096 41920
rect 7032 41860 7036 41916
rect 7036 41860 7092 41916
rect 7092 41860 7096 41916
rect 7032 41856 7096 41860
rect 7112 41916 7176 41920
rect 7112 41860 7116 41916
rect 7116 41860 7172 41916
rect 7172 41860 7176 41916
rect 7112 41856 7176 41860
rect 7192 41916 7256 41920
rect 7192 41860 7196 41916
rect 7196 41860 7252 41916
rect 7252 41860 7256 41916
rect 7192 41856 7256 41860
rect 11952 41916 12016 41920
rect 11952 41860 11956 41916
rect 11956 41860 12012 41916
rect 12012 41860 12016 41916
rect 11952 41856 12016 41860
rect 12032 41916 12096 41920
rect 12032 41860 12036 41916
rect 12036 41860 12092 41916
rect 12092 41860 12096 41916
rect 12032 41856 12096 41860
rect 12112 41916 12176 41920
rect 12112 41860 12116 41916
rect 12116 41860 12172 41916
rect 12172 41860 12176 41916
rect 12112 41856 12176 41860
rect 12192 41916 12256 41920
rect 12192 41860 12196 41916
rect 12196 41860 12252 41916
rect 12252 41860 12256 41916
rect 12192 41856 12256 41860
rect 16952 41916 17016 41920
rect 16952 41860 16956 41916
rect 16956 41860 17012 41916
rect 17012 41860 17016 41916
rect 16952 41856 17016 41860
rect 17032 41916 17096 41920
rect 17032 41860 17036 41916
rect 17036 41860 17092 41916
rect 17092 41860 17096 41916
rect 17032 41856 17096 41860
rect 17112 41916 17176 41920
rect 17112 41860 17116 41916
rect 17116 41860 17172 41916
rect 17172 41860 17176 41916
rect 17112 41856 17176 41860
rect 17192 41916 17256 41920
rect 17192 41860 17196 41916
rect 17196 41860 17252 41916
rect 17252 41860 17256 41916
rect 17192 41856 17256 41860
rect 21952 41916 22016 41920
rect 21952 41860 21956 41916
rect 21956 41860 22012 41916
rect 22012 41860 22016 41916
rect 21952 41856 22016 41860
rect 22032 41916 22096 41920
rect 22032 41860 22036 41916
rect 22036 41860 22092 41916
rect 22092 41860 22096 41916
rect 22032 41856 22096 41860
rect 22112 41916 22176 41920
rect 22112 41860 22116 41916
rect 22116 41860 22172 41916
rect 22172 41860 22176 41916
rect 22112 41856 22176 41860
rect 22192 41916 22256 41920
rect 22192 41860 22196 41916
rect 22196 41860 22252 41916
rect 22252 41860 22256 41916
rect 22192 41856 22256 41860
rect 26952 41916 27016 41920
rect 26952 41860 26956 41916
rect 26956 41860 27012 41916
rect 27012 41860 27016 41916
rect 26952 41856 27016 41860
rect 27032 41916 27096 41920
rect 27032 41860 27036 41916
rect 27036 41860 27092 41916
rect 27092 41860 27096 41916
rect 27032 41856 27096 41860
rect 27112 41916 27176 41920
rect 27112 41860 27116 41916
rect 27116 41860 27172 41916
rect 27172 41860 27176 41916
rect 27112 41856 27176 41860
rect 27192 41916 27256 41920
rect 27192 41860 27196 41916
rect 27196 41860 27252 41916
rect 27252 41860 27256 41916
rect 27192 41856 27256 41860
rect 31952 41916 32016 41920
rect 31952 41860 31956 41916
rect 31956 41860 32012 41916
rect 32012 41860 32016 41916
rect 31952 41856 32016 41860
rect 32032 41916 32096 41920
rect 32032 41860 32036 41916
rect 32036 41860 32092 41916
rect 32092 41860 32096 41916
rect 32032 41856 32096 41860
rect 32112 41916 32176 41920
rect 32112 41860 32116 41916
rect 32116 41860 32172 41916
rect 32172 41860 32176 41916
rect 32112 41856 32176 41860
rect 32192 41916 32256 41920
rect 32192 41860 32196 41916
rect 32196 41860 32252 41916
rect 32252 41860 32256 41916
rect 32192 41856 32256 41860
rect 36952 41916 37016 41920
rect 36952 41860 36956 41916
rect 36956 41860 37012 41916
rect 37012 41860 37016 41916
rect 36952 41856 37016 41860
rect 37032 41916 37096 41920
rect 37032 41860 37036 41916
rect 37036 41860 37092 41916
rect 37092 41860 37096 41916
rect 37032 41856 37096 41860
rect 37112 41916 37176 41920
rect 37112 41860 37116 41916
rect 37116 41860 37172 41916
rect 37172 41860 37176 41916
rect 37112 41856 37176 41860
rect 37192 41916 37256 41920
rect 37192 41860 37196 41916
rect 37196 41860 37252 41916
rect 37252 41860 37256 41916
rect 37192 41856 37256 41860
rect 41952 41916 42016 41920
rect 41952 41860 41956 41916
rect 41956 41860 42012 41916
rect 42012 41860 42016 41916
rect 41952 41856 42016 41860
rect 42032 41916 42096 41920
rect 42032 41860 42036 41916
rect 42036 41860 42092 41916
rect 42092 41860 42096 41916
rect 42032 41856 42096 41860
rect 42112 41916 42176 41920
rect 42112 41860 42116 41916
rect 42116 41860 42172 41916
rect 42172 41860 42176 41916
rect 42112 41856 42176 41860
rect 42192 41916 42256 41920
rect 42192 41860 42196 41916
rect 42196 41860 42252 41916
rect 42252 41860 42256 41916
rect 42192 41856 42256 41860
rect 46952 41916 47016 41920
rect 46952 41860 46956 41916
rect 46956 41860 47012 41916
rect 47012 41860 47016 41916
rect 46952 41856 47016 41860
rect 47032 41916 47096 41920
rect 47032 41860 47036 41916
rect 47036 41860 47092 41916
rect 47092 41860 47096 41916
rect 47032 41856 47096 41860
rect 47112 41916 47176 41920
rect 47112 41860 47116 41916
rect 47116 41860 47172 41916
rect 47172 41860 47176 41916
rect 47112 41856 47176 41860
rect 47192 41916 47256 41920
rect 47192 41860 47196 41916
rect 47196 41860 47252 41916
rect 47252 41860 47256 41916
rect 47192 41856 47256 41860
rect 51952 41916 52016 41920
rect 51952 41860 51956 41916
rect 51956 41860 52012 41916
rect 52012 41860 52016 41916
rect 51952 41856 52016 41860
rect 52032 41916 52096 41920
rect 52032 41860 52036 41916
rect 52036 41860 52092 41916
rect 52092 41860 52096 41916
rect 52032 41856 52096 41860
rect 52112 41916 52176 41920
rect 52112 41860 52116 41916
rect 52116 41860 52172 41916
rect 52172 41860 52176 41916
rect 52112 41856 52176 41860
rect 52192 41916 52256 41920
rect 52192 41860 52196 41916
rect 52196 41860 52252 41916
rect 52252 41860 52256 41916
rect 52192 41856 52256 41860
rect 56952 41916 57016 41920
rect 56952 41860 56956 41916
rect 56956 41860 57012 41916
rect 57012 41860 57016 41916
rect 56952 41856 57016 41860
rect 57032 41916 57096 41920
rect 57032 41860 57036 41916
rect 57036 41860 57092 41916
rect 57092 41860 57096 41916
rect 57032 41856 57096 41860
rect 57112 41916 57176 41920
rect 57112 41860 57116 41916
rect 57116 41860 57172 41916
rect 57172 41860 57176 41916
rect 57112 41856 57176 41860
rect 57192 41916 57256 41920
rect 57192 41860 57196 41916
rect 57196 41860 57252 41916
rect 57252 41860 57256 41916
rect 57192 41856 57256 41860
rect 2612 41372 2676 41376
rect 2612 41316 2616 41372
rect 2616 41316 2672 41372
rect 2672 41316 2676 41372
rect 2612 41312 2676 41316
rect 2692 41372 2756 41376
rect 2692 41316 2696 41372
rect 2696 41316 2752 41372
rect 2752 41316 2756 41372
rect 2692 41312 2756 41316
rect 2772 41372 2836 41376
rect 2772 41316 2776 41372
rect 2776 41316 2832 41372
rect 2832 41316 2836 41372
rect 2772 41312 2836 41316
rect 2852 41372 2916 41376
rect 2852 41316 2856 41372
rect 2856 41316 2912 41372
rect 2912 41316 2916 41372
rect 2852 41312 2916 41316
rect 7612 41372 7676 41376
rect 7612 41316 7616 41372
rect 7616 41316 7672 41372
rect 7672 41316 7676 41372
rect 7612 41312 7676 41316
rect 7692 41372 7756 41376
rect 7692 41316 7696 41372
rect 7696 41316 7752 41372
rect 7752 41316 7756 41372
rect 7692 41312 7756 41316
rect 7772 41372 7836 41376
rect 7772 41316 7776 41372
rect 7776 41316 7832 41372
rect 7832 41316 7836 41372
rect 7772 41312 7836 41316
rect 7852 41372 7916 41376
rect 7852 41316 7856 41372
rect 7856 41316 7912 41372
rect 7912 41316 7916 41372
rect 7852 41312 7916 41316
rect 12612 41372 12676 41376
rect 12612 41316 12616 41372
rect 12616 41316 12672 41372
rect 12672 41316 12676 41372
rect 12612 41312 12676 41316
rect 12692 41372 12756 41376
rect 12692 41316 12696 41372
rect 12696 41316 12752 41372
rect 12752 41316 12756 41372
rect 12692 41312 12756 41316
rect 12772 41372 12836 41376
rect 12772 41316 12776 41372
rect 12776 41316 12832 41372
rect 12832 41316 12836 41372
rect 12772 41312 12836 41316
rect 12852 41372 12916 41376
rect 12852 41316 12856 41372
rect 12856 41316 12912 41372
rect 12912 41316 12916 41372
rect 12852 41312 12916 41316
rect 17612 41372 17676 41376
rect 17612 41316 17616 41372
rect 17616 41316 17672 41372
rect 17672 41316 17676 41372
rect 17612 41312 17676 41316
rect 17692 41372 17756 41376
rect 17692 41316 17696 41372
rect 17696 41316 17752 41372
rect 17752 41316 17756 41372
rect 17692 41312 17756 41316
rect 17772 41372 17836 41376
rect 17772 41316 17776 41372
rect 17776 41316 17832 41372
rect 17832 41316 17836 41372
rect 17772 41312 17836 41316
rect 17852 41372 17916 41376
rect 17852 41316 17856 41372
rect 17856 41316 17912 41372
rect 17912 41316 17916 41372
rect 17852 41312 17916 41316
rect 22612 41372 22676 41376
rect 22612 41316 22616 41372
rect 22616 41316 22672 41372
rect 22672 41316 22676 41372
rect 22612 41312 22676 41316
rect 22692 41372 22756 41376
rect 22692 41316 22696 41372
rect 22696 41316 22752 41372
rect 22752 41316 22756 41372
rect 22692 41312 22756 41316
rect 22772 41372 22836 41376
rect 22772 41316 22776 41372
rect 22776 41316 22832 41372
rect 22832 41316 22836 41372
rect 22772 41312 22836 41316
rect 22852 41372 22916 41376
rect 22852 41316 22856 41372
rect 22856 41316 22912 41372
rect 22912 41316 22916 41372
rect 22852 41312 22916 41316
rect 27612 41372 27676 41376
rect 27612 41316 27616 41372
rect 27616 41316 27672 41372
rect 27672 41316 27676 41372
rect 27612 41312 27676 41316
rect 27692 41372 27756 41376
rect 27692 41316 27696 41372
rect 27696 41316 27752 41372
rect 27752 41316 27756 41372
rect 27692 41312 27756 41316
rect 27772 41372 27836 41376
rect 27772 41316 27776 41372
rect 27776 41316 27832 41372
rect 27832 41316 27836 41372
rect 27772 41312 27836 41316
rect 27852 41372 27916 41376
rect 27852 41316 27856 41372
rect 27856 41316 27912 41372
rect 27912 41316 27916 41372
rect 27852 41312 27916 41316
rect 32612 41372 32676 41376
rect 32612 41316 32616 41372
rect 32616 41316 32672 41372
rect 32672 41316 32676 41372
rect 32612 41312 32676 41316
rect 32692 41372 32756 41376
rect 32692 41316 32696 41372
rect 32696 41316 32752 41372
rect 32752 41316 32756 41372
rect 32692 41312 32756 41316
rect 32772 41372 32836 41376
rect 32772 41316 32776 41372
rect 32776 41316 32832 41372
rect 32832 41316 32836 41372
rect 32772 41312 32836 41316
rect 32852 41372 32916 41376
rect 32852 41316 32856 41372
rect 32856 41316 32912 41372
rect 32912 41316 32916 41372
rect 32852 41312 32916 41316
rect 37612 41372 37676 41376
rect 37612 41316 37616 41372
rect 37616 41316 37672 41372
rect 37672 41316 37676 41372
rect 37612 41312 37676 41316
rect 37692 41372 37756 41376
rect 37692 41316 37696 41372
rect 37696 41316 37752 41372
rect 37752 41316 37756 41372
rect 37692 41312 37756 41316
rect 37772 41372 37836 41376
rect 37772 41316 37776 41372
rect 37776 41316 37832 41372
rect 37832 41316 37836 41372
rect 37772 41312 37836 41316
rect 37852 41372 37916 41376
rect 37852 41316 37856 41372
rect 37856 41316 37912 41372
rect 37912 41316 37916 41372
rect 37852 41312 37916 41316
rect 42612 41372 42676 41376
rect 42612 41316 42616 41372
rect 42616 41316 42672 41372
rect 42672 41316 42676 41372
rect 42612 41312 42676 41316
rect 42692 41372 42756 41376
rect 42692 41316 42696 41372
rect 42696 41316 42752 41372
rect 42752 41316 42756 41372
rect 42692 41312 42756 41316
rect 42772 41372 42836 41376
rect 42772 41316 42776 41372
rect 42776 41316 42832 41372
rect 42832 41316 42836 41372
rect 42772 41312 42836 41316
rect 42852 41372 42916 41376
rect 42852 41316 42856 41372
rect 42856 41316 42912 41372
rect 42912 41316 42916 41372
rect 42852 41312 42916 41316
rect 47612 41372 47676 41376
rect 47612 41316 47616 41372
rect 47616 41316 47672 41372
rect 47672 41316 47676 41372
rect 47612 41312 47676 41316
rect 47692 41372 47756 41376
rect 47692 41316 47696 41372
rect 47696 41316 47752 41372
rect 47752 41316 47756 41372
rect 47692 41312 47756 41316
rect 47772 41372 47836 41376
rect 47772 41316 47776 41372
rect 47776 41316 47832 41372
rect 47832 41316 47836 41372
rect 47772 41312 47836 41316
rect 47852 41372 47916 41376
rect 47852 41316 47856 41372
rect 47856 41316 47912 41372
rect 47912 41316 47916 41372
rect 47852 41312 47916 41316
rect 52612 41372 52676 41376
rect 52612 41316 52616 41372
rect 52616 41316 52672 41372
rect 52672 41316 52676 41372
rect 52612 41312 52676 41316
rect 52692 41372 52756 41376
rect 52692 41316 52696 41372
rect 52696 41316 52752 41372
rect 52752 41316 52756 41372
rect 52692 41312 52756 41316
rect 52772 41372 52836 41376
rect 52772 41316 52776 41372
rect 52776 41316 52832 41372
rect 52832 41316 52836 41372
rect 52772 41312 52836 41316
rect 52852 41372 52916 41376
rect 52852 41316 52856 41372
rect 52856 41316 52912 41372
rect 52912 41316 52916 41372
rect 52852 41312 52916 41316
rect 57612 41372 57676 41376
rect 57612 41316 57616 41372
rect 57616 41316 57672 41372
rect 57672 41316 57676 41372
rect 57612 41312 57676 41316
rect 57692 41372 57756 41376
rect 57692 41316 57696 41372
rect 57696 41316 57752 41372
rect 57752 41316 57756 41372
rect 57692 41312 57756 41316
rect 57772 41372 57836 41376
rect 57772 41316 57776 41372
rect 57776 41316 57832 41372
rect 57832 41316 57836 41372
rect 57772 41312 57836 41316
rect 57852 41372 57916 41376
rect 57852 41316 57856 41372
rect 57856 41316 57912 41372
rect 57912 41316 57916 41372
rect 57852 41312 57916 41316
rect 1952 40828 2016 40832
rect 1952 40772 1956 40828
rect 1956 40772 2012 40828
rect 2012 40772 2016 40828
rect 1952 40768 2016 40772
rect 2032 40828 2096 40832
rect 2032 40772 2036 40828
rect 2036 40772 2092 40828
rect 2092 40772 2096 40828
rect 2032 40768 2096 40772
rect 2112 40828 2176 40832
rect 2112 40772 2116 40828
rect 2116 40772 2172 40828
rect 2172 40772 2176 40828
rect 2112 40768 2176 40772
rect 2192 40828 2256 40832
rect 2192 40772 2196 40828
rect 2196 40772 2252 40828
rect 2252 40772 2256 40828
rect 2192 40768 2256 40772
rect 6952 40828 7016 40832
rect 6952 40772 6956 40828
rect 6956 40772 7012 40828
rect 7012 40772 7016 40828
rect 6952 40768 7016 40772
rect 7032 40828 7096 40832
rect 7032 40772 7036 40828
rect 7036 40772 7092 40828
rect 7092 40772 7096 40828
rect 7032 40768 7096 40772
rect 7112 40828 7176 40832
rect 7112 40772 7116 40828
rect 7116 40772 7172 40828
rect 7172 40772 7176 40828
rect 7112 40768 7176 40772
rect 7192 40828 7256 40832
rect 7192 40772 7196 40828
rect 7196 40772 7252 40828
rect 7252 40772 7256 40828
rect 7192 40768 7256 40772
rect 11952 40828 12016 40832
rect 11952 40772 11956 40828
rect 11956 40772 12012 40828
rect 12012 40772 12016 40828
rect 11952 40768 12016 40772
rect 12032 40828 12096 40832
rect 12032 40772 12036 40828
rect 12036 40772 12092 40828
rect 12092 40772 12096 40828
rect 12032 40768 12096 40772
rect 12112 40828 12176 40832
rect 12112 40772 12116 40828
rect 12116 40772 12172 40828
rect 12172 40772 12176 40828
rect 12112 40768 12176 40772
rect 12192 40828 12256 40832
rect 12192 40772 12196 40828
rect 12196 40772 12252 40828
rect 12252 40772 12256 40828
rect 12192 40768 12256 40772
rect 16952 40828 17016 40832
rect 16952 40772 16956 40828
rect 16956 40772 17012 40828
rect 17012 40772 17016 40828
rect 16952 40768 17016 40772
rect 17032 40828 17096 40832
rect 17032 40772 17036 40828
rect 17036 40772 17092 40828
rect 17092 40772 17096 40828
rect 17032 40768 17096 40772
rect 17112 40828 17176 40832
rect 17112 40772 17116 40828
rect 17116 40772 17172 40828
rect 17172 40772 17176 40828
rect 17112 40768 17176 40772
rect 17192 40828 17256 40832
rect 17192 40772 17196 40828
rect 17196 40772 17252 40828
rect 17252 40772 17256 40828
rect 17192 40768 17256 40772
rect 21952 40828 22016 40832
rect 21952 40772 21956 40828
rect 21956 40772 22012 40828
rect 22012 40772 22016 40828
rect 21952 40768 22016 40772
rect 22032 40828 22096 40832
rect 22032 40772 22036 40828
rect 22036 40772 22092 40828
rect 22092 40772 22096 40828
rect 22032 40768 22096 40772
rect 22112 40828 22176 40832
rect 22112 40772 22116 40828
rect 22116 40772 22172 40828
rect 22172 40772 22176 40828
rect 22112 40768 22176 40772
rect 22192 40828 22256 40832
rect 22192 40772 22196 40828
rect 22196 40772 22252 40828
rect 22252 40772 22256 40828
rect 22192 40768 22256 40772
rect 26952 40828 27016 40832
rect 26952 40772 26956 40828
rect 26956 40772 27012 40828
rect 27012 40772 27016 40828
rect 26952 40768 27016 40772
rect 27032 40828 27096 40832
rect 27032 40772 27036 40828
rect 27036 40772 27092 40828
rect 27092 40772 27096 40828
rect 27032 40768 27096 40772
rect 27112 40828 27176 40832
rect 27112 40772 27116 40828
rect 27116 40772 27172 40828
rect 27172 40772 27176 40828
rect 27112 40768 27176 40772
rect 27192 40828 27256 40832
rect 27192 40772 27196 40828
rect 27196 40772 27252 40828
rect 27252 40772 27256 40828
rect 27192 40768 27256 40772
rect 31952 40828 32016 40832
rect 31952 40772 31956 40828
rect 31956 40772 32012 40828
rect 32012 40772 32016 40828
rect 31952 40768 32016 40772
rect 32032 40828 32096 40832
rect 32032 40772 32036 40828
rect 32036 40772 32092 40828
rect 32092 40772 32096 40828
rect 32032 40768 32096 40772
rect 32112 40828 32176 40832
rect 32112 40772 32116 40828
rect 32116 40772 32172 40828
rect 32172 40772 32176 40828
rect 32112 40768 32176 40772
rect 32192 40828 32256 40832
rect 32192 40772 32196 40828
rect 32196 40772 32252 40828
rect 32252 40772 32256 40828
rect 32192 40768 32256 40772
rect 36952 40828 37016 40832
rect 36952 40772 36956 40828
rect 36956 40772 37012 40828
rect 37012 40772 37016 40828
rect 36952 40768 37016 40772
rect 37032 40828 37096 40832
rect 37032 40772 37036 40828
rect 37036 40772 37092 40828
rect 37092 40772 37096 40828
rect 37032 40768 37096 40772
rect 37112 40828 37176 40832
rect 37112 40772 37116 40828
rect 37116 40772 37172 40828
rect 37172 40772 37176 40828
rect 37112 40768 37176 40772
rect 37192 40828 37256 40832
rect 37192 40772 37196 40828
rect 37196 40772 37252 40828
rect 37252 40772 37256 40828
rect 37192 40768 37256 40772
rect 41952 40828 42016 40832
rect 41952 40772 41956 40828
rect 41956 40772 42012 40828
rect 42012 40772 42016 40828
rect 41952 40768 42016 40772
rect 42032 40828 42096 40832
rect 42032 40772 42036 40828
rect 42036 40772 42092 40828
rect 42092 40772 42096 40828
rect 42032 40768 42096 40772
rect 42112 40828 42176 40832
rect 42112 40772 42116 40828
rect 42116 40772 42172 40828
rect 42172 40772 42176 40828
rect 42112 40768 42176 40772
rect 42192 40828 42256 40832
rect 42192 40772 42196 40828
rect 42196 40772 42252 40828
rect 42252 40772 42256 40828
rect 42192 40768 42256 40772
rect 46952 40828 47016 40832
rect 46952 40772 46956 40828
rect 46956 40772 47012 40828
rect 47012 40772 47016 40828
rect 46952 40768 47016 40772
rect 47032 40828 47096 40832
rect 47032 40772 47036 40828
rect 47036 40772 47092 40828
rect 47092 40772 47096 40828
rect 47032 40768 47096 40772
rect 47112 40828 47176 40832
rect 47112 40772 47116 40828
rect 47116 40772 47172 40828
rect 47172 40772 47176 40828
rect 47112 40768 47176 40772
rect 47192 40828 47256 40832
rect 47192 40772 47196 40828
rect 47196 40772 47252 40828
rect 47252 40772 47256 40828
rect 47192 40768 47256 40772
rect 51952 40828 52016 40832
rect 51952 40772 51956 40828
rect 51956 40772 52012 40828
rect 52012 40772 52016 40828
rect 51952 40768 52016 40772
rect 52032 40828 52096 40832
rect 52032 40772 52036 40828
rect 52036 40772 52092 40828
rect 52092 40772 52096 40828
rect 52032 40768 52096 40772
rect 52112 40828 52176 40832
rect 52112 40772 52116 40828
rect 52116 40772 52172 40828
rect 52172 40772 52176 40828
rect 52112 40768 52176 40772
rect 52192 40828 52256 40832
rect 52192 40772 52196 40828
rect 52196 40772 52252 40828
rect 52252 40772 52256 40828
rect 52192 40768 52256 40772
rect 56952 40828 57016 40832
rect 56952 40772 56956 40828
rect 56956 40772 57012 40828
rect 57012 40772 57016 40828
rect 56952 40768 57016 40772
rect 57032 40828 57096 40832
rect 57032 40772 57036 40828
rect 57036 40772 57092 40828
rect 57092 40772 57096 40828
rect 57032 40768 57096 40772
rect 57112 40828 57176 40832
rect 57112 40772 57116 40828
rect 57116 40772 57172 40828
rect 57172 40772 57176 40828
rect 57112 40768 57176 40772
rect 57192 40828 57256 40832
rect 57192 40772 57196 40828
rect 57196 40772 57252 40828
rect 57252 40772 57256 40828
rect 57192 40768 57256 40772
rect 2612 40284 2676 40288
rect 2612 40228 2616 40284
rect 2616 40228 2672 40284
rect 2672 40228 2676 40284
rect 2612 40224 2676 40228
rect 2692 40284 2756 40288
rect 2692 40228 2696 40284
rect 2696 40228 2752 40284
rect 2752 40228 2756 40284
rect 2692 40224 2756 40228
rect 2772 40284 2836 40288
rect 2772 40228 2776 40284
rect 2776 40228 2832 40284
rect 2832 40228 2836 40284
rect 2772 40224 2836 40228
rect 2852 40284 2916 40288
rect 2852 40228 2856 40284
rect 2856 40228 2912 40284
rect 2912 40228 2916 40284
rect 2852 40224 2916 40228
rect 7612 40284 7676 40288
rect 7612 40228 7616 40284
rect 7616 40228 7672 40284
rect 7672 40228 7676 40284
rect 7612 40224 7676 40228
rect 7692 40284 7756 40288
rect 7692 40228 7696 40284
rect 7696 40228 7752 40284
rect 7752 40228 7756 40284
rect 7692 40224 7756 40228
rect 7772 40284 7836 40288
rect 7772 40228 7776 40284
rect 7776 40228 7832 40284
rect 7832 40228 7836 40284
rect 7772 40224 7836 40228
rect 7852 40284 7916 40288
rect 7852 40228 7856 40284
rect 7856 40228 7912 40284
rect 7912 40228 7916 40284
rect 7852 40224 7916 40228
rect 12612 40284 12676 40288
rect 12612 40228 12616 40284
rect 12616 40228 12672 40284
rect 12672 40228 12676 40284
rect 12612 40224 12676 40228
rect 12692 40284 12756 40288
rect 12692 40228 12696 40284
rect 12696 40228 12752 40284
rect 12752 40228 12756 40284
rect 12692 40224 12756 40228
rect 12772 40284 12836 40288
rect 12772 40228 12776 40284
rect 12776 40228 12832 40284
rect 12832 40228 12836 40284
rect 12772 40224 12836 40228
rect 12852 40284 12916 40288
rect 12852 40228 12856 40284
rect 12856 40228 12912 40284
rect 12912 40228 12916 40284
rect 12852 40224 12916 40228
rect 17612 40284 17676 40288
rect 17612 40228 17616 40284
rect 17616 40228 17672 40284
rect 17672 40228 17676 40284
rect 17612 40224 17676 40228
rect 17692 40284 17756 40288
rect 17692 40228 17696 40284
rect 17696 40228 17752 40284
rect 17752 40228 17756 40284
rect 17692 40224 17756 40228
rect 17772 40284 17836 40288
rect 17772 40228 17776 40284
rect 17776 40228 17832 40284
rect 17832 40228 17836 40284
rect 17772 40224 17836 40228
rect 17852 40284 17916 40288
rect 17852 40228 17856 40284
rect 17856 40228 17912 40284
rect 17912 40228 17916 40284
rect 17852 40224 17916 40228
rect 22612 40284 22676 40288
rect 22612 40228 22616 40284
rect 22616 40228 22672 40284
rect 22672 40228 22676 40284
rect 22612 40224 22676 40228
rect 22692 40284 22756 40288
rect 22692 40228 22696 40284
rect 22696 40228 22752 40284
rect 22752 40228 22756 40284
rect 22692 40224 22756 40228
rect 22772 40284 22836 40288
rect 22772 40228 22776 40284
rect 22776 40228 22832 40284
rect 22832 40228 22836 40284
rect 22772 40224 22836 40228
rect 22852 40284 22916 40288
rect 22852 40228 22856 40284
rect 22856 40228 22912 40284
rect 22912 40228 22916 40284
rect 22852 40224 22916 40228
rect 27612 40284 27676 40288
rect 27612 40228 27616 40284
rect 27616 40228 27672 40284
rect 27672 40228 27676 40284
rect 27612 40224 27676 40228
rect 27692 40284 27756 40288
rect 27692 40228 27696 40284
rect 27696 40228 27752 40284
rect 27752 40228 27756 40284
rect 27692 40224 27756 40228
rect 27772 40284 27836 40288
rect 27772 40228 27776 40284
rect 27776 40228 27832 40284
rect 27832 40228 27836 40284
rect 27772 40224 27836 40228
rect 27852 40284 27916 40288
rect 27852 40228 27856 40284
rect 27856 40228 27912 40284
rect 27912 40228 27916 40284
rect 27852 40224 27916 40228
rect 32612 40284 32676 40288
rect 32612 40228 32616 40284
rect 32616 40228 32672 40284
rect 32672 40228 32676 40284
rect 32612 40224 32676 40228
rect 32692 40284 32756 40288
rect 32692 40228 32696 40284
rect 32696 40228 32752 40284
rect 32752 40228 32756 40284
rect 32692 40224 32756 40228
rect 32772 40284 32836 40288
rect 32772 40228 32776 40284
rect 32776 40228 32832 40284
rect 32832 40228 32836 40284
rect 32772 40224 32836 40228
rect 32852 40284 32916 40288
rect 32852 40228 32856 40284
rect 32856 40228 32912 40284
rect 32912 40228 32916 40284
rect 32852 40224 32916 40228
rect 37612 40284 37676 40288
rect 37612 40228 37616 40284
rect 37616 40228 37672 40284
rect 37672 40228 37676 40284
rect 37612 40224 37676 40228
rect 37692 40284 37756 40288
rect 37692 40228 37696 40284
rect 37696 40228 37752 40284
rect 37752 40228 37756 40284
rect 37692 40224 37756 40228
rect 37772 40284 37836 40288
rect 37772 40228 37776 40284
rect 37776 40228 37832 40284
rect 37832 40228 37836 40284
rect 37772 40224 37836 40228
rect 37852 40284 37916 40288
rect 37852 40228 37856 40284
rect 37856 40228 37912 40284
rect 37912 40228 37916 40284
rect 37852 40224 37916 40228
rect 42612 40284 42676 40288
rect 42612 40228 42616 40284
rect 42616 40228 42672 40284
rect 42672 40228 42676 40284
rect 42612 40224 42676 40228
rect 42692 40284 42756 40288
rect 42692 40228 42696 40284
rect 42696 40228 42752 40284
rect 42752 40228 42756 40284
rect 42692 40224 42756 40228
rect 42772 40284 42836 40288
rect 42772 40228 42776 40284
rect 42776 40228 42832 40284
rect 42832 40228 42836 40284
rect 42772 40224 42836 40228
rect 42852 40284 42916 40288
rect 42852 40228 42856 40284
rect 42856 40228 42912 40284
rect 42912 40228 42916 40284
rect 42852 40224 42916 40228
rect 47612 40284 47676 40288
rect 47612 40228 47616 40284
rect 47616 40228 47672 40284
rect 47672 40228 47676 40284
rect 47612 40224 47676 40228
rect 47692 40284 47756 40288
rect 47692 40228 47696 40284
rect 47696 40228 47752 40284
rect 47752 40228 47756 40284
rect 47692 40224 47756 40228
rect 47772 40284 47836 40288
rect 47772 40228 47776 40284
rect 47776 40228 47832 40284
rect 47832 40228 47836 40284
rect 47772 40224 47836 40228
rect 47852 40284 47916 40288
rect 47852 40228 47856 40284
rect 47856 40228 47912 40284
rect 47912 40228 47916 40284
rect 47852 40224 47916 40228
rect 52612 40284 52676 40288
rect 52612 40228 52616 40284
rect 52616 40228 52672 40284
rect 52672 40228 52676 40284
rect 52612 40224 52676 40228
rect 52692 40284 52756 40288
rect 52692 40228 52696 40284
rect 52696 40228 52752 40284
rect 52752 40228 52756 40284
rect 52692 40224 52756 40228
rect 52772 40284 52836 40288
rect 52772 40228 52776 40284
rect 52776 40228 52832 40284
rect 52832 40228 52836 40284
rect 52772 40224 52836 40228
rect 52852 40284 52916 40288
rect 52852 40228 52856 40284
rect 52856 40228 52912 40284
rect 52912 40228 52916 40284
rect 52852 40224 52916 40228
rect 57612 40284 57676 40288
rect 57612 40228 57616 40284
rect 57616 40228 57672 40284
rect 57672 40228 57676 40284
rect 57612 40224 57676 40228
rect 57692 40284 57756 40288
rect 57692 40228 57696 40284
rect 57696 40228 57752 40284
rect 57752 40228 57756 40284
rect 57692 40224 57756 40228
rect 57772 40284 57836 40288
rect 57772 40228 57776 40284
rect 57776 40228 57832 40284
rect 57832 40228 57836 40284
rect 57772 40224 57836 40228
rect 57852 40284 57916 40288
rect 57852 40228 57856 40284
rect 57856 40228 57912 40284
rect 57912 40228 57916 40284
rect 57852 40224 57916 40228
rect 1952 39740 2016 39744
rect 1952 39684 1956 39740
rect 1956 39684 2012 39740
rect 2012 39684 2016 39740
rect 1952 39680 2016 39684
rect 2032 39740 2096 39744
rect 2032 39684 2036 39740
rect 2036 39684 2092 39740
rect 2092 39684 2096 39740
rect 2032 39680 2096 39684
rect 2112 39740 2176 39744
rect 2112 39684 2116 39740
rect 2116 39684 2172 39740
rect 2172 39684 2176 39740
rect 2112 39680 2176 39684
rect 2192 39740 2256 39744
rect 2192 39684 2196 39740
rect 2196 39684 2252 39740
rect 2252 39684 2256 39740
rect 2192 39680 2256 39684
rect 6952 39740 7016 39744
rect 6952 39684 6956 39740
rect 6956 39684 7012 39740
rect 7012 39684 7016 39740
rect 6952 39680 7016 39684
rect 7032 39740 7096 39744
rect 7032 39684 7036 39740
rect 7036 39684 7092 39740
rect 7092 39684 7096 39740
rect 7032 39680 7096 39684
rect 7112 39740 7176 39744
rect 7112 39684 7116 39740
rect 7116 39684 7172 39740
rect 7172 39684 7176 39740
rect 7112 39680 7176 39684
rect 7192 39740 7256 39744
rect 7192 39684 7196 39740
rect 7196 39684 7252 39740
rect 7252 39684 7256 39740
rect 7192 39680 7256 39684
rect 11952 39740 12016 39744
rect 11952 39684 11956 39740
rect 11956 39684 12012 39740
rect 12012 39684 12016 39740
rect 11952 39680 12016 39684
rect 12032 39740 12096 39744
rect 12032 39684 12036 39740
rect 12036 39684 12092 39740
rect 12092 39684 12096 39740
rect 12032 39680 12096 39684
rect 12112 39740 12176 39744
rect 12112 39684 12116 39740
rect 12116 39684 12172 39740
rect 12172 39684 12176 39740
rect 12112 39680 12176 39684
rect 12192 39740 12256 39744
rect 12192 39684 12196 39740
rect 12196 39684 12252 39740
rect 12252 39684 12256 39740
rect 12192 39680 12256 39684
rect 16952 39740 17016 39744
rect 16952 39684 16956 39740
rect 16956 39684 17012 39740
rect 17012 39684 17016 39740
rect 16952 39680 17016 39684
rect 17032 39740 17096 39744
rect 17032 39684 17036 39740
rect 17036 39684 17092 39740
rect 17092 39684 17096 39740
rect 17032 39680 17096 39684
rect 17112 39740 17176 39744
rect 17112 39684 17116 39740
rect 17116 39684 17172 39740
rect 17172 39684 17176 39740
rect 17112 39680 17176 39684
rect 17192 39740 17256 39744
rect 17192 39684 17196 39740
rect 17196 39684 17252 39740
rect 17252 39684 17256 39740
rect 17192 39680 17256 39684
rect 21952 39740 22016 39744
rect 21952 39684 21956 39740
rect 21956 39684 22012 39740
rect 22012 39684 22016 39740
rect 21952 39680 22016 39684
rect 22032 39740 22096 39744
rect 22032 39684 22036 39740
rect 22036 39684 22092 39740
rect 22092 39684 22096 39740
rect 22032 39680 22096 39684
rect 22112 39740 22176 39744
rect 22112 39684 22116 39740
rect 22116 39684 22172 39740
rect 22172 39684 22176 39740
rect 22112 39680 22176 39684
rect 22192 39740 22256 39744
rect 22192 39684 22196 39740
rect 22196 39684 22252 39740
rect 22252 39684 22256 39740
rect 22192 39680 22256 39684
rect 26952 39740 27016 39744
rect 26952 39684 26956 39740
rect 26956 39684 27012 39740
rect 27012 39684 27016 39740
rect 26952 39680 27016 39684
rect 27032 39740 27096 39744
rect 27032 39684 27036 39740
rect 27036 39684 27092 39740
rect 27092 39684 27096 39740
rect 27032 39680 27096 39684
rect 27112 39740 27176 39744
rect 27112 39684 27116 39740
rect 27116 39684 27172 39740
rect 27172 39684 27176 39740
rect 27112 39680 27176 39684
rect 27192 39740 27256 39744
rect 27192 39684 27196 39740
rect 27196 39684 27252 39740
rect 27252 39684 27256 39740
rect 27192 39680 27256 39684
rect 31952 39740 32016 39744
rect 31952 39684 31956 39740
rect 31956 39684 32012 39740
rect 32012 39684 32016 39740
rect 31952 39680 32016 39684
rect 32032 39740 32096 39744
rect 32032 39684 32036 39740
rect 32036 39684 32092 39740
rect 32092 39684 32096 39740
rect 32032 39680 32096 39684
rect 32112 39740 32176 39744
rect 32112 39684 32116 39740
rect 32116 39684 32172 39740
rect 32172 39684 32176 39740
rect 32112 39680 32176 39684
rect 32192 39740 32256 39744
rect 32192 39684 32196 39740
rect 32196 39684 32252 39740
rect 32252 39684 32256 39740
rect 32192 39680 32256 39684
rect 36952 39740 37016 39744
rect 36952 39684 36956 39740
rect 36956 39684 37012 39740
rect 37012 39684 37016 39740
rect 36952 39680 37016 39684
rect 37032 39740 37096 39744
rect 37032 39684 37036 39740
rect 37036 39684 37092 39740
rect 37092 39684 37096 39740
rect 37032 39680 37096 39684
rect 37112 39740 37176 39744
rect 37112 39684 37116 39740
rect 37116 39684 37172 39740
rect 37172 39684 37176 39740
rect 37112 39680 37176 39684
rect 37192 39740 37256 39744
rect 37192 39684 37196 39740
rect 37196 39684 37252 39740
rect 37252 39684 37256 39740
rect 37192 39680 37256 39684
rect 41952 39740 42016 39744
rect 41952 39684 41956 39740
rect 41956 39684 42012 39740
rect 42012 39684 42016 39740
rect 41952 39680 42016 39684
rect 42032 39740 42096 39744
rect 42032 39684 42036 39740
rect 42036 39684 42092 39740
rect 42092 39684 42096 39740
rect 42032 39680 42096 39684
rect 42112 39740 42176 39744
rect 42112 39684 42116 39740
rect 42116 39684 42172 39740
rect 42172 39684 42176 39740
rect 42112 39680 42176 39684
rect 42192 39740 42256 39744
rect 42192 39684 42196 39740
rect 42196 39684 42252 39740
rect 42252 39684 42256 39740
rect 42192 39680 42256 39684
rect 46952 39740 47016 39744
rect 46952 39684 46956 39740
rect 46956 39684 47012 39740
rect 47012 39684 47016 39740
rect 46952 39680 47016 39684
rect 47032 39740 47096 39744
rect 47032 39684 47036 39740
rect 47036 39684 47092 39740
rect 47092 39684 47096 39740
rect 47032 39680 47096 39684
rect 47112 39740 47176 39744
rect 47112 39684 47116 39740
rect 47116 39684 47172 39740
rect 47172 39684 47176 39740
rect 47112 39680 47176 39684
rect 47192 39740 47256 39744
rect 47192 39684 47196 39740
rect 47196 39684 47252 39740
rect 47252 39684 47256 39740
rect 47192 39680 47256 39684
rect 51952 39740 52016 39744
rect 51952 39684 51956 39740
rect 51956 39684 52012 39740
rect 52012 39684 52016 39740
rect 51952 39680 52016 39684
rect 52032 39740 52096 39744
rect 52032 39684 52036 39740
rect 52036 39684 52092 39740
rect 52092 39684 52096 39740
rect 52032 39680 52096 39684
rect 52112 39740 52176 39744
rect 52112 39684 52116 39740
rect 52116 39684 52172 39740
rect 52172 39684 52176 39740
rect 52112 39680 52176 39684
rect 52192 39740 52256 39744
rect 52192 39684 52196 39740
rect 52196 39684 52252 39740
rect 52252 39684 52256 39740
rect 52192 39680 52256 39684
rect 56952 39740 57016 39744
rect 56952 39684 56956 39740
rect 56956 39684 57012 39740
rect 57012 39684 57016 39740
rect 56952 39680 57016 39684
rect 57032 39740 57096 39744
rect 57032 39684 57036 39740
rect 57036 39684 57092 39740
rect 57092 39684 57096 39740
rect 57032 39680 57096 39684
rect 57112 39740 57176 39744
rect 57112 39684 57116 39740
rect 57116 39684 57172 39740
rect 57172 39684 57176 39740
rect 57112 39680 57176 39684
rect 57192 39740 57256 39744
rect 57192 39684 57196 39740
rect 57196 39684 57252 39740
rect 57252 39684 57256 39740
rect 57192 39680 57256 39684
rect 2612 39196 2676 39200
rect 2612 39140 2616 39196
rect 2616 39140 2672 39196
rect 2672 39140 2676 39196
rect 2612 39136 2676 39140
rect 2692 39196 2756 39200
rect 2692 39140 2696 39196
rect 2696 39140 2752 39196
rect 2752 39140 2756 39196
rect 2692 39136 2756 39140
rect 2772 39196 2836 39200
rect 2772 39140 2776 39196
rect 2776 39140 2832 39196
rect 2832 39140 2836 39196
rect 2772 39136 2836 39140
rect 2852 39196 2916 39200
rect 2852 39140 2856 39196
rect 2856 39140 2912 39196
rect 2912 39140 2916 39196
rect 2852 39136 2916 39140
rect 7612 39196 7676 39200
rect 7612 39140 7616 39196
rect 7616 39140 7672 39196
rect 7672 39140 7676 39196
rect 7612 39136 7676 39140
rect 7692 39196 7756 39200
rect 7692 39140 7696 39196
rect 7696 39140 7752 39196
rect 7752 39140 7756 39196
rect 7692 39136 7756 39140
rect 7772 39196 7836 39200
rect 7772 39140 7776 39196
rect 7776 39140 7832 39196
rect 7832 39140 7836 39196
rect 7772 39136 7836 39140
rect 7852 39196 7916 39200
rect 7852 39140 7856 39196
rect 7856 39140 7912 39196
rect 7912 39140 7916 39196
rect 7852 39136 7916 39140
rect 12612 39196 12676 39200
rect 12612 39140 12616 39196
rect 12616 39140 12672 39196
rect 12672 39140 12676 39196
rect 12612 39136 12676 39140
rect 12692 39196 12756 39200
rect 12692 39140 12696 39196
rect 12696 39140 12752 39196
rect 12752 39140 12756 39196
rect 12692 39136 12756 39140
rect 12772 39196 12836 39200
rect 12772 39140 12776 39196
rect 12776 39140 12832 39196
rect 12832 39140 12836 39196
rect 12772 39136 12836 39140
rect 12852 39196 12916 39200
rect 12852 39140 12856 39196
rect 12856 39140 12912 39196
rect 12912 39140 12916 39196
rect 12852 39136 12916 39140
rect 17612 39196 17676 39200
rect 17612 39140 17616 39196
rect 17616 39140 17672 39196
rect 17672 39140 17676 39196
rect 17612 39136 17676 39140
rect 17692 39196 17756 39200
rect 17692 39140 17696 39196
rect 17696 39140 17752 39196
rect 17752 39140 17756 39196
rect 17692 39136 17756 39140
rect 17772 39196 17836 39200
rect 17772 39140 17776 39196
rect 17776 39140 17832 39196
rect 17832 39140 17836 39196
rect 17772 39136 17836 39140
rect 17852 39196 17916 39200
rect 17852 39140 17856 39196
rect 17856 39140 17912 39196
rect 17912 39140 17916 39196
rect 17852 39136 17916 39140
rect 22612 39196 22676 39200
rect 22612 39140 22616 39196
rect 22616 39140 22672 39196
rect 22672 39140 22676 39196
rect 22612 39136 22676 39140
rect 22692 39196 22756 39200
rect 22692 39140 22696 39196
rect 22696 39140 22752 39196
rect 22752 39140 22756 39196
rect 22692 39136 22756 39140
rect 22772 39196 22836 39200
rect 22772 39140 22776 39196
rect 22776 39140 22832 39196
rect 22832 39140 22836 39196
rect 22772 39136 22836 39140
rect 22852 39196 22916 39200
rect 22852 39140 22856 39196
rect 22856 39140 22912 39196
rect 22912 39140 22916 39196
rect 22852 39136 22916 39140
rect 27612 39196 27676 39200
rect 27612 39140 27616 39196
rect 27616 39140 27672 39196
rect 27672 39140 27676 39196
rect 27612 39136 27676 39140
rect 27692 39196 27756 39200
rect 27692 39140 27696 39196
rect 27696 39140 27752 39196
rect 27752 39140 27756 39196
rect 27692 39136 27756 39140
rect 27772 39196 27836 39200
rect 27772 39140 27776 39196
rect 27776 39140 27832 39196
rect 27832 39140 27836 39196
rect 27772 39136 27836 39140
rect 27852 39196 27916 39200
rect 27852 39140 27856 39196
rect 27856 39140 27912 39196
rect 27912 39140 27916 39196
rect 27852 39136 27916 39140
rect 32612 39196 32676 39200
rect 32612 39140 32616 39196
rect 32616 39140 32672 39196
rect 32672 39140 32676 39196
rect 32612 39136 32676 39140
rect 32692 39196 32756 39200
rect 32692 39140 32696 39196
rect 32696 39140 32752 39196
rect 32752 39140 32756 39196
rect 32692 39136 32756 39140
rect 32772 39196 32836 39200
rect 32772 39140 32776 39196
rect 32776 39140 32832 39196
rect 32832 39140 32836 39196
rect 32772 39136 32836 39140
rect 32852 39196 32916 39200
rect 32852 39140 32856 39196
rect 32856 39140 32912 39196
rect 32912 39140 32916 39196
rect 32852 39136 32916 39140
rect 37612 39196 37676 39200
rect 37612 39140 37616 39196
rect 37616 39140 37672 39196
rect 37672 39140 37676 39196
rect 37612 39136 37676 39140
rect 37692 39196 37756 39200
rect 37692 39140 37696 39196
rect 37696 39140 37752 39196
rect 37752 39140 37756 39196
rect 37692 39136 37756 39140
rect 37772 39196 37836 39200
rect 37772 39140 37776 39196
rect 37776 39140 37832 39196
rect 37832 39140 37836 39196
rect 37772 39136 37836 39140
rect 37852 39196 37916 39200
rect 37852 39140 37856 39196
rect 37856 39140 37912 39196
rect 37912 39140 37916 39196
rect 37852 39136 37916 39140
rect 42612 39196 42676 39200
rect 42612 39140 42616 39196
rect 42616 39140 42672 39196
rect 42672 39140 42676 39196
rect 42612 39136 42676 39140
rect 42692 39196 42756 39200
rect 42692 39140 42696 39196
rect 42696 39140 42752 39196
rect 42752 39140 42756 39196
rect 42692 39136 42756 39140
rect 42772 39196 42836 39200
rect 42772 39140 42776 39196
rect 42776 39140 42832 39196
rect 42832 39140 42836 39196
rect 42772 39136 42836 39140
rect 42852 39196 42916 39200
rect 42852 39140 42856 39196
rect 42856 39140 42912 39196
rect 42912 39140 42916 39196
rect 42852 39136 42916 39140
rect 47612 39196 47676 39200
rect 47612 39140 47616 39196
rect 47616 39140 47672 39196
rect 47672 39140 47676 39196
rect 47612 39136 47676 39140
rect 47692 39196 47756 39200
rect 47692 39140 47696 39196
rect 47696 39140 47752 39196
rect 47752 39140 47756 39196
rect 47692 39136 47756 39140
rect 47772 39196 47836 39200
rect 47772 39140 47776 39196
rect 47776 39140 47832 39196
rect 47832 39140 47836 39196
rect 47772 39136 47836 39140
rect 47852 39196 47916 39200
rect 47852 39140 47856 39196
rect 47856 39140 47912 39196
rect 47912 39140 47916 39196
rect 47852 39136 47916 39140
rect 52612 39196 52676 39200
rect 52612 39140 52616 39196
rect 52616 39140 52672 39196
rect 52672 39140 52676 39196
rect 52612 39136 52676 39140
rect 52692 39196 52756 39200
rect 52692 39140 52696 39196
rect 52696 39140 52752 39196
rect 52752 39140 52756 39196
rect 52692 39136 52756 39140
rect 52772 39196 52836 39200
rect 52772 39140 52776 39196
rect 52776 39140 52832 39196
rect 52832 39140 52836 39196
rect 52772 39136 52836 39140
rect 52852 39196 52916 39200
rect 52852 39140 52856 39196
rect 52856 39140 52912 39196
rect 52912 39140 52916 39196
rect 52852 39136 52916 39140
rect 57612 39196 57676 39200
rect 57612 39140 57616 39196
rect 57616 39140 57672 39196
rect 57672 39140 57676 39196
rect 57612 39136 57676 39140
rect 57692 39196 57756 39200
rect 57692 39140 57696 39196
rect 57696 39140 57752 39196
rect 57752 39140 57756 39196
rect 57692 39136 57756 39140
rect 57772 39196 57836 39200
rect 57772 39140 57776 39196
rect 57776 39140 57832 39196
rect 57832 39140 57836 39196
rect 57772 39136 57836 39140
rect 57852 39196 57916 39200
rect 57852 39140 57856 39196
rect 57856 39140 57912 39196
rect 57912 39140 57916 39196
rect 57852 39136 57916 39140
rect 1952 38652 2016 38656
rect 1952 38596 1956 38652
rect 1956 38596 2012 38652
rect 2012 38596 2016 38652
rect 1952 38592 2016 38596
rect 2032 38652 2096 38656
rect 2032 38596 2036 38652
rect 2036 38596 2092 38652
rect 2092 38596 2096 38652
rect 2032 38592 2096 38596
rect 2112 38652 2176 38656
rect 2112 38596 2116 38652
rect 2116 38596 2172 38652
rect 2172 38596 2176 38652
rect 2112 38592 2176 38596
rect 2192 38652 2256 38656
rect 2192 38596 2196 38652
rect 2196 38596 2252 38652
rect 2252 38596 2256 38652
rect 2192 38592 2256 38596
rect 6952 38652 7016 38656
rect 6952 38596 6956 38652
rect 6956 38596 7012 38652
rect 7012 38596 7016 38652
rect 6952 38592 7016 38596
rect 7032 38652 7096 38656
rect 7032 38596 7036 38652
rect 7036 38596 7092 38652
rect 7092 38596 7096 38652
rect 7032 38592 7096 38596
rect 7112 38652 7176 38656
rect 7112 38596 7116 38652
rect 7116 38596 7172 38652
rect 7172 38596 7176 38652
rect 7112 38592 7176 38596
rect 7192 38652 7256 38656
rect 7192 38596 7196 38652
rect 7196 38596 7252 38652
rect 7252 38596 7256 38652
rect 7192 38592 7256 38596
rect 11952 38652 12016 38656
rect 11952 38596 11956 38652
rect 11956 38596 12012 38652
rect 12012 38596 12016 38652
rect 11952 38592 12016 38596
rect 12032 38652 12096 38656
rect 12032 38596 12036 38652
rect 12036 38596 12092 38652
rect 12092 38596 12096 38652
rect 12032 38592 12096 38596
rect 12112 38652 12176 38656
rect 12112 38596 12116 38652
rect 12116 38596 12172 38652
rect 12172 38596 12176 38652
rect 12112 38592 12176 38596
rect 12192 38652 12256 38656
rect 12192 38596 12196 38652
rect 12196 38596 12252 38652
rect 12252 38596 12256 38652
rect 12192 38592 12256 38596
rect 16952 38652 17016 38656
rect 16952 38596 16956 38652
rect 16956 38596 17012 38652
rect 17012 38596 17016 38652
rect 16952 38592 17016 38596
rect 17032 38652 17096 38656
rect 17032 38596 17036 38652
rect 17036 38596 17092 38652
rect 17092 38596 17096 38652
rect 17032 38592 17096 38596
rect 17112 38652 17176 38656
rect 17112 38596 17116 38652
rect 17116 38596 17172 38652
rect 17172 38596 17176 38652
rect 17112 38592 17176 38596
rect 17192 38652 17256 38656
rect 17192 38596 17196 38652
rect 17196 38596 17252 38652
rect 17252 38596 17256 38652
rect 17192 38592 17256 38596
rect 21952 38652 22016 38656
rect 21952 38596 21956 38652
rect 21956 38596 22012 38652
rect 22012 38596 22016 38652
rect 21952 38592 22016 38596
rect 22032 38652 22096 38656
rect 22032 38596 22036 38652
rect 22036 38596 22092 38652
rect 22092 38596 22096 38652
rect 22032 38592 22096 38596
rect 22112 38652 22176 38656
rect 22112 38596 22116 38652
rect 22116 38596 22172 38652
rect 22172 38596 22176 38652
rect 22112 38592 22176 38596
rect 22192 38652 22256 38656
rect 22192 38596 22196 38652
rect 22196 38596 22252 38652
rect 22252 38596 22256 38652
rect 22192 38592 22256 38596
rect 26952 38652 27016 38656
rect 26952 38596 26956 38652
rect 26956 38596 27012 38652
rect 27012 38596 27016 38652
rect 26952 38592 27016 38596
rect 27032 38652 27096 38656
rect 27032 38596 27036 38652
rect 27036 38596 27092 38652
rect 27092 38596 27096 38652
rect 27032 38592 27096 38596
rect 27112 38652 27176 38656
rect 27112 38596 27116 38652
rect 27116 38596 27172 38652
rect 27172 38596 27176 38652
rect 27112 38592 27176 38596
rect 27192 38652 27256 38656
rect 27192 38596 27196 38652
rect 27196 38596 27252 38652
rect 27252 38596 27256 38652
rect 27192 38592 27256 38596
rect 31952 38652 32016 38656
rect 31952 38596 31956 38652
rect 31956 38596 32012 38652
rect 32012 38596 32016 38652
rect 31952 38592 32016 38596
rect 32032 38652 32096 38656
rect 32032 38596 32036 38652
rect 32036 38596 32092 38652
rect 32092 38596 32096 38652
rect 32032 38592 32096 38596
rect 32112 38652 32176 38656
rect 32112 38596 32116 38652
rect 32116 38596 32172 38652
rect 32172 38596 32176 38652
rect 32112 38592 32176 38596
rect 32192 38652 32256 38656
rect 32192 38596 32196 38652
rect 32196 38596 32252 38652
rect 32252 38596 32256 38652
rect 32192 38592 32256 38596
rect 36952 38652 37016 38656
rect 36952 38596 36956 38652
rect 36956 38596 37012 38652
rect 37012 38596 37016 38652
rect 36952 38592 37016 38596
rect 37032 38652 37096 38656
rect 37032 38596 37036 38652
rect 37036 38596 37092 38652
rect 37092 38596 37096 38652
rect 37032 38592 37096 38596
rect 37112 38652 37176 38656
rect 37112 38596 37116 38652
rect 37116 38596 37172 38652
rect 37172 38596 37176 38652
rect 37112 38592 37176 38596
rect 37192 38652 37256 38656
rect 37192 38596 37196 38652
rect 37196 38596 37252 38652
rect 37252 38596 37256 38652
rect 37192 38592 37256 38596
rect 41952 38652 42016 38656
rect 41952 38596 41956 38652
rect 41956 38596 42012 38652
rect 42012 38596 42016 38652
rect 41952 38592 42016 38596
rect 42032 38652 42096 38656
rect 42032 38596 42036 38652
rect 42036 38596 42092 38652
rect 42092 38596 42096 38652
rect 42032 38592 42096 38596
rect 42112 38652 42176 38656
rect 42112 38596 42116 38652
rect 42116 38596 42172 38652
rect 42172 38596 42176 38652
rect 42112 38592 42176 38596
rect 42192 38652 42256 38656
rect 42192 38596 42196 38652
rect 42196 38596 42252 38652
rect 42252 38596 42256 38652
rect 42192 38592 42256 38596
rect 46952 38652 47016 38656
rect 46952 38596 46956 38652
rect 46956 38596 47012 38652
rect 47012 38596 47016 38652
rect 46952 38592 47016 38596
rect 47032 38652 47096 38656
rect 47032 38596 47036 38652
rect 47036 38596 47092 38652
rect 47092 38596 47096 38652
rect 47032 38592 47096 38596
rect 47112 38652 47176 38656
rect 47112 38596 47116 38652
rect 47116 38596 47172 38652
rect 47172 38596 47176 38652
rect 47112 38592 47176 38596
rect 47192 38652 47256 38656
rect 47192 38596 47196 38652
rect 47196 38596 47252 38652
rect 47252 38596 47256 38652
rect 47192 38592 47256 38596
rect 51952 38652 52016 38656
rect 51952 38596 51956 38652
rect 51956 38596 52012 38652
rect 52012 38596 52016 38652
rect 51952 38592 52016 38596
rect 52032 38652 52096 38656
rect 52032 38596 52036 38652
rect 52036 38596 52092 38652
rect 52092 38596 52096 38652
rect 52032 38592 52096 38596
rect 52112 38652 52176 38656
rect 52112 38596 52116 38652
rect 52116 38596 52172 38652
rect 52172 38596 52176 38652
rect 52112 38592 52176 38596
rect 52192 38652 52256 38656
rect 52192 38596 52196 38652
rect 52196 38596 52252 38652
rect 52252 38596 52256 38652
rect 52192 38592 52256 38596
rect 56952 38652 57016 38656
rect 56952 38596 56956 38652
rect 56956 38596 57012 38652
rect 57012 38596 57016 38652
rect 56952 38592 57016 38596
rect 57032 38652 57096 38656
rect 57032 38596 57036 38652
rect 57036 38596 57092 38652
rect 57092 38596 57096 38652
rect 57032 38592 57096 38596
rect 57112 38652 57176 38656
rect 57112 38596 57116 38652
rect 57116 38596 57172 38652
rect 57172 38596 57176 38652
rect 57112 38592 57176 38596
rect 57192 38652 57256 38656
rect 57192 38596 57196 38652
rect 57196 38596 57252 38652
rect 57252 38596 57256 38652
rect 57192 38592 57256 38596
rect 2612 38108 2676 38112
rect 2612 38052 2616 38108
rect 2616 38052 2672 38108
rect 2672 38052 2676 38108
rect 2612 38048 2676 38052
rect 2692 38108 2756 38112
rect 2692 38052 2696 38108
rect 2696 38052 2752 38108
rect 2752 38052 2756 38108
rect 2692 38048 2756 38052
rect 2772 38108 2836 38112
rect 2772 38052 2776 38108
rect 2776 38052 2832 38108
rect 2832 38052 2836 38108
rect 2772 38048 2836 38052
rect 2852 38108 2916 38112
rect 2852 38052 2856 38108
rect 2856 38052 2912 38108
rect 2912 38052 2916 38108
rect 2852 38048 2916 38052
rect 7612 38108 7676 38112
rect 7612 38052 7616 38108
rect 7616 38052 7672 38108
rect 7672 38052 7676 38108
rect 7612 38048 7676 38052
rect 7692 38108 7756 38112
rect 7692 38052 7696 38108
rect 7696 38052 7752 38108
rect 7752 38052 7756 38108
rect 7692 38048 7756 38052
rect 7772 38108 7836 38112
rect 7772 38052 7776 38108
rect 7776 38052 7832 38108
rect 7832 38052 7836 38108
rect 7772 38048 7836 38052
rect 7852 38108 7916 38112
rect 7852 38052 7856 38108
rect 7856 38052 7912 38108
rect 7912 38052 7916 38108
rect 7852 38048 7916 38052
rect 12612 38108 12676 38112
rect 12612 38052 12616 38108
rect 12616 38052 12672 38108
rect 12672 38052 12676 38108
rect 12612 38048 12676 38052
rect 12692 38108 12756 38112
rect 12692 38052 12696 38108
rect 12696 38052 12752 38108
rect 12752 38052 12756 38108
rect 12692 38048 12756 38052
rect 12772 38108 12836 38112
rect 12772 38052 12776 38108
rect 12776 38052 12832 38108
rect 12832 38052 12836 38108
rect 12772 38048 12836 38052
rect 12852 38108 12916 38112
rect 12852 38052 12856 38108
rect 12856 38052 12912 38108
rect 12912 38052 12916 38108
rect 12852 38048 12916 38052
rect 17612 38108 17676 38112
rect 17612 38052 17616 38108
rect 17616 38052 17672 38108
rect 17672 38052 17676 38108
rect 17612 38048 17676 38052
rect 17692 38108 17756 38112
rect 17692 38052 17696 38108
rect 17696 38052 17752 38108
rect 17752 38052 17756 38108
rect 17692 38048 17756 38052
rect 17772 38108 17836 38112
rect 17772 38052 17776 38108
rect 17776 38052 17832 38108
rect 17832 38052 17836 38108
rect 17772 38048 17836 38052
rect 17852 38108 17916 38112
rect 17852 38052 17856 38108
rect 17856 38052 17912 38108
rect 17912 38052 17916 38108
rect 17852 38048 17916 38052
rect 22612 38108 22676 38112
rect 22612 38052 22616 38108
rect 22616 38052 22672 38108
rect 22672 38052 22676 38108
rect 22612 38048 22676 38052
rect 22692 38108 22756 38112
rect 22692 38052 22696 38108
rect 22696 38052 22752 38108
rect 22752 38052 22756 38108
rect 22692 38048 22756 38052
rect 22772 38108 22836 38112
rect 22772 38052 22776 38108
rect 22776 38052 22832 38108
rect 22832 38052 22836 38108
rect 22772 38048 22836 38052
rect 22852 38108 22916 38112
rect 22852 38052 22856 38108
rect 22856 38052 22912 38108
rect 22912 38052 22916 38108
rect 22852 38048 22916 38052
rect 27612 38108 27676 38112
rect 27612 38052 27616 38108
rect 27616 38052 27672 38108
rect 27672 38052 27676 38108
rect 27612 38048 27676 38052
rect 27692 38108 27756 38112
rect 27692 38052 27696 38108
rect 27696 38052 27752 38108
rect 27752 38052 27756 38108
rect 27692 38048 27756 38052
rect 27772 38108 27836 38112
rect 27772 38052 27776 38108
rect 27776 38052 27832 38108
rect 27832 38052 27836 38108
rect 27772 38048 27836 38052
rect 27852 38108 27916 38112
rect 27852 38052 27856 38108
rect 27856 38052 27912 38108
rect 27912 38052 27916 38108
rect 27852 38048 27916 38052
rect 32612 38108 32676 38112
rect 32612 38052 32616 38108
rect 32616 38052 32672 38108
rect 32672 38052 32676 38108
rect 32612 38048 32676 38052
rect 32692 38108 32756 38112
rect 32692 38052 32696 38108
rect 32696 38052 32752 38108
rect 32752 38052 32756 38108
rect 32692 38048 32756 38052
rect 32772 38108 32836 38112
rect 32772 38052 32776 38108
rect 32776 38052 32832 38108
rect 32832 38052 32836 38108
rect 32772 38048 32836 38052
rect 32852 38108 32916 38112
rect 32852 38052 32856 38108
rect 32856 38052 32912 38108
rect 32912 38052 32916 38108
rect 32852 38048 32916 38052
rect 37612 38108 37676 38112
rect 37612 38052 37616 38108
rect 37616 38052 37672 38108
rect 37672 38052 37676 38108
rect 37612 38048 37676 38052
rect 37692 38108 37756 38112
rect 37692 38052 37696 38108
rect 37696 38052 37752 38108
rect 37752 38052 37756 38108
rect 37692 38048 37756 38052
rect 37772 38108 37836 38112
rect 37772 38052 37776 38108
rect 37776 38052 37832 38108
rect 37832 38052 37836 38108
rect 37772 38048 37836 38052
rect 37852 38108 37916 38112
rect 37852 38052 37856 38108
rect 37856 38052 37912 38108
rect 37912 38052 37916 38108
rect 37852 38048 37916 38052
rect 42612 38108 42676 38112
rect 42612 38052 42616 38108
rect 42616 38052 42672 38108
rect 42672 38052 42676 38108
rect 42612 38048 42676 38052
rect 42692 38108 42756 38112
rect 42692 38052 42696 38108
rect 42696 38052 42752 38108
rect 42752 38052 42756 38108
rect 42692 38048 42756 38052
rect 42772 38108 42836 38112
rect 42772 38052 42776 38108
rect 42776 38052 42832 38108
rect 42832 38052 42836 38108
rect 42772 38048 42836 38052
rect 42852 38108 42916 38112
rect 42852 38052 42856 38108
rect 42856 38052 42912 38108
rect 42912 38052 42916 38108
rect 42852 38048 42916 38052
rect 47612 38108 47676 38112
rect 47612 38052 47616 38108
rect 47616 38052 47672 38108
rect 47672 38052 47676 38108
rect 47612 38048 47676 38052
rect 47692 38108 47756 38112
rect 47692 38052 47696 38108
rect 47696 38052 47752 38108
rect 47752 38052 47756 38108
rect 47692 38048 47756 38052
rect 47772 38108 47836 38112
rect 47772 38052 47776 38108
rect 47776 38052 47832 38108
rect 47832 38052 47836 38108
rect 47772 38048 47836 38052
rect 47852 38108 47916 38112
rect 47852 38052 47856 38108
rect 47856 38052 47912 38108
rect 47912 38052 47916 38108
rect 47852 38048 47916 38052
rect 52612 38108 52676 38112
rect 52612 38052 52616 38108
rect 52616 38052 52672 38108
rect 52672 38052 52676 38108
rect 52612 38048 52676 38052
rect 52692 38108 52756 38112
rect 52692 38052 52696 38108
rect 52696 38052 52752 38108
rect 52752 38052 52756 38108
rect 52692 38048 52756 38052
rect 52772 38108 52836 38112
rect 52772 38052 52776 38108
rect 52776 38052 52832 38108
rect 52832 38052 52836 38108
rect 52772 38048 52836 38052
rect 52852 38108 52916 38112
rect 52852 38052 52856 38108
rect 52856 38052 52912 38108
rect 52912 38052 52916 38108
rect 52852 38048 52916 38052
rect 57612 38108 57676 38112
rect 57612 38052 57616 38108
rect 57616 38052 57672 38108
rect 57672 38052 57676 38108
rect 57612 38048 57676 38052
rect 57692 38108 57756 38112
rect 57692 38052 57696 38108
rect 57696 38052 57752 38108
rect 57752 38052 57756 38108
rect 57692 38048 57756 38052
rect 57772 38108 57836 38112
rect 57772 38052 57776 38108
rect 57776 38052 57832 38108
rect 57832 38052 57836 38108
rect 57772 38048 57836 38052
rect 57852 38108 57916 38112
rect 57852 38052 57856 38108
rect 57856 38052 57912 38108
rect 57912 38052 57916 38108
rect 57852 38048 57916 38052
rect 1952 37564 2016 37568
rect 1952 37508 1956 37564
rect 1956 37508 2012 37564
rect 2012 37508 2016 37564
rect 1952 37504 2016 37508
rect 2032 37564 2096 37568
rect 2032 37508 2036 37564
rect 2036 37508 2092 37564
rect 2092 37508 2096 37564
rect 2032 37504 2096 37508
rect 2112 37564 2176 37568
rect 2112 37508 2116 37564
rect 2116 37508 2172 37564
rect 2172 37508 2176 37564
rect 2112 37504 2176 37508
rect 2192 37564 2256 37568
rect 2192 37508 2196 37564
rect 2196 37508 2252 37564
rect 2252 37508 2256 37564
rect 2192 37504 2256 37508
rect 6952 37564 7016 37568
rect 6952 37508 6956 37564
rect 6956 37508 7012 37564
rect 7012 37508 7016 37564
rect 6952 37504 7016 37508
rect 7032 37564 7096 37568
rect 7032 37508 7036 37564
rect 7036 37508 7092 37564
rect 7092 37508 7096 37564
rect 7032 37504 7096 37508
rect 7112 37564 7176 37568
rect 7112 37508 7116 37564
rect 7116 37508 7172 37564
rect 7172 37508 7176 37564
rect 7112 37504 7176 37508
rect 7192 37564 7256 37568
rect 7192 37508 7196 37564
rect 7196 37508 7252 37564
rect 7252 37508 7256 37564
rect 7192 37504 7256 37508
rect 11952 37564 12016 37568
rect 11952 37508 11956 37564
rect 11956 37508 12012 37564
rect 12012 37508 12016 37564
rect 11952 37504 12016 37508
rect 12032 37564 12096 37568
rect 12032 37508 12036 37564
rect 12036 37508 12092 37564
rect 12092 37508 12096 37564
rect 12032 37504 12096 37508
rect 12112 37564 12176 37568
rect 12112 37508 12116 37564
rect 12116 37508 12172 37564
rect 12172 37508 12176 37564
rect 12112 37504 12176 37508
rect 12192 37564 12256 37568
rect 12192 37508 12196 37564
rect 12196 37508 12252 37564
rect 12252 37508 12256 37564
rect 12192 37504 12256 37508
rect 16952 37564 17016 37568
rect 16952 37508 16956 37564
rect 16956 37508 17012 37564
rect 17012 37508 17016 37564
rect 16952 37504 17016 37508
rect 17032 37564 17096 37568
rect 17032 37508 17036 37564
rect 17036 37508 17092 37564
rect 17092 37508 17096 37564
rect 17032 37504 17096 37508
rect 17112 37564 17176 37568
rect 17112 37508 17116 37564
rect 17116 37508 17172 37564
rect 17172 37508 17176 37564
rect 17112 37504 17176 37508
rect 17192 37564 17256 37568
rect 17192 37508 17196 37564
rect 17196 37508 17252 37564
rect 17252 37508 17256 37564
rect 17192 37504 17256 37508
rect 21952 37564 22016 37568
rect 21952 37508 21956 37564
rect 21956 37508 22012 37564
rect 22012 37508 22016 37564
rect 21952 37504 22016 37508
rect 22032 37564 22096 37568
rect 22032 37508 22036 37564
rect 22036 37508 22092 37564
rect 22092 37508 22096 37564
rect 22032 37504 22096 37508
rect 22112 37564 22176 37568
rect 22112 37508 22116 37564
rect 22116 37508 22172 37564
rect 22172 37508 22176 37564
rect 22112 37504 22176 37508
rect 22192 37564 22256 37568
rect 22192 37508 22196 37564
rect 22196 37508 22252 37564
rect 22252 37508 22256 37564
rect 22192 37504 22256 37508
rect 26952 37564 27016 37568
rect 26952 37508 26956 37564
rect 26956 37508 27012 37564
rect 27012 37508 27016 37564
rect 26952 37504 27016 37508
rect 27032 37564 27096 37568
rect 27032 37508 27036 37564
rect 27036 37508 27092 37564
rect 27092 37508 27096 37564
rect 27032 37504 27096 37508
rect 27112 37564 27176 37568
rect 27112 37508 27116 37564
rect 27116 37508 27172 37564
rect 27172 37508 27176 37564
rect 27112 37504 27176 37508
rect 27192 37564 27256 37568
rect 27192 37508 27196 37564
rect 27196 37508 27252 37564
rect 27252 37508 27256 37564
rect 27192 37504 27256 37508
rect 31952 37564 32016 37568
rect 31952 37508 31956 37564
rect 31956 37508 32012 37564
rect 32012 37508 32016 37564
rect 31952 37504 32016 37508
rect 32032 37564 32096 37568
rect 32032 37508 32036 37564
rect 32036 37508 32092 37564
rect 32092 37508 32096 37564
rect 32032 37504 32096 37508
rect 32112 37564 32176 37568
rect 32112 37508 32116 37564
rect 32116 37508 32172 37564
rect 32172 37508 32176 37564
rect 32112 37504 32176 37508
rect 32192 37564 32256 37568
rect 32192 37508 32196 37564
rect 32196 37508 32252 37564
rect 32252 37508 32256 37564
rect 32192 37504 32256 37508
rect 36952 37564 37016 37568
rect 36952 37508 36956 37564
rect 36956 37508 37012 37564
rect 37012 37508 37016 37564
rect 36952 37504 37016 37508
rect 37032 37564 37096 37568
rect 37032 37508 37036 37564
rect 37036 37508 37092 37564
rect 37092 37508 37096 37564
rect 37032 37504 37096 37508
rect 37112 37564 37176 37568
rect 37112 37508 37116 37564
rect 37116 37508 37172 37564
rect 37172 37508 37176 37564
rect 37112 37504 37176 37508
rect 37192 37564 37256 37568
rect 37192 37508 37196 37564
rect 37196 37508 37252 37564
rect 37252 37508 37256 37564
rect 37192 37504 37256 37508
rect 41952 37564 42016 37568
rect 41952 37508 41956 37564
rect 41956 37508 42012 37564
rect 42012 37508 42016 37564
rect 41952 37504 42016 37508
rect 42032 37564 42096 37568
rect 42032 37508 42036 37564
rect 42036 37508 42092 37564
rect 42092 37508 42096 37564
rect 42032 37504 42096 37508
rect 42112 37564 42176 37568
rect 42112 37508 42116 37564
rect 42116 37508 42172 37564
rect 42172 37508 42176 37564
rect 42112 37504 42176 37508
rect 42192 37564 42256 37568
rect 42192 37508 42196 37564
rect 42196 37508 42252 37564
rect 42252 37508 42256 37564
rect 42192 37504 42256 37508
rect 46952 37564 47016 37568
rect 46952 37508 46956 37564
rect 46956 37508 47012 37564
rect 47012 37508 47016 37564
rect 46952 37504 47016 37508
rect 47032 37564 47096 37568
rect 47032 37508 47036 37564
rect 47036 37508 47092 37564
rect 47092 37508 47096 37564
rect 47032 37504 47096 37508
rect 47112 37564 47176 37568
rect 47112 37508 47116 37564
rect 47116 37508 47172 37564
rect 47172 37508 47176 37564
rect 47112 37504 47176 37508
rect 47192 37564 47256 37568
rect 47192 37508 47196 37564
rect 47196 37508 47252 37564
rect 47252 37508 47256 37564
rect 47192 37504 47256 37508
rect 51952 37564 52016 37568
rect 51952 37508 51956 37564
rect 51956 37508 52012 37564
rect 52012 37508 52016 37564
rect 51952 37504 52016 37508
rect 52032 37564 52096 37568
rect 52032 37508 52036 37564
rect 52036 37508 52092 37564
rect 52092 37508 52096 37564
rect 52032 37504 52096 37508
rect 52112 37564 52176 37568
rect 52112 37508 52116 37564
rect 52116 37508 52172 37564
rect 52172 37508 52176 37564
rect 52112 37504 52176 37508
rect 52192 37564 52256 37568
rect 52192 37508 52196 37564
rect 52196 37508 52252 37564
rect 52252 37508 52256 37564
rect 52192 37504 52256 37508
rect 56952 37564 57016 37568
rect 56952 37508 56956 37564
rect 56956 37508 57012 37564
rect 57012 37508 57016 37564
rect 56952 37504 57016 37508
rect 57032 37564 57096 37568
rect 57032 37508 57036 37564
rect 57036 37508 57092 37564
rect 57092 37508 57096 37564
rect 57032 37504 57096 37508
rect 57112 37564 57176 37568
rect 57112 37508 57116 37564
rect 57116 37508 57172 37564
rect 57172 37508 57176 37564
rect 57112 37504 57176 37508
rect 57192 37564 57256 37568
rect 57192 37508 57196 37564
rect 57196 37508 57252 37564
rect 57252 37508 57256 37564
rect 57192 37504 57256 37508
rect 2612 37020 2676 37024
rect 2612 36964 2616 37020
rect 2616 36964 2672 37020
rect 2672 36964 2676 37020
rect 2612 36960 2676 36964
rect 2692 37020 2756 37024
rect 2692 36964 2696 37020
rect 2696 36964 2752 37020
rect 2752 36964 2756 37020
rect 2692 36960 2756 36964
rect 2772 37020 2836 37024
rect 2772 36964 2776 37020
rect 2776 36964 2832 37020
rect 2832 36964 2836 37020
rect 2772 36960 2836 36964
rect 2852 37020 2916 37024
rect 2852 36964 2856 37020
rect 2856 36964 2912 37020
rect 2912 36964 2916 37020
rect 2852 36960 2916 36964
rect 7612 37020 7676 37024
rect 7612 36964 7616 37020
rect 7616 36964 7672 37020
rect 7672 36964 7676 37020
rect 7612 36960 7676 36964
rect 7692 37020 7756 37024
rect 7692 36964 7696 37020
rect 7696 36964 7752 37020
rect 7752 36964 7756 37020
rect 7692 36960 7756 36964
rect 7772 37020 7836 37024
rect 7772 36964 7776 37020
rect 7776 36964 7832 37020
rect 7832 36964 7836 37020
rect 7772 36960 7836 36964
rect 7852 37020 7916 37024
rect 7852 36964 7856 37020
rect 7856 36964 7912 37020
rect 7912 36964 7916 37020
rect 7852 36960 7916 36964
rect 12612 37020 12676 37024
rect 12612 36964 12616 37020
rect 12616 36964 12672 37020
rect 12672 36964 12676 37020
rect 12612 36960 12676 36964
rect 12692 37020 12756 37024
rect 12692 36964 12696 37020
rect 12696 36964 12752 37020
rect 12752 36964 12756 37020
rect 12692 36960 12756 36964
rect 12772 37020 12836 37024
rect 12772 36964 12776 37020
rect 12776 36964 12832 37020
rect 12832 36964 12836 37020
rect 12772 36960 12836 36964
rect 12852 37020 12916 37024
rect 12852 36964 12856 37020
rect 12856 36964 12912 37020
rect 12912 36964 12916 37020
rect 12852 36960 12916 36964
rect 17612 37020 17676 37024
rect 17612 36964 17616 37020
rect 17616 36964 17672 37020
rect 17672 36964 17676 37020
rect 17612 36960 17676 36964
rect 17692 37020 17756 37024
rect 17692 36964 17696 37020
rect 17696 36964 17752 37020
rect 17752 36964 17756 37020
rect 17692 36960 17756 36964
rect 17772 37020 17836 37024
rect 17772 36964 17776 37020
rect 17776 36964 17832 37020
rect 17832 36964 17836 37020
rect 17772 36960 17836 36964
rect 17852 37020 17916 37024
rect 17852 36964 17856 37020
rect 17856 36964 17912 37020
rect 17912 36964 17916 37020
rect 17852 36960 17916 36964
rect 22612 37020 22676 37024
rect 22612 36964 22616 37020
rect 22616 36964 22672 37020
rect 22672 36964 22676 37020
rect 22612 36960 22676 36964
rect 22692 37020 22756 37024
rect 22692 36964 22696 37020
rect 22696 36964 22752 37020
rect 22752 36964 22756 37020
rect 22692 36960 22756 36964
rect 22772 37020 22836 37024
rect 22772 36964 22776 37020
rect 22776 36964 22832 37020
rect 22832 36964 22836 37020
rect 22772 36960 22836 36964
rect 22852 37020 22916 37024
rect 22852 36964 22856 37020
rect 22856 36964 22912 37020
rect 22912 36964 22916 37020
rect 22852 36960 22916 36964
rect 27612 37020 27676 37024
rect 27612 36964 27616 37020
rect 27616 36964 27672 37020
rect 27672 36964 27676 37020
rect 27612 36960 27676 36964
rect 27692 37020 27756 37024
rect 27692 36964 27696 37020
rect 27696 36964 27752 37020
rect 27752 36964 27756 37020
rect 27692 36960 27756 36964
rect 27772 37020 27836 37024
rect 27772 36964 27776 37020
rect 27776 36964 27832 37020
rect 27832 36964 27836 37020
rect 27772 36960 27836 36964
rect 27852 37020 27916 37024
rect 27852 36964 27856 37020
rect 27856 36964 27912 37020
rect 27912 36964 27916 37020
rect 27852 36960 27916 36964
rect 32612 37020 32676 37024
rect 32612 36964 32616 37020
rect 32616 36964 32672 37020
rect 32672 36964 32676 37020
rect 32612 36960 32676 36964
rect 32692 37020 32756 37024
rect 32692 36964 32696 37020
rect 32696 36964 32752 37020
rect 32752 36964 32756 37020
rect 32692 36960 32756 36964
rect 32772 37020 32836 37024
rect 32772 36964 32776 37020
rect 32776 36964 32832 37020
rect 32832 36964 32836 37020
rect 32772 36960 32836 36964
rect 32852 37020 32916 37024
rect 32852 36964 32856 37020
rect 32856 36964 32912 37020
rect 32912 36964 32916 37020
rect 32852 36960 32916 36964
rect 37612 37020 37676 37024
rect 37612 36964 37616 37020
rect 37616 36964 37672 37020
rect 37672 36964 37676 37020
rect 37612 36960 37676 36964
rect 37692 37020 37756 37024
rect 37692 36964 37696 37020
rect 37696 36964 37752 37020
rect 37752 36964 37756 37020
rect 37692 36960 37756 36964
rect 37772 37020 37836 37024
rect 37772 36964 37776 37020
rect 37776 36964 37832 37020
rect 37832 36964 37836 37020
rect 37772 36960 37836 36964
rect 37852 37020 37916 37024
rect 37852 36964 37856 37020
rect 37856 36964 37912 37020
rect 37912 36964 37916 37020
rect 37852 36960 37916 36964
rect 42612 37020 42676 37024
rect 42612 36964 42616 37020
rect 42616 36964 42672 37020
rect 42672 36964 42676 37020
rect 42612 36960 42676 36964
rect 42692 37020 42756 37024
rect 42692 36964 42696 37020
rect 42696 36964 42752 37020
rect 42752 36964 42756 37020
rect 42692 36960 42756 36964
rect 42772 37020 42836 37024
rect 42772 36964 42776 37020
rect 42776 36964 42832 37020
rect 42832 36964 42836 37020
rect 42772 36960 42836 36964
rect 42852 37020 42916 37024
rect 42852 36964 42856 37020
rect 42856 36964 42912 37020
rect 42912 36964 42916 37020
rect 42852 36960 42916 36964
rect 47612 37020 47676 37024
rect 47612 36964 47616 37020
rect 47616 36964 47672 37020
rect 47672 36964 47676 37020
rect 47612 36960 47676 36964
rect 47692 37020 47756 37024
rect 47692 36964 47696 37020
rect 47696 36964 47752 37020
rect 47752 36964 47756 37020
rect 47692 36960 47756 36964
rect 47772 37020 47836 37024
rect 47772 36964 47776 37020
rect 47776 36964 47832 37020
rect 47832 36964 47836 37020
rect 47772 36960 47836 36964
rect 47852 37020 47916 37024
rect 47852 36964 47856 37020
rect 47856 36964 47912 37020
rect 47912 36964 47916 37020
rect 47852 36960 47916 36964
rect 52612 37020 52676 37024
rect 52612 36964 52616 37020
rect 52616 36964 52672 37020
rect 52672 36964 52676 37020
rect 52612 36960 52676 36964
rect 52692 37020 52756 37024
rect 52692 36964 52696 37020
rect 52696 36964 52752 37020
rect 52752 36964 52756 37020
rect 52692 36960 52756 36964
rect 52772 37020 52836 37024
rect 52772 36964 52776 37020
rect 52776 36964 52832 37020
rect 52832 36964 52836 37020
rect 52772 36960 52836 36964
rect 52852 37020 52916 37024
rect 52852 36964 52856 37020
rect 52856 36964 52912 37020
rect 52912 36964 52916 37020
rect 52852 36960 52916 36964
rect 57612 37020 57676 37024
rect 57612 36964 57616 37020
rect 57616 36964 57672 37020
rect 57672 36964 57676 37020
rect 57612 36960 57676 36964
rect 57692 37020 57756 37024
rect 57692 36964 57696 37020
rect 57696 36964 57752 37020
rect 57752 36964 57756 37020
rect 57692 36960 57756 36964
rect 57772 37020 57836 37024
rect 57772 36964 57776 37020
rect 57776 36964 57832 37020
rect 57832 36964 57836 37020
rect 57772 36960 57836 36964
rect 57852 37020 57916 37024
rect 57852 36964 57856 37020
rect 57856 36964 57912 37020
rect 57912 36964 57916 37020
rect 57852 36960 57916 36964
rect 1952 36476 2016 36480
rect 1952 36420 1956 36476
rect 1956 36420 2012 36476
rect 2012 36420 2016 36476
rect 1952 36416 2016 36420
rect 2032 36476 2096 36480
rect 2032 36420 2036 36476
rect 2036 36420 2092 36476
rect 2092 36420 2096 36476
rect 2032 36416 2096 36420
rect 2112 36476 2176 36480
rect 2112 36420 2116 36476
rect 2116 36420 2172 36476
rect 2172 36420 2176 36476
rect 2112 36416 2176 36420
rect 2192 36476 2256 36480
rect 2192 36420 2196 36476
rect 2196 36420 2252 36476
rect 2252 36420 2256 36476
rect 2192 36416 2256 36420
rect 6952 36476 7016 36480
rect 6952 36420 6956 36476
rect 6956 36420 7012 36476
rect 7012 36420 7016 36476
rect 6952 36416 7016 36420
rect 7032 36476 7096 36480
rect 7032 36420 7036 36476
rect 7036 36420 7092 36476
rect 7092 36420 7096 36476
rect 7032 36416 7096 36420
rect 7112 36476 7176 36480
rect 7112 36420 7116 36476
rect 7116 36420 7172 36476
rect 7172 36420 7176 36476
rect 7112 36416 7176 36420
rect 7192 36476 7256 36480
rect 7192 36420 7196 36476
rect 7196 36420 7252 36476
rect 7252 36420 7256 36476
rect 7192 36416 7256 36420
rect 11952 36476 12016 36480
rect 11952 36420 11956 36476
rect 11956 36420 12012 36476
rect 12012 36420 12016 36476
rect 11952 36416 12016 36420
rect 12032 36476 12096 36480
rect 12032 36420 12036 36476
rect 12036 36420 12092 36476
rect 12092 36420 12096 36476
rect 12032 36416 12096 36420
rect 12112 36476 12176 36480
rect 12112 36420 12116 36476
rect 12116 36420 12172 36476
rect 12172 36420 12176 36476
rect 12112 36416 12176 36420
rect 12192 36476 12256 36480
rect 12192 36420 12196 36476
rect 12196 36420 12252 36476
rect 12252 36420 12256 36476
rect 12192 36416 12256 36420
rect 16952 36476 17016 36480
rect 16952 36420 16956 36476
rect 16956 36420 17012 36476
rect 17012 36420 17016 36476
rect 16952 36416 17016 36420
rect 17032 36476 17096 36480
rect 17032 36420 17036 36476
rect 17036 36420 17092 36476
rect 17092 36420 17096 36476
rect 17032 36416 17096 36420
rect 17112 36476 17176 36480
rect 17112 36420 17116 36476
rect 17116 36420 17172 36476
rect 17172 36420 17176 36476
rect 17112 36416 17176 36420
rect 17192 36476 17256 36480
rect 17192 36420 17196 36476
rect 17196 36420 17252 36476
rect 17252 36420 17256 36476
rect 17192 36416 17256 36420
rect 21952 36476 22016 36480
rect 21952 36420 21956 36476
rect 21956 36420 22012 36476
rect 22012 36420 22016 36476
rect 21952 36416 22016 36420
rect 22032 36476 22096 36480
rect 22032 36420 22036 36476
rect 22036 36420 22092 36476
rect 22092 36420 22096 36476
rect 22032 36416 22096 36420
rect 22112 36476 22176 36480
rect 22112 36420 22116 36476
rect 22116 36420 22172 36476
rect 22172 36420 22176 36476
rect 22112 36416 22176 36420
rect 22192 36476 22256 36480
rect 22192 36420 22196 36476
rect 22196 36420 22252 36476
rect 22252 36420 22256 36476
rect 22192 36416 22256 36420
rect 26952 36476 27016 36480
rect 26952 36420 26956 36476
rect 26956 36420 27012 36476
rect 27012 36420 27016 36476
rect 26952 36416 27016 36420
rect 27032 36476 27096 36480
rect 27032 36420 27036 36476
rect 27036 36420 27092 36476
rect 27092 36420 27096 36476
rect 27032 36416 27096 36420
rect 27112 36476 27176 36480
rect 27112 36420 27116 36476
rect 27116 36420 27172 36476
rect 27172 36420 27176 36476
rect 27112 36416 27176 36420
rect 27192 36476 27256 36480
rect 27192 36420 27196 36476
rect 27196 36420 27252 36476
rect 27252 36420 27256 36476
rect 27192 36416 27256 36420
rect 31952 36476 32016 36480
rect 31952 36420 31956 36476
rect 31956 36420 32012 36476
rect 32012 36420 32016 36476
rect 31952 36416 32016 36420
rect 32032 36476 32096 36480
rect 32032 36420 32036 36476
rect 32036 36420 32092 36476
rect 32092 36420 32096 36476
rect 32032 36416 32096 36420
rect 32112 36476 32176 36480
rect 32112 36420 32116 36476
rect 32116 36420 32172 36476
rect 32172 36420 32176 36476
rect 32112 36416 32176 36420
rect 32192 36476 32256 36480
rect 32192 36420 32196 36476
rect 32196 36420 32252 36476
rect 32252 36420 32256 36476
rect 32192 36416 32256 36420
rect 36952 36476 37016 36480
rect 36952 36420 36956 36476
rect 36956 36420 37012 36476
rect 37012 36420 37016 36476
rect 36952 36416 37016 36420
rect 37032 36476 37096 36480
rect 37032 36420 37036 36476
rect 37036 36420 37092 36476
rect 37092 36420 37096 36476
rect 37032 36416 37096 36420
rect 37112 36476 37176 36480
rect 37112 36420 37116 36476
rect 37116 36420 37172 36476
rect 37172 36420 37176 36476
rect 37112 36416 37176 36420
rect 37192 36476 37256 36480
rect 37192 36420 37196 36476
rect 37196 36420 37252 36476
rect 37252 36420 37256 36476
rect 37192 36416 37256 36420
rect 41952 36476 42016 36480
rect 41952 36420 41956 36476
rect 41956 36420 42012 36476
rect 42012 36420 42016 36476
rect 41952 36416 42016 36420
rect 42032 36476 42096 36480
rect 42032 36420 42036 36476
rect 42036 36420 42092 36476
rect 42092 36420 42096 36476
rect 42032 36416 42096 36420
rect 42112 36476 42176 36480
rect 42112 36420 42116 36476
rect 42116 36420 42172 36476
rect 42172 36420 42176 36476
rect 42112 36416 42176 36420
rect 42192 36476 42256 36480
rect 42192 36420 42196 36476
rect 42196 36420 42252 36476
rect 42252 36420 42256 36476
rect 42192 36416 42256 36420
rect 46952 36476 47016 36480
rect 46952 36420 46956 36476
rect 46956 36420 47012 36476
rect 47012 36420 47016 36476
rect 46952 36416 47016 36420
rect 47032 36476 47096 36480
rect 47032 36420 47036 36476
rect 47036 36420 47092 36476
rect 47092 36420 47096 36476
rect 47032 36416 47096 36420
rect 47112 36476 47176 36480
rect 47112 36420 47116 36476
rect 47116 36420 47172 36476
rect 47172 36420 47176 36476
rect 47112 36416 47176 36420
rect 47192 36476 47256 36480
rect 47192 36420 47196 36476
rect 47196 36420 47252 36476
rect 47252 36420 47256 36476
rect 47192 36416 47256 36420
rect 51952 36476 52016 36480
rect 51952 36420 51956 36476
rect 51956 36420 52012 36476
rect 52012 36420 52016 36476
rect 51952 36416 52016 36420
rect 52032 36476 52096 36480
rect 52032 36420 52036 36476
rect 52036 36420 52092 36476
rect 52092 36420 52096 36476
rect 52032 36416 52096 36420
rect 52112 36476 52176 36480
rect 52112 36420 52116 36476
rect 52116 36420 52172 36476
rect 52172 36420 52176 36476
rect 52112 36416 52176 36420
rect 52192 36476 52256 36480
rect 52192 36420 52196 36476
rect 52196 36420 52252 36476
rect 52252 36420 52256 36476
rect 52192 36416 52256 36420
rect 56952 36476 57016 36480
rect 56952 36420 56956 36476
rect 56956 36420 57012 36476
rect 57012 36420 57016 36476
rect 56952 36416 57016 36420
rect 57032 36476 57096 36480
rect 57032 36420 57036 36476
rect 57036 36420 57092 36476
rect 57092 36420 57096 36476
rect 57032 36416 57096 36420
rect 57112 36476 57176 36480
rect 57112 36420 57116 36476
rect 57116 36420 57172 36476
rect 57172 36420 57176 36476
rect 57112 36416 57176 36420
rect 57192 36476 57256 36480
rect 57192 36420 57196 36476
rect 57196 36420 57252 36476
rect 57252 36420 57256 36476
rect 57192 36416 57256 36420
rect 2612 35932 2676 35936
rect 2612 35876 2616 35932
rect 2616 35876 2672 35932
rect 2672 35876 2676 35932
rect 2612 35872 2676 35876
rect 2692 35932 2756 35936
rect 2692 35876 2696 35932
rect 2696 35876 2752 35932
rect 2752 35876 2756 35932
rect 2692 35872 2756 35876
rect 2772 35932 2836 35936
rect 2772 35876 2776 35932
rect 2776 35876 2832 35932
rect 2832 35876 2836 35932
rect 2772 35872 2836 35876
rect 2852 35932 2916 35936
rect 2852 35876 2856 35932
rect 2856 35876 2912 35932
rect 2912 35876 2916 35932
rect 2852 35872 2916 35876
rect 7612 35932 7676 35936
rect 7612 35876 7616 35932
rect 7616 35876 7672 35932
rect 7672 35876 7676 35932
rect 7612 35872 7676 35876
rect 7692 35932 7756 35936
rect 7692 35876 7696 35932
rect 7696 35876 7752 35932
rect 7752 35876 7756 35932
rect 7692 35872 7756 35876
rect 7772 35932 7836 35936
rect 7772 35876 7776 35932
rect 7776 35876 7832 35932
rect 7832 35876 7836 35932
rect 7772 35872 7836 35876
rect 7852 35932 7916 35936
rect 7852 35876 7856 35932
rect 7856 35876 7912 35932
rect 7912 35876 7916 35932
rect 7852 35872 7916 35876
rect 12612 35932 12676 35936
rect 12612 35876 12616 35932
rect 12616 35876 12672 35932
rect 12672 35876 12676 35932
rect 12612 35872 12676 35876
rect 12692 35932 12756 35936
rect 12692 35876 12696 35932
rect 12696 35876 12752 35932
rect 12752 35876 12756 35932
rect 12692 35872 12756 35876
rect 12772 35932 12836 35936
rect 12772 35876 12776 35932
rect 12776 35876 12832 35932
rect 12832 35876 12836 35932
rect 12772 35872 12836 35876
rect 12852 35932 12916 35936
rect 12852 35876 12856 35932
rect 12856 35876 12912 35932
rect 12912 35876 12916 35932
rect 12852 35872 12916 35876
rect 17612 35932 17676 35936
rect 17612 35876 17616 35932
rect 17616 35876 17672 35932
rect 17672 35876 17676 35932
rect 17612 35872 17676 35876
rect 17692 35932 17756 35936
rect 17692 35876 17696 35932
rect 17696 35876 17752 35932
rect 17752 35876 17756 35932
rect 17692 35872 17756 35876
rect 17772 35932 17836 35936
rect 17772 35876 17776 35932
rect 17776 35876 17832 35932
rect 17832 35876 17836 35932
rect 17772 35872 17836 35876
rect 17852 35932 17916 35936
rect 17852 35876 17856 35932
rect 17856 35876 17912 35932
rect 17912 35876 17916 35932
rect 17852 35872 17916 35876
rect 22612 35932 22676 35936
rect 22612 35876 22616 35932
rect 22616 35876 22672 35932
rect 22672 35876 22676 35932
rect 22612 35872 22676 35876
rect 22692 35932 22756 35936
rect 22692 35876 22696 35932
rect 22696 35876 22752 35932
rect 22752 35876 22756 35932
rect 22692 35872 22756 35876
rect 22772 35932 22836 35936
rect 22772 35876 22776 35932
rect 22776 35876 22832 35932
rect 22832 35876 22836 35932
rect 22772 35872 22836 35876
rect 22852 35932 22916 35936
rect 22852 35876 22856 35932
rect 22856 35876 22912 35932
rect 22912 35876 22916 35932
rect 22852 35872 22916 35876
rect 27612 35932 27676 35936
rect 27612 35876 27616 35932
rect 27616 35876 27672 35932
rect 27672 35876 27676 35932
rect 27612 35872 27676 35876
rect 27692 35932 27756 35936
rect 27692 35876 27696 35932
rect 27696 35876 27752 35932
rect 27752 35876 27756 35932
rect 27692 35872 27756 35876
rect 27772 35932 27836 35936
rect 27772 35876 27776 35932
rect 27776 35876 27832 35932
rect 27832 35876 27836 35932
rect 27772 35872 27836 35876
rect 27852 35932 27916 35936
rect 27852 35876 27856 35932
rect 27856 35876 27912 35932
rect 27912 35876 27916 35932
rect 27852 35872 27916 35876
rect 32612 35932 32676 35936
rect 32612 35876 32616 35932
rect 32616 35876 32672 35932
rect 32672 35876 32676 35932
rect 32612 35872 32676 35876
rect 32692 35932 32756 35936
rect 32692 35876 32696 35932
rect 32696 35876 32752 35932
rect 32752 35876 32756 35932
rect 32692 35872 32756 35876
rect 32772 35932 32836 35936
rect 32772 35876 32776 35932
rect 32776 35876 32832 35932
rect 32832 35876 32836 35932
rect 32772 35872 32836 35876
rect 32852 35932 32916 35936
rect 32852 35876 32856 35932
rect 32856 35876 32912 35932
rect 32912 35876 32916 35932
rect 32852 35872 32916 35876
rect 37612 35932 37676 35936
rect 37612 35876 37616 35932
rect 37616 35876 37672 35932
rect 37672 35876 37676 35932
rect 37612 35872 37676 35876
rect 37692 35932 37756 35936
rect 37692 35876 37696 35932
rect 37696 35876 37752 35932
rect 37752 35876 37756 35932
rect 37692 35872 37756 35876
rect 37772 35932 37836 35936
rect 37772 35876 37776 35932
rect 37776 35876 37832 35932
rect 37832 35876 37836 35932
rect 37772 35872 37836 35876
rect 37852 35932 37916 35936
rect 37852 35876 37856 35932
rect 37856 35876 37912 35932
rect 37912 35876 37916 35932
rect 37852 35872 37916 35876
rect 42612 35932 42676 35936
rect 42612 35876 42616 35932
rect 42616 35876 42672 35932
rect 42672 35876 42676 35932
rect 42612 35872 42676 35876
rect 42692 35932 42756 35936
rect 42692 35876 42696 35932
rect 42696 35876 42752 35932
rect 42752 35876 42756 35932
rect 42692 35872 42756 35876
rect 42772 35932 42836 35936
rect 42772 35876 42776 35932
rect 42776 35876 42832 35932
rect 42832 35876 42836 35932
rect 42772 35872 42836 35876
rect 42852 35932 42916 35936
rect 42852 35876 42856 35932
rect 42856 35876 42912 35932
rect 42912 35876 42916 35932
rect 42852 35872 42916 35876
rect 47612 35932 47676 35936
rect 47612 35876 47616 35932
rect 47616 35876 47672 35932
rect 47672 35876 47676 35932
rect 47612 35872 47676 35876
rect 47692 35932 47756 35936
rect 47692 35876 47696 35932
rect 47696 35876 47752 35932
rect 47752 35876 47756 35932
rect 47692 35872 47756 35876
rect 47772 35932 47836 35936
rect 47772 35876 47776 35932
rect 47776 35876 47832 35932
rect 47832 35876 47836 35932
rect 47772 35872 47836 35876
rect 47852 35932 47916 35936
rect 47852 35876 47856 35932
rect 47856 35876 47912 35932
rect 47912 35876 47916 35932
rect 47852 35872 47916 35876
rect 52612 35932 52676 35936
rect 52612 35876 52616 35932
rect 52616 35876 52672 35932
rect 52672 35876 52676 35932
rect 52612 35872 52676 35876
rect 52692 35932 52756 35936
rect 52692 35876 52696 35932
rect 52696 35876 52752 35932
rect 52752 35876 52756 35932
rect 52692 35872 52756 35876
rect 52772 35932 52836 35936
rect 52772 35876 52776 35932
rect 52776 35876 52832 35932
rect 52832 35876 52836 35932
rect 52772 35872 52836 35876
rect 52852 35932 52916 35936
rect 52852 35876 52856 35932
rect 52856 35876 52912 35932
rect 52912 35876 52916 35932
rect 52852 35872 52916 35876
rect 57612 35932 57676 35936
rect 57612 35876 57616 35932
rect 57616 35876 57672 35932
rect 57672 35876 57676 35932
rect 57612 35872 57676 35876
rect 57692 35932 57756 35936
rect 57692 35876 57696 35932
rect 57696 35876 57752 35932
rect 57752 35876 57756 35932
rect 57692 35872 57756 35876
rect 57772 35932 57836 35936
rect 57772 35876 57776 35932
rect 57776 35876 57832 35932
rect 57832 35876 57836 35932
rect 57772 35872 57836 35876
rect 57852 35932 57916 35936
rect 57852 35876 57856 35932
rect 57856 35876 57912 35932
rect 57912 35876 57916 35932
rect 57852 35872 57916 35876
rect 1952 35388 2016 35392
rect 1952 35332 1956 35388
rect 1956 35332 2012 35388
rect 2012 35332 2016 35388
rect 1952 35328 2016 35332
rect 2032 35388 2096 35392
rect 2032 35332 2036 35388
rect 2036 35332 2092 35388
rect 2092 35332 2096 35388
rect 2032 35328 2096 35332
rect 2112 35388 2176 35392
rect 2112 35332 2116 35388
rect 2116 35332 2172 35388
rect 2172 35332 2176 35388
rect 2112 35328 2176 35332
rect 2192 35388 2256 35392
rect 2192 35332 2196 35388
rect 2196 35332 2252 35388
rect 2252 35332 2256 35388
rect 2192 35328 2256 35332
rect 6952 35388 7016 35392
rect 6952 35332 6956 35388
rect 6956 35332 7012 35388
rect 7012 35332 7016 35388
rect 6952 35328 7016 35332
rect 7032 35388 7096 35392
rect 7032 35332 7036 35388
rect 7036 35332 7092 35388
rect 7092 35332 7096 35388
rect 7032 35328 7096 35332
rect 7112 35388 7176 35392
rect 7112 35332 7116 35388
rect 7116 35332 7172 35388
rect 7172 35332 7176 35388
rect 7112 35328 7176 35332
rect 7192 35388 7256 35392
rect 7192 35332 7196 35388
rect 7196 35332 7252 35388
rect 7252 35332 7256 35388
rect 7192 35328 7256 35332
rect 11952 35388 12016 35392
rect 11952 35332 11956 35388
rect 11956 35332 12012 35388
rect 12012 35332 12016 35388
rect 11952 35328 12016 35332
rect 12032 35388 12096 35392
rect 12032 35332 12036 35388
rect 12036 35332 12092 35388
rect 12092 35332 12096 35388
rect 12032 35328 12096 35332
rect 12112 35388 12176 35392
rect 12112 35332 12116 35388
rect 12116 35332 12172 35388
rect 12172 35332 12176 35388
rect 12112 35328 12176 35332
rect 12192 35388 12256 35392
rect 12192 35332 12196 35388
rect 12196 35332 12252 35388
rect 12252 35332 12256 35388
rect 12192 35328 12256 35332
rect 16952 35388 17016 35392
rect 16952 35332 16956 35388
rect 16956 35332 17012 35388
rect 17012 35332 17016 35388
rect 16952 35328 17016 35332
rect 17032 35388 17096 35392
rect 17032 35332 17036 35388
rect 17036 35332 17092 35388
rect 17092 35332 17096 35388
rect 17032 35328 17096 35332
rect 17112 35388 17176 35392
rect 17112 35332 17116 35388
rect 17116 35332 17172 35388
rect 17172 35332 17176 35388
rect 17112 35328 17176 35332
rect 17192 35388 17256 35392
rect 17192 35332 17196 35388
rect 17196 35332 17252 35388
rect 17252 35332 17256 35388
rect 17192 35328 17256 35332
rect 21952 35388 22016 35392
rect 21952 35332 21956 35388
rect 21956 35332 22012 35388
rect 22012 35332 22016 35388
rect 21952 35328 22016 35332
rect 22032 35388 22096 35392
rect 22032 35332 22036 35388
rect 22036 35332 22092 35388
rect 22092 35332 22096 35388
rect 22032 35328 22096 35332
rect 22112 35388 22176 35392
rect 22112 35332 22116 35388
rect 22116 35332 22172 35388
rect 22172 35332 22176 35388
rect 22112 35328 22176 35332
rect 22192 35388 22256 35392
rect 22192 35332 22196 35388
rect 22196 35332 22252 35388
rect 22252 35332 22256 35388
rect 22192 35328 22256 35332
rect 26952 35388 27016 35392
rect 26952 35332 26956 35388
rect 26956 35332 27012 35388
rect 27012 35332 27016 35388
rect 26952 35328 27016 35332
rect 27032 35388 27096 35392
rect 27032 35332 27036 35388
rect 27036 35332 27092 35388
rect 27092 35332 27096 35388
rect 27032 35328 27096 35332
rect 27112 35388 27176 35392
rect 27112 35332 27116 35388
rect 27116 35332 27172 35388
rect 27172 35332 27176 35388
rect 27112 35328 27176 35332
rect 27192 35388 27256 35392
rect 27192 35332 27196 35388
rect 27196 35332 27252 35388
rect 27252 35332 27256 35388
rect 27192 35328 27256 35332
rect 31952 35388 32016 35392
rect 31952 35332 31956 35388
rect 31956 35332 32012 35388
rect 32012 35332 32016 35388
rect 31952 35328 32016 35332
rect 32032 35388 32096 35392
rect 32032 35332 32036 35388
rect 32036 35332 32092 35388
rect 32092 35332 32096 35388
rect 32032 35328 32096 35332
rect 32112 35388 32176 35392
rect 32112 35332 32116 35388
rect 32116 35332 32172 35388
rect 32172 35332 32176 35388
rect 32112 35328 32176 35332
rect 32192 35388 32256 35392
rect 32192 35332 32196 35388
rect 32196 35332 32252 35388
rect 32252 35332 32256 35388
rect 32192 35328 32256 35332
rect 36952 35388 37016 35392
rect 36952 35332 36956 35388
rect 36956 35332 37012 35388
rect 37012 35332 37016 35388
rect 36952 35328 37016 35332
rect 37032 35388 37096 35392
rect 37032 35332 37036 35388
rect 37036 35332 37092 35388
rect 37092 35332 37096 35388
rect 37032 35328 37096 35332
rect 37112 35388 37176 35392
rect 37112 35332 37116 35388
rect 37116 35332 37172 35388
rect 37172 35332 37176 35388
rect 37112 35328 37176 35332
rect 37192 35388 37256 35392
rect 37192 35332 37196 35388
rect 37196 35332 37252 35388
rect 37252 35332 37256 35388
rect 37192 35328 37256 35332
rect 41952 35388 42016 35392
rect 41952 35332 41956 35388
rect 41956 35332 42012 35388
rect 42012 35332 42016 35388
rect 41952 35328 42016 35332
rect 42032 35388 42096 35392
rect 42032 35332 42036 35388
rect 42036 35332 42092 35388
rect 42092 35332 42096 35388
rect 42032 35328 42096 35332
rect 42112 35388 42176 35392
rect 42112 35332 42116 35388
rect 42116 35332 42172 35388
rect 42172 35332 42176 35388
rect 42112 35328 42176 35332
rect 42192 35388 42256 35392
rect 42192 35332 42196 35388
rect 42196 35332 42252 35388
rect 42252 35332 42256 35388
rect 42192 35328 42256 35332
rect 46952 35388 47016 35392
rect 46952 35332 46956 35388
rect 46956 35332 47012 35388
rect 47012 35332 47016 35388
rect 46952 35328 47016 35332
rect 47032 35388 47096 35392
rect 47032 35332 47036 35388
rect 47036 35332 47092 35388
rect 47092 35332 47096 35388
rect 47032 35328 47096 35332
rect 47112 35388 47176 35392
rect 47112 35332 47116 35388
rect 47116 35332 47172 35388
rect 47172 35332 47176 35388
rect 47112 35328 47176 35332
rect 47192 35388 47256 35392
rect 47192 35332 47196 35388
rect 47196 35332 47252 35388
rect 47252 35332 47256 35388
rect 47192 35328 47256 35332
rect 51952 35388 52016 35392
rect 51952 35332 51956 35388
rect 51956 35332 52012 35388
rect 52012 35332 52016 35388
rect 51952 35328 52016 35332
rect 52032 35388 52096 35392
rect 52032 35332 52036 35388
rect 52036 35332 52092 35388
rect 52092 35332 52096 35388
rect 52032 35328 52096 35332
rect 52112 35388 52176 35392
rect 52112 35332 52116 35388
rect 52116 35332 52172 35388
rect 52172 35332 52176 35388
rect 52112 35328 52176 35332
rect 52192 35388 52256 35392
rect 52192 35332 52196 35388
rect 52196 35332 52252 35388
rect 52252 35332 52256 35388
rect 52192 35328 52256 35332
rect 56952 35388 57016 35392
rect 56952 35332 56956 35388
rect 56956 35332 57012 35388
rect 57012 35332 57016 35388
rect 56952 35328 57016 35332
rect 57032 35388 57096 35392
rect 57032 35332 57036 35388
rect 57036 35332 57092 35388
rect 57092 35332 57096 35388
rect 57032 35328 57096 35332
rect 57112 35388 57176 35392
rect 57112 35332 57116 35388
rect 57116 35332 57172 35388
rect 57172 35332 57176 35388
rect 57112 35328 57176 35332
rect 57192 35388 57256 35392
rect 57192 35332 57196 35388
rect 57196 35332 57252 35388
rect 57252 35332 57256 35388
rect 57192 35328 57256 35332
rect 2612 34844 2676 34848
rect 2612 34788 2616 34844
rect 2616 34788 2672 34844
rect 2672 34788 2676 34844
rect 2612 34784 2676 34788
rect 2692 34844 2756 34848
rect 2692 34788 2696 34844
rect 2696 34788 2752 34844
rect 2752 34788 2756 34844
rect 2692 34784 2756 34788
rect 2772 34844 2836 34848
rect 2772 34788 2776 34844
rect 2776 34788 2832 34844
rect 2832 34788 2836 34844
rect 2772 34784 2836 34788
rect 2852 34844 2916 34848
rect 2852 34788 2856 34844
rect 2856 34788 2912 34844
rect 2912 34788 2916 34844
rect 2852 34784 2916 34788
rect 7612 34844 7676 34848
rect 7612 34788 7616 34844
rect 7616 34788 7672 34844
rect 7672 34788 7676 34844
rect 7612 34784 7676 34788
rect 7692 34844 7756 34848
rect 7692 34788 7696 34844
rect 7696 34788 7752 34844
rect 7752 34788 7756 34844
rect 7692 34784 7756 34788
rect 7772 34844 7836 34848
rect 7772 34788 7776 34844
rect 7776 34788 7832 34844
rect 7832 34788 7836 34844
rect 7772 34784 7836 34788
rect 7852 34844 7916 34848
rect 7852 34788 7856 34844
rect 7856 34788 7912 34844
rect 7912 34788 7916 34844
rect 7852 34784 7916 34788
rect 12612 34844 12676 34848
rect 12612 34788 12616 34844
rect 12616 34788 12672 34844
rect 12672 34788 12676 34844
rect 12612 34784 12676 34788
rect 12692 34844 12756 34848
rect 12692 34788 12696 34844
rect 12696 34788 12752 34844
rect 12752 34788 12756 34844
rect 12692 34784 12756 34788
rect 12772 34844 12836 34848
rect 12772 34788 12776 34844
rect 12776 34788 12832 34844
rect 12832 34788 12836 34844
rect 12772 34784 12836 34788
rect 12852 34844 12916 34848
rect 12852 34788 12856 34844
rect 12856 34788 12912 34844
rect 12912 34788 12916 34844
rect 12852 34784 12916 34788
rect 17612 34844 17676 34848
rect 17612 34788 17616 34844
rect 17616 34788 17672 34844
rect 17672 34788 17676 34844
rect 17612 34784 17676 34788
rect 17692 34844 17756 34848
rect 17692 34788 17696 34844
rect 17696 34788 17752 34844
rect 17752 34788 17756 34844
rect 17692 34784 17756 34788
rect 17772 34844 17836 34848
rect 17772 34788 17776 34844
rect 17776 34788 17832 34844
rect 17832 34788 17836 34844
rect 17772 34784 17836 34788
rect 17852 34844 17916 34848
rect 17852 34788 17856 34844
rect 17856 34788 17912 34844
rect 17912 34788 17916 34844
rect 17852 34784 17916 34788
rect 22612 34844 22676 34848
rect 22612 34788 22616 34844
rect 22616 34788 22672 34844
rect 22672 34788 22676 34844
rect 22612 34784 22676 34788
rect 22692 34844 22756 34848
rect 22692 34788 22696 34844
rect 22696 34788 22752 34844
rect 22752 34788 22756 34844
rect 22692 34784 22756 34788
rect 22772 34844 22836 34848
rect 22772 34788 22776 34844
rect 22776 34788 22832 34844
rect 22832 34788 22836 34844
rect 22772 34784 22836 34788
rect 22852 34844 22916 34848
rect 22852 34788 22856 34844
rect 22856 34788 22912 34844
rect 22912 34788 22916 34844
rect 22852 34784 22916 34788
rect 27612 34844 27676 34848
rect 27612 34788 27616 34844
rect 27616 34788 27672 34844
rect 27672 34788 27676 34844
rect 27612 34784 27676 34788
rect 27692 34844 27756 34848
rect 27692 34788 27696 34844
rect 27696 34788 27752 34844
rect 27752 34788 27756 34844
rect 27692 34784 27756 34788
rect 27772 34844 27836 34848
rect 27772 34788 27776 34844
rect 27776 34788 27832 34844
rect 27832 34788 27836 34844
rect 27772 34784 27836 34788
rect 27852 34844 27916 34848
rect 27852 34788 27856 34844
rect 27856 34788 27912 34844
rect 27912 34788 27916 34844
rect 27852 34784 27916 34788
rect 32612 34844 32676 34848
rect 32612 34788 32616 34844
rect 32616 34788 32672 34844
rect 32672 34788 32676 34844
rect 32612 34784 32676 34788
rect 32692 34844 32756 34848
rect 32692 34788 32696 34844
rect 32696 34788 32752 34844
rect 32752 34788 32756 34844
rect 32692 34784 32756 34788
rect 32772 34844 32836 34848
rect 32772 34788 32776 34844
rect 32776 34788 32832 34844
rect 32832 34788 32836 34844
rect 32772 34784 32836 34788
rect 32852 34844 32916 34848
rect 32852 34788 32856 34844
rect 32856 34788 32912 34844
rect 32912 34788 32916 34844
rect 32852 34784 32916 34788
rect 37612 34844 37676 34848
rect 37612 34788 37616 34844
rect 37616 34788 37672 34844
rect 37672 34788 37676 34844
rect 37612 34784 37676 34788
rect 37692 34844 37756 34848
rect 37692 34788 37696 34844
rect 37696 34788 37752 34844
rect 37752 34788 37756 34844
rect 37692 34784 37756 34788
rect 37772 34844 37836 34848
rect 37772 34788 37776 34844
rect 37776 34788 37832 34844
rect 37832 34788 37836 34844
rect 37772 34784 37836 34788
rect 37852 34844 37916 34848
rect 37852 34788 37856 34844
rect 37856 34788 37912 34844
rect 37912 34788 37916 34844
rect 37852 34784 37916 34788
rect 42612 34844 42676 34848
rect 42612 34788 42616 34844
rect 42616 34788 42672 34844
rect 42672 34788 42676 34844
rect 42612 34784 42676 34788
rect 42692 34844 42756 34848
rect 42692 34788 42696 34844
rect 42696 34788 42752 34844
rect 42752 34788 42756 34844
rect 42692 34784 42756 34788
rect 42772 34844 42836 34848
rect 42772 34788 42776 34844
rect 42776 34788 42832 34844
rect 42832 34788 42836 34844
rect 42772 34784 42836 34788
rect 42852 34844 42916 34848
rect 42852 34788 42856 34844
rect 42856 34788 42912 34844
rect 42912 34788 42916 34844
rect 42852 34784 42916 34788
rect 47612 34844 47676 34848
rect 47612 34788 47616 34844
rect 47616 34788 47672 34844
rect 47672 34788 47676 34844
rect 47612 34784 47676 34788
rect 47692 34844 47756 34848
rect 47692 34788 47696 34844
rect 47696 34788 47752 34844
rect 47752 34788 47756 34844
rect 47692 34784 47756 34788
rect 47772 34844 47836 34848
rect 47772 34788 47776 34844
rect 47776 34788 47832 34844
rect 47832 34788 47836 34844
rect 47772 34784 47836 34788
rect 47852 34844 47916 34848
rect 47852 34788 47856 34844
rect 47856 34788 47912 34844
rect 47912 34788 47916 34844
rect 47852 34784 47916 34788
rect 52612 34844 52676 34848
rect 52612 34788 52616 34844
rect 52616 34788 52672 34844
rect 52672 34788 52676 34844
rect 52612 34784 52676 34788
rect 52692 34844 52756 34848
rect 52692 34788 52696 34844
rect 52696 34788 52752 34844
rect 52752 34788 52756 34844
rect 52692 34784 52756 34788
rect 52772 34844 52836 34848
rect 52772 34788 52776 34844
rect 52776 34788 52832 34844
rect 52832 34788 52836 34844
rect 52772 34784 52836 34788
rect 52852 34844 52916 34848
rect 52852 34788 52856 34844
rect 52856 34788 52912 34844
rect 52912 34788 52916 34844
rect 52852 34784 52916 34788
rect 57612 34844 57676 34848
rect 57612 34788 57616 34844
rect 57616 34788 57672 34844
rect 57672 34788 57676 34844
rect 57612 34784 57676 34788
rect 57692 34844 57756 34848
rect 57692 34788 57696 34844
rect 57696 34788 57752 34844
rect 57752 34788 57756 34844
rect 57692 34784 57756 34788
rect 57772 34844 57836 34848
rect 57772 34788 57776 34844
rect 57776 34788 57832 34844
rect 57832 34788 57836 34844
rect 57772 34784 57836 34788
rect 57852 34844 57916 34848
rect 57852 34788 57856 34844
rect 57856 34788 57912 34844
rect 57912 34788 57916 34844
rect 57852 34784 57916 34788
rect 1952 34300 2016 34304
rect 1952 34244 1956 34300
rect 1956 34244 2012 34300
rect 2012 34244 2016 34300
rect 1952 34240 2016 34244
rect 2032 34300 2096 34304
rect 2032 34244 2036 34300
rect 2036 34244 2092 34300
rect 2092 34244 2096 34300
rect 2032 34240 2096 34244
rect 2112 34300 2176 34304
rect 2112 34244 2116 34300
rect 2116 34244 2172 34300
rect 2172 34244 2176 34300
rect 2112 34240 2176 34244
rect 2192 34300 2256 34304
rect 2192 34244 2196 34300
rect 2196 34244 2252 34300
rect 2252 34244 2256 34300
rect 2192 34240 2256 34244
rect 6952 34300 7016 34304
rect 6952 34244 6956 34300
rect 6956 34244 7012 34300
rect 7012 34244 7016 34300
rect 6952 34240 7016 34244
rect 7032 34300 7096 34304
rect 7032 34244 7036 34300
rect 7036 34244 7092 34300
rect 7092 34244 7096 34300
rect 7032 34240 7096 34244
rect 7112 34300 7176 34304
rect 7112 34244 7116 34300
rect 7116 34244 7172 34300
rect 7172 34244 7176 34300
rect 7112 34240 7176 34244
rect 7192 34300 7256 34304
rect 7192 34244 7196 34300
rect 7196 34244 7252 34300
rect 7252 34244 7256 34300
rect 7192 34240 7256 34244
rect 11952 34300 12016 34304
rect 11952 34244 11956 34300
rect 11956 34244 12012 34300
rect 12012 34244 12016 34300
rect 11952 34240 12016 34244
rect 12032 34300 12096 34304
rect 12032 34244 12036 34300
rect 12036 34244 12092 34300
rect 12092 34244 12096 34300
rect 12032 34240 12096 34244
rect 12112 34300 12176 34304
rect 12112 34244 12116 34300
rect 12116 34244 12172 34300
rect 12172 34244 12176 34300
rect 12112 34240 12176 34244
rect 12192 34300 12256 34304
rect 12192 34244 12196 34300
rect 12196 34244 12252 34300
rect 12252 34244 12256 34300
rect 12192 34240 12256 34244
rect 16952 34300 17016 34304
rect 16952 34244 16956 34300
rect 16956 34244 17012 34300
rect 17012 34244 17016 34300
rect 16952 34240 17016 34244
rect 17032 34300 17096 34304
rect 17032 34244 17036 34300
rect 17036 34244 17092 34300
rect 17092 34244 17096 34300
rect 17032 34240 17096 34244
rect 17112 34300 17176 34304
rect 17112 34244 17116 34300
rect 17116 34244 17172 34300
rect 17172 34244 17176 34300
rect 17112 34240 17176 34244
rect 17192 34300 17256 34304
rect 17192 34244 17196 34300
rect 17196 34244 17252 34300
rect 17252 34244 17256 34300
rect 17192 34240 17256 34244
rect 21952 34300 22016 34304
rect 21952 34244 21956 34300
rect 21956 34244 22012 34300
rect 22012 34244 22016 34300
rect 21952 34240 22016 34244
rect 22032 34300 22096 34304
rect 22032 34244 22036 34300
rect 22036 34244 22092 34300
rect 22092 34244 22096 34300
rect 22032 34240 22096 34244
rect 22112 34300 22176 34304
rect 22112 34244 22116 34300
rect 22116 34244 22172 34300
rect 22172 34244 22176 34300
rect 22112 34240 22176 34244
rect 22192 34300 22256 34304
rect 22192 34244 22196 34300
rect 22196 34244 22252 34300
rect 22252 34244 22256 34300
rect 22192 34240 22256 34244
rect 26952 34300 27016 34304
rect 26952 34244 26956 34300
rect 26956 34244 27012 34300
rect 27012 34244 27016 34300
rect 26952 34240 27016 34244
rect 27032 34300 27096 34304
rect 27032 34244 27036 34300
rect 27036 34244 27092 34300
rect 27092 34244 27096 34300
rect 27032 34240 27096 34244
rect 27112 34300 27176 34304
rect 27112 34244 27116 34300
rect 27116 34244 27172 34300
rect 27172 34244 27176 34300
rect 27112 34240 27176 34244
rect 27192 34300 27256 34304
rect 27192 34244 27196 34300
rect 27196 34244 27252 34300
rect 27252 34244 27256 34300
rect 27192 34240 27256 34244
rect 31952 34300 32016 34304
rect 31952 34244 31956 34300
rect 31956 34244 32012 34300
rect 32012 34244 32016 34300
rect 31952 34240 32016 34244
rect 32032 34300 32096 34304
rect 32032 34244 32036 34300
rect 32036 34244 32092 34300
rect 32092 34244 32096 34300
rect 32032 34240 32096 34244
rect 32112 34300 32176 34304
rect 32112 34244 32116 34300
rect 32116 34244 32172 34300
rect 32172 34244 32176 34300
rect 32112 34240 32176 34244
rect 32192 34300 32256 34304
rect 32192 34244 32196 34300
rect 32196 34244 32252 34300
rect 32252 34244 32256 34300
rect 32192 34240 32256 34244
rect 36952 34300 37016 34304
rect 36952 34244 36956 34300
rect 36956 34244 37012 34300
rect 37012 34244 37016 34300
rect 36952 34240 37016 34244
rect 37032 34300 37096 34304
rect 37032 34244 37036 34300
rect 37036 34244 37092 34300
rect 37092 34244 37096 34300
rect 37032 34240 37096 34244
rect 37112 34300 37176 34304
rect 37112 34244 37116 34300
rect 37116 34244 37172 34300
rect 37172 34244 37176 34300
rect 37112 34240 37176 34244
rect 37192 34300 37256 34304
rect 37192 34244 37196 34300
rect 37196 34244 37252 34300
rect 37252 34244 37256 34300
rect 37192 34240 37256 34244
rect 41952 34300 42016 34304
rect 41952 34244 41956 34300
rect 41956 34244 42012 34300
rect 42012 34244 42016 34300
rect 41952 34240 42016 34244
rect 42032 34300 42096 34304
rect 42032 34244 42036 34300
rect 42036 34244 42092 34300
rect 42092 34244 42096 34300
rect 42032 34240 42096 34244
rect 42112 34300 42176 34304
rect 42112 34244 42116 34300
rect 42116 34244 42172 34300
rect 42172 34244 42176 34300
rect 42112 34240 42176 34244
rect 42192 34300 42256 34304
rect 42192 34244 42196 34300
rect 42196 34244 42252 34300
rect 42252 34244 42256 34300
rect 42192 34240 42256 34244
rect 46952 34300 47016 34304
rect 46952 34244 46956 34300
rect 46956 34244 47012 34300
rect 47012 34244 47016 34300
rect 46952 34240 47016 34244
rect 47032 34300 47096 34304
rect 47032 34244 47036 34300
rect 47036 34244 47092 34300
rect 47092 34244 47096 34300
rect 47032 34240 47096 34244
rect 47112 34300 47176 34304
rect 47112 34244 47116 34300
rect 47116 34244 47172 34300
rect 47172 34244 47176 34300
rect 47112 34240 47176 34244
rect 47192 34300 47256 34304
rect 47192 34244 47196 34300
rect 47196 34244 47252 34300
rect 47252 34244 47256 34300
rect 47192 34240 47256 34244
rect 51952 34300 52016 34304
rect 51952 34244 51956 34300
rect 51956 34244 52012 34300
rect 52012 34244 52016 34300
rect 51952 34240 52016 34244
rect 52032 34300 52096 34304
rect 52032 34244 52036 34300
rect 52036 34244 52092 34300
rect 52092 34244 52096 34300
rect 52032 34240 52096 34244
rect 52112 34300 52176 34304
rect 52112 34244 52116 34300
rect 52116 34244 52172 34300
rect 52172 34244 52176 34300
rect 52112 34240 52176 34244
rect 52192 34300 52256 34304
rect 52192 34244 52196 34300
rect 52196 34244 52252 34300
rect 52252 34244 52256 34300
rect 52192 34240 52256 34244
rect 56952 34300 57016 34304
rect 56952 34244 56956 34300
rect 56956 34244 57012 34300
rect 57012 34244 57016 34300
rect 56952 34240 57016 34244
rect 57032 34300 57096 34304
rect 57032 34244 57036 34300
rect 57036 34244 57092 34300
rect 57092 34244 57096 34300
rect 57032 34240 57096 34244
rect 57112 34300 57176 34304
rect 57112 34244 57116 34300
rect 57116 34244 57172 34300
rect 57172 34244 57176 34300
rect 57112 34240 57176 34244
rect 57192 34300 57256 34304
rect 57192 34244 57196 34300
rect 57196 34244 57252 34300
rect 57252 34244 57256 34300
rect 57192 34240 57256 34244
rect 2612 33756 2676 33760
rect 2612 33700 2616 33756
rect 2616 33700 2672 33756
rect 2672 33700 2676 33756
rect 2612 33696 2676 33700
rect 2692 33756 2756 33760
rect 2692 33700 2696 33756
rect 2696 33700 2752 33756
rect 2752 33700 2756 33756
rect 2692 33696 2756 33700
rect 2772 33756 2836 33760
rect 2772 33700 2776 33756
rect 2776 33700 2832 33756
rect 2832 33700 2836 33756
rect 2772 33696 2836 33700
rect 2852 33756 2916 33760
rect 2852 33700 2856 33756
rect 2856 33700 2912 33756
rect 2912 33700 2916 33756
rect 2852 33696 2916 33700
rect 7612 33756 7676 33760
rect 7612 33700 7616 33756
rect 7616 33700 7672 33756
rect 7672 33700 7676 33756
rect 7612 33696 7676 33700
rect 7692 33756 7756 33760
rect 7692 33700 7696 33756
rect 7696 33700 7752 33756
rect 7752 33700 7756 33756
rect 7692 33696 7756 33700
rect 7772 33756 7836 33760
rect 7772 33700 7776 33756
rect 7776 33700 7832 33756
rect 7832 33700 7836 33756
rect 7772 33696 7836 33700
rect 7852 33756 7916 33760
rect 7852 33700 7856 33756
rect 7856 33700 7912 33756
rect 7912 33700 7916 33756
rect 7852 33696 7916 33700
rect 12612 33756 12676 33760
rect 12612 33700 12616 33756
rect 12616 33700 12672 33756
rect 12672 33700 12676 33756
rect 12612 33696 12676 33700
rect 12692 33756 12756 33760
rect 12692 33700 12696 33756
rect 12696 33700 12752 33756
rect 12752 33700 12756 33756
rect 12692 33696 12756 33700
rect 12772 33756 12836 33760
rect 12772 33700 12776 33756
rect 12776 33700 12832 33756
rect 12832 33700 12836 33756
rect 12772 33696 12836 33700
rect 12852 33756 12916 33760
rect 12852 33700 12856 33756
rect 12856 33700 12912 33756
rect 12912 33700 12916 33756
rect 12852 33696 12916 33700
rect 17612 33756 17676 33760
rect 17612 33700 17616 33756
rect 17616 33700 17672 33756
rect 17672 33700 17676 33756
rect 17612 33696 17676 33700
rect 17692 33756 17756 33760
rect 17692 33700 17696 33756
rect 17696 33700 17752 33756
rect 17752 33700 17756 33756
rect 17692 33696 17756 33700
rect 17772 33756 17836 33760
rect 17772 33700 17776 33756
rect 17776 33700 17832 33756
rect 17832 33700 17836 33756
rect 17772 33696 17836 33700
rect 17852 33756 17916 33760
rect 17852 33700 17856 33756
rect 17856 33700 17912 33756
rect 17912 33700 17916 33756
rect 17852 33696 17916 33700
rect 22612 33756 22676 33760
rect 22612 33700 22616 33756
rect 22616 33700 22672 33756
rect 22672 33700 22676 33756
rect 22612 33696 22676 33700
rect 22692 33756 22756 33760
rect 22692 33700 22696 33756
rect 22696 33700 22752 33756
rect 22752 33700 22756 33756
rect 22692 33696 22756 33700
rect 22772 33756 22836 33760
rect 22772 33700 22776 33756
rect 22776 33700 22832 33756
rect 22832 33700 22836 33756
rect 22772 33696 22836 33700
rect 22852 33756 22916 33760
rect 22852 33700 22856 33756
rect 22856 33700 22912 33756
rect 22912 33700 22916 33756
rect 22852 33696 22916 33700
rect 27612 33756 27676 33760
rect 27612 33700 27616 33756
rect 27616 33700 27672 33756
rect 27672 33700 27676 33756
rect 27612 33696 27676 33700
rect 27692 33756 27756 33760
rect 27692 33700 27696 33756
rect 27696 33700 27752 33756
rect 27752 33700 27756 33756
rect 27692 33696 27756 33700
rect 27772 33756 27836 33760
rect 27772 33700 27776 33756
rect 27776 33700 27832 33756
rect 27832 33700 27836 33756
rect 27772 33696 27836 33700
rect 27852 33756 27916 33760
rect 27852 33700 27856 33756
rect 27856 33700 27912 33756
rect 27912 33700 27916 33756
rect 27852 33696 27916 33700
rect 32612 33756 32676 33760
rect 32612 33700 32616 33756
rect 32616 33700 32672 33756
rect 32672 33700 32676 33756
rect 32612 33696 32676 33700
rect 32692 33756 32756 33760
rect 32692 33700 32696 33756
rect 32696 33700 32752 33756
rect 32752 33700 32756 33756
rect 32692 33696 32756 33700
rect 32772 33756 32836 33760
rect 32772 33700 32776 33756
rect 32776 33700 32832 33756
rect 32832 33700 32836 33756
rect 32772 33696 32836 33700
rect 32852 33756 32916 33760
rect 32852 33700 32856 33756
rect 32856 33700 32912 33756
rect 32912 33700 32916 33756
rect 32852 33696 32916 33700
rect 37612 33756 37676 33760
rect 37612 33700 37616 33756
rect 37616 33700 37672 33756
rect 37672 33700 37676 33756
rect 37612 33696 37676 33700
rect 37692 33756 37756 33760
rect 37692 33700 37696 33756
rect 37696 33700 37752 33756
rect 37752 33700 37756 33756
rect 37692 33696 37756 33700
rect 37772 33756 37836 33760
rect 37772 33700 37776 33756
rect 37776 33700 37832 33756
rect 37832 33700 37836 33756
rect 37772 33696 37836 33700
rect 37852 33756 37916 33760
rect 37852 33700 37856 33756
rect 37856 33700 37912 33756
rect 37912 33700 37916 33756
rect 37852 33696 37916 33700
rect 42612 33756 42676 33760
rect 42612 33700 42616 33756
rect 42616 33700 42672 33756
rect 42672 33700 42676 33756
rect 42612 33696 42676 33700
rect 42692 33756 42756 33760
rect 42692 33700 42696 33756
rect 42696 33700 42752 33756
rect 42752 33700 42756 33756
rect 42692 33696 42756 33700
rect 42772 33756 42836 33760
rect 42772 33700 42776 33756
rect 42776 33700 42832 33756
rect 42832 33700 42836 33756
rect 42772 33696 42836 33700
rect 42852 33756 42916 33760
rect 42852 33700 42856 33756
rect 42856 33700 42912 33756
rect 42912 33700 42916 33756
rect 42852 33696 42916 33700
rect 47612 33756 47676 33760
rect 47612 33700 47616 33756
rect 47616 33700 47672 33756
rect 47672 33700 47676 33756
rect 47612 33696 47676 33700
rect 47692 33756 47756 33760
rect 47692 33700 47696 33756
rect 47696 33700 47752 33756
rect 47752 33700 47756 33756
rect 47692 33696 47756 33700
rect 47772 33756 47836 33760
rect 47772 33700 47776 33756
rect 47776 33700 47832 33756
rect 47832 33700 47836 33756
rect 47772 33696 47836 33700
rect 47852 33756 47916 33760
rect 47852 33700 47856 33756
rect 47856 33700 47912 33756
rect 47912 33700 47916 33756
rect 47852 33696 47916 33700
rect 52612 33756 52676 33760
rect 52612 33700 52616 33756
rect 52616 33700 52672 33756
rect 52672 33700 52676 33756
rect 52612 33696 52676 33700
rect 52692 33756 52756 33760
rect 52692 33700 52696 33756
rect 52696 33700 52752 33756
rect 52752 33700 52756 33756
rect 52692 33696 52756 33700
rect 52772 33756 52836 33760
rect 52772 33700 52776 33756
rect 52776 33700 52832 33756
rect 52832 33700 52836 33756
rect 52772 33696 52836 33700
rect 52852 33756 52916 33760
rect 52852 33700 52856 33756
rect 52856 33700 52912 33756
rect 52912 33700 52916 33756
rect 52852 33696 52916 33700
rect 57612 33756 57676 33760
rect 57612 33700 57616 33756
rect 57616 33700 57672 33756
rect 57672 33700 57676 33756
rect 57612 33696 57676 33700
rect 57692 33756 57756 33760
rect 57692 33700 57696 33756
rect 57696 33700 57752 33756
rect 57752 33700 57756 33756
rect 57692 33696 57756 33700
rect 57772 33756 57836 33760
rect 57772 33700 57776 33756
rect 57776 33700 57832 33756
rect 57832 33700 57836 33756
rect 57772 33696 57836 33700
rect 57852 33756 57916 33760
rect 57852 33700 57856 33756
rect 57856 33700 57912 33756
rect 57912 33700 57916 33756
rect 57852 33696 57916 33700
rect 1952 33212 2016 33216
rect 1952 33156 1956 33212
rect 1956 33156 2012 33212
rect 2012 33156 2016 33212
rect 1952 33152 2016 33156
rect 2032 33212 2096 33216
rect 2032 33156 2036 33212
rect 2036 33156 2092 33212
rect 2092 33156 2096 33212
rect 2032 33152 2096 33156
rect 2112 33212 2176 33216
rect 2112 33156 2116 33212
rect 2116 33156 2172 33212
rect 2172 33156 2176 33212
rect 2112 33152 2176 33156
rect 2192 33212 2256 33216
rect 2192 33156 2196 33212
rect 2196 33156 2252 33212
rect 2252 33156 2256 33212
rect 2192 33152 2256 33156
rect 6952 33212 7016 33216
rect 6952 33156 6956 33212
rect 6956 33156 7012 33212
rect 7012 33156 7016 33212
rect 6952 33152 7016 33156
rect 7032 33212 7096 33216
rect 7032 33156 7036 33212
rect 7036 33156 7092 33212
rect 7092 33156 7096 33212
rect 7032 33152 7096 33156
rect 7112 33212 7176 33216
rect 7112 33156 7116 33212
rect 7116 33156 7172 33212
rect 7172 33156 7176 33212
rect 7112 33152 7176 33156
rect 7192 33212 7256 33216
rect 7192 33156 7196 33212
rect 7196 33156 7252 33212
rect 7252 33156 7256 33212
rect 7192 33152 7256 33156
rect 11952 33212 12016 33216
rect 11952 33156 11956 33212
rect 11956 33156 12012 33212
rect 12012 33156 12016 33212
rect 11952 33152 12016 33156
rect 12032 33212 12096 33216
rect 12032 33156 12036 33212
rect 12036 33156 12092 33212
rect 12092 33156 12096 33212
rect 12032 33152 12096 33156
rect 12112 33212 12176 33216
rect 12112 33156 12116 33212
rect 12116 33156 12172 33212
rect 12172 33156 12176 33212
rect 12112 33152 12176 33156
rect 12192 33212 12256 33216
rect 12192 33156 12196 33212
rect 12196 33156 12252 33212
rect 12252 33156 12256 33212
rect 12192 33152 12256 33156
rect 16952 33212 17016 33216
rect 16952 33156 16956 33212
rect 16956 33156 17012 33212
rect 17012 33156 17016 33212
rect 16952 33152 17016 33156
rect 17032 33212 17096 33216
rect 17032 33156 17036 33212
rect 17036 33156 17092 33212
rect 17092 33156 17096 33212
rect 17032 33152 17096 33156
rect 17112 33212 17176 33216
rect 17112 33156 17116 33212
rect 17116 33156 17172 33212
rect 17172 33156 17176 33212
rect 17112 33152 17176 33156
rect 17192 33212 17256 33216
rect 17192 33156 17196 33212
rect 17196 33156 17252 33212
rect 17252 33156 17256 33212
rect 17192 33152 17256 33156
rect 21952 33212 22016 33216
rect 21952 33156 21956 33212
rect 21956 33156 22012 33212
rect 22012 33156 22016 33212
rect 21952 33152 22016 33156
rect 22032 33212 22096 33216
rect 22032 33156 22036 33212
rect 22036 33156 22092 33212
rect 22092 33156 22096 33212
rect 22032 33152 22096 33156
rect 22112 33212 22176 33216
rect 22112 33156 22116 33212
rect 22116 33156 22172 33212
rect 22172 33156 22176 33212
rect 22112 33152 22176 33156
rect 22192 33212 22256 33216
rect 22192 33156 22196 33212
rect 22196 33156 22252 33212
rect 22252 33156 22256 33212
rect 22192 33152 22256 33156
rect 26952 33212 27016 33216
rect 26952 33156 26956 33212
rect 26956 33156 27012 33212
rect 27012 33156 27016 33212
rect 26952 33152 27016 33156
rect 27032 33212 27096 33216
rect 27032 33156 27036 33212
rect 27036 33156 27092 33212
rect 27092 33156 27096 33212
rect 27032 33152 27096 33156
rect 27112 33212 27176 33216
rect 27112 33156 27116 33212
rect 27116 33156 27172 33212
rect 27172 33156 27176 33212
rect 27112 33152 27176 33156
rect 27192 33212 27256 33216
rect 27192 33156 27196 33212
rect 27196 33156 27252 33212
rect 27252 33156 27256 33212
rect 27192 33152 27256 33156
rect 31952 33212 32016 33216
rect 31952 33156 31956 33212
rect 31956 33156 32012 33212
rect 32012 33156 32016 33212
rect 31952 33152 32016 33156
rect 32032 33212 32096 33216
rect 32032 33156 32036 33212
rect 32036 33156 32092 33212
rect 32092 33156 32096 33212
rect 32032 33152 32096 33156
rect 32112 33212 32176 33216
rect 32112 33156 32116 33212
rect 32116 33156 32172 33212
rect 32172 33156 32176 33212
rect 32112 33152 32176 33156
rect 32192 33212 32256 33216
rect 32192 33156 32196 33212
rect 32196 33156 32252 33212
rect 32252 33156 32256 33212
rect 32192 33152 32256 33156
rect 36952 33212 37016 33216
rect 36952 33156 36956 33212
rect 36956 33156 37012 33212
rect 37012 33156 37016 33212
rect 36952 33152 37016 33156
rect 37032 33212 37096 33216
rect 37032 33156 37036 33212
rect 37036 33156 37092 33212
rect 37092 33156 37096 33212
rect 37032 33152 37096 33156
rect 37112 33212 37176 33216
rect 37112 33156 37116 33212
rect 37116 33156 37172 33212
rect 37172 33156 37176 33212
rect 37112 33152 37176 33156
rect 37192 33212 37256 33216
rect 37192 33156 37196 33212
rect 37196 33156 37252 33212
rect 37252 33156 37256 33212
rect 37192 33152 37256 33156
rect 41952 33212 42016 33216
rect 41952 33156 41956 33212
rect 41956 33156 42012 33212
rect 42012 33156 42016 33212
rect 41952 33152 42016 33156
rect 42032 33212 42096 33216
rect 42032 33156 42036 33212
rect 42036 33156 42092 33212
rect 42092 33156 42096 33212
rect 42032 33152 42096 33156
rect 42112 33212 42176 33216
rect 42112 33156 42116 33212
rect 42116 33156 42172 33212
rect 42172 33156 42176 33212
rect 42112 33152 42176 33156
rect 42192 33212 42256 33216
rect 42192 33156 42196 33212
rect 42196 33156 42252 33212
rect 42252 33156 42256 33212
rect 42192 33152 42256 33156
rect 46952 33212 47016 33216
rect 46952 33156 46956 33212
rect 46956 33156 47012 33212
rect 47012 33156 47016 33212
rect 46952 33152 47016 33156
rect 47032 33212 47096 33216
rect 47032 33156 47036 33212
rect 47036 33156 47092 33212
rect 47092 33156 47096 33212
rect 47032 33152 47096 33156
rect 47112 33212 47176 33216
rect 47112 33156 47116 33212
rect 47116 33156 47172 33212
rect 47172 33156 47176 33212
rect 47112 33152 47176 33156
rect 47192 33212 47256 33216
rect 47192 33156 47196 33212
rect 47196 33156 47252 33212
rect 47252 33156 47256 33212
rect 47192 33152 47256 33156
rect 51952 33212 52016 33216
rect 51952 33156 51956 33212
rect 51956 33156 52012 33212
rect 52012 33156 52016 33212
rect 51952 33152 52016 33156
rect 52032 33212 52096 33216
rect 52032 33156 52036 33212
rect 52036 33156 52092 33212
rect 52092 33156 52096 33212
rect 52032 33152 52096 33156
rect 52112 33212 52176 33216
rect 52112 33156 52116 33212
rect 52116 33156 52172 33212
rect 52172 33156 52176 33212
rect 52112 33152 52176 33156
rect 52192 33212 52256 33216
rect 52192 33156 52196 33212
rect 52196 33156 52252 33212
rect 52252 33156 52256 33212
rect 52192 33152 52256 33156
rect 56952 33212 57016 33216
rect 56952 33156 56956 33212
rect 56956 33156 57012 33212
rect 57012 33156 57016 33212
rect 56952 33152 57016 33156
rect 57032 33212 57096 33216
rect 57032 33156 57036 33212
rect 57036 33156 57092 33212
rect 57092 33156 57096 33212
rect 57032 33152 57096 33156
rect 57112 33212 57176 33216
rect 57112 33156 57116 33212
rect 57116 33156 57172 33212
rect 57172 33156 57176 33212
rect 57112 33152 57176 33156
rect 57192 33212 57256 33216
rect 57192 33156 57196 33212
rect 57196 33156 57252 33212
rect 57252 33156 57256 33212
rect 57192 33152 57256 33156
rect 2612 32668 2676 32672
rect 2612 32612 2616 32668
rect 2616 32612 2672 32668
rect 2672 32612 2676 32668
rect 2612 32608 2676 32612
rect 2692 32668 2756 32672
rect 2692 32612 2696 32668
rect 2696 32612 2752 32668
rect 2752 32612 2756 32668
rect 2692 32608 2756 32612
rect 2772 32668 2836 32672
rect 2772 32612 2776 32668
rect 2776 32612 2832 32668
rect 2832 32612 2836 32668
rect 2772 32608 2836 32612
rect 2852 32668 2916 32672
rect 2852 32612 2856 32668
rect 2856 32612 2912 32668
rect 2912 32612 2916 32668
rect 2852 32608 2916 32612
rect 7612 32668 7676 32672
rect 7612 32612 7616 32668
rect 7616 32612 7672 32668
rect 7672 32612 7676 32668
rect 7612 32608 7676 32612
rect 7692 32668 7756 32672
rect 7692 32612 7696 32668
rect 7696 32612 7752 32668
rect 7752 32612 7756 32668
rect 7692 32608 7756 32612
rect 7772 32668 7836 32672
rect 7772 32612 7776 32668
rect 7776 32612 7832 32668
rect 7832 32612 7836 32668
rect 7772 32608 7836 32612
rect 7852 32668 7916 32672
rect 7852 32612 7856 32668
rect 7856 32612 7912 32668
rect 7912 32612 7916 32668
rect 7852 32608 7916 32612
rect 12612 32668 12676 32672
rect 12612 32612 12616 32668
rect 12616 32612 12672 32668
rect 12672 32612 12676 32668
rect 12612 32608 12676 32612
rect 12692 32668 12756 32672
rect 12692 32612 12696 32668
rect 12696 32612 12752 32668
rect 12752 32612 12756 32668
rect 12692 32608 12756 32612
rect 12772 32668 12836 32672
rect 12772 32612 12776 32668
rect 12776 32612 12832 32668
rect 12832 32612 12836 32668
rect 12772 32608 12836 32612
rect 12852 32668 12916 32672
rect 12852 32612 12856 32668
rect 12856 32612 12912 32668
rect 12912 32612 12916 32668
rect 12852 32608 12916 32612
rect 17612 32668 17676 32672
rect 17612 32612 17616 32668
rect 17616 32612 17672 32668
rect 17672 32612 17676 32668
rect 17612 32608 17676 32612
rect 17692 32668 17756 32672
rect 17692 32612 17696 32668
rect 17696 32612 17752 32668
rect 17752 32612 17756 32668
rect 17692 32608 17756 32612
rect 17772 32668 17836 32672
rect 17772 32612 17776 32668
rect 17776 32612 17832 32668
rect 17832 32612 17836 32668
rect 17772 32608 17836 32612
rect 17852 32668 17916 32672
rect 17852 32612 17856 32668
rect 17856 32612 17912 32668
rect 17912 32612 17916 32668
rect 17852 32608 17916 32612
rect 22612 32668 22676 32672
rect 22612 32612 22616 32668
rect 22616 32612 22672 32668
rect 22672 32612 22676 32668
rect 22612 32608 22676 32612
rect 22692 32668 22756 32672
rect 22692 32612 22696 32668
rect 22696 32612 22752 32668
rect 22752 32612 22756 32668
rect 22692 32608 22756 32612
rect 22772 32668 22836 32672
rect 22772 32612 22776 32668
rect 22776 32612 22832 32668
rect 22832 32612 22836 32668
rect 22772 32608 22836 32612
rect 22852 32668 22916 32672
rect 22852 32612 22856 32668
rect 22856 32612 22912 32668
rect 22912 32612 22916 32668
rect 22852 32608 22916 32612
rect 27612 32668 27676 32672
rect 27612 32612 27616 32668
rect 27616 32612 27672 32668
rect 27672 32612 27676 32668
rect 27612 32608 27676 32612
rect 27692 32668 27756 32672
rect 27692 32612 27696 32668
rect 27696 32612 27752 32668
rect 27752 32612 27756 32668
rect 27692 32608 27756 32612
rect 27772 32668 27836 32672
rect 27772 32612 27776 32668
rect 27776 32612 27832 32668
rect 27832 32612 27836 32668
rect 27772 32608 27836 32612
rect 27852 32668 27916 32672
rect 27852 32612 27856 32668
rect 27856 32612 27912 32668
rect 27912 32612 27916 32668
rect 27852 32608 27916 32612
rect 32612 32668 32676 32672
rect 32612 32612 32616 32668
rect 32616 32612 32672 32668
rect 32672 32612 32676 32668
rect 32612 32608 32676 32612
rect 32692 32668 32756 32672
rect 32692 32612 32696 32668
rect 32696 32612 32752 32668
rect 32752 32612 32756 32668
rect 32692 32608 32756 32612
rect 32772 32668 32836 32672
rect 32772 32612 32776 32668
rect 32776 32612 32832 32668
rect 32832 32612 32836 32668
rect 32772 32608 32836 32612
rect 32852 32668 32916 32672
rect 32852 32612 32856 32668
rect 32856 32612 32912 32668
rect 32912 32612 32916 32668
rect 32852 32608 32916 32612
rect 37612 32668 37676 32672
rect 37612 32612 37616 32668
rect 37616 32612 37672 32668
rect 37672 32612 37676 32668
rect 37612 32608 37676 32612
rect 37692 32668 37756 32672
rect 37692 32612 37696 32668
rect 37696 32612 37752 32668
rect 37752 32612 37756 32668
rect 37692 32608 37756 32612
rect 37772 32668 37836 32672
rect 37772 32612 37776 32668
rect 37776 32612 37832 32668
rect 37832 32612 37836 32668
rect 37772 32608 37836 32612
rect 37852 32668 37916 32672
rect 37852 32612 37856 32668
rect 37856 32612 37912 32668
rect 37912 32612 37916 32668
rect 37852 32608 37916 32612
rect 42612 32668 42676 32672
rect 42612 32612 42616 32668
rect 42616 32612 42672 32668
rect 42672 32612 42676 32668
rect 42612 32608 42676 32612
rect 42692 32668 42756 32672
rect 42692 32612 42696 32668
rect 42696 32612 42752 32668
rect 42752 32612 42756 32668
rect 42692 32608 42756 32612
rect 42772 32668 42836 32672
rect 42772 32612 42776 32668
rect 42776 32612 42832 32668
rect 42832 32612 42836 32668
rect 42772 32608 42836 32612
rect 42852 32668 42916 32672
rect 42852 32612 42856 32668
rect 42856 32612 42912 32668
rect 42912 32612 42916 32668
rect 42852 32608 42916 32612
rect 47612 32668 47676 32672
rect 47612 32612 47616 32668
rect 47616 32612 47672 32668
rect 47672 32612 47676 32668
rect 47612 32608 47676 32612
rect 47692 32668 47756 32672
rect 47692 32612 47696 32668
rect 47696 32612 47752 32668
rect 47752 32612 47756 32668
rect 47692 32608 47756 32612
rect 47772 32668 47836 32672
rect 47772 32612 47776 32668
rect 47776 32612 47832 32668
rect 47832 32612 47836 32668
rect 47772 32608 47836 32612
rect 47852 32668 47916 32672
rect 47852 32612 47856 32668
rect 47856 32612 47912 32668
rect 47912 32612 47916 32668
rect 47852 32608 47916 32612
rect 52612 32668 52676 32672
rect 52612 32612 52616 32668
rect 52616 32612 52672 32668
rect 52672 32612 52676 32668
rect 52612 32608 52676 32612
rect 52692 32668 52756 32672
rect 52692 32612 52696 32668
rect 52696 32612 52752 32668
rect 52752 32612 52756 32668
rect 52692 32608 52756 32612
rect 52772 32668 52836 32672
rect 52772 32612 52776 32668
rect 52776 32612 52832 32668
rect 52832 32612 52836 32668
rect 52772 32608 52836 32612
rect 52852 32668 52916 32672
rect 52852 32612 52856 32668
rect 52856 32612 52912 32668
rect 52912 32612 52916 32668
rect 52852 32608 52916 32612
rect 57612 32668 57676 32672
rect 57612 32612 57616 32668
rect 57616 32612 57672 32668
rect 57672 32612 57676 32668
rect 57612 32608 57676 32612
rect 57692 32668 57756 32672
rect 57692 32612 57696 32668
rect 57696 32612 57752 32668
rect 57752 32612 57756 32668
rect 57692 32608 57756 32612
rect 57772 32668 57836 32672
rect 57772 32612 57776 32668
rect 57776 32612 57832 32668
rect 57832 32612 57836 32668
rect 57772 32608 57836 32612
rect 57852 32668 57916 32672
rect 57852 32612 57856 32668
rect 57856 32612 57912 32668
rect 57912 32612 57916 32668
rect 57852 32608 57916 32612
rect 1952 32124 2016 32128
rect 1952 32068 1956 32124
rect 1956 32068 2012 32124
rect 2012 32068 2016 32124
rect 1952 32064 2016 32068
rect 2032 32124 2096 32128
rect 2032 32068 2036 32124
rect 2036 32068 2092 32124
rect 2092 32068 2096 32124
rect 2032 32064 2096 32068
rect 2112 32124 2176 32128
rect 2112 32068 2116 32124
rect 2116 32068 2172 32124
rect 2172 32068 2176 32124
rect 2112 32064 2176 32068
rect 2192 32124 2256 32128
rect 2192 32068 2196 32124
rect 2196 32068 2252 32124
rect 2252 32068 2256 32124
rect 2192 32064 2256 32068
rect 6952 32124 7016 32128
rect 6952 32068 6956 32124
rect 6956 32068 7012 32124
rect 7012 32068 7016 32124
rect 6952 32064 7016 32068
rect 7032 32124 7096 32128
rect 7032 32068 7036 32124
rect 7036 32068 7092 32124
rect 7092 32068 7096 32124
rect 7032 32064 7096 32068
rect 7112 32124 7176 32128
rect 7112 32068 7116 32124
rect 7116 32068 7172 32124
rect 7172 32068 7176 32124
rect 7112 32064 7176 32068
rect 7192 32124 7256 32128
rect 7192 32068 7196 32124
rect 7196 32068 7252 32124
rect 7252 32068 7256 32124
rect 7192 32064 7256 32068
rect 11952 32124 12016 32128
rect 11952 32068 11956 32124
rect 11956 32068 12012 32124
rect 12012 32068 12016 32124
rect 11952 32064 12016 32068
rect 12032 32124 12096 32128
rect 12032 32068 12036 32124
rect 12036 32068 12092 32124
rect 12092 32068 12096 32124
rect 12032 32064 12096 32068
rect 12112 32124 12176 32128
rect 12112 32068 12116 32124
rect 12116 32068 12172 32124
rect 12172 32068 12176 32124
rect 12112 32064 12176 32068
rect 12192 32124 12256 32128
rect 12192 32068 12196 32124
rect 12196 32068 12252 32124
rect 12252 32068 12256 32124
rect 12192 32064 12256 32068
rect 16952 32124 17016 32128
rect 16952 32068 16956 32124
rect 16956 32068 17012 32124
rect 17012 32068 17016 32124
rect 16952 32064 17016 32068
rect 17032 32124 17096 32128
rect 17032 32068 17036 32124
rect 17036 32068 17092 32124
rect 17092 32068 17096 32124
rect 17032 32064 17096 32068
rect 17112 32124 17176 32128
rect 17112 32068 17116 32124
rect 17116 32068 17172 32124
rect 17172 32068 17176 32124
rect 17112 32064 17176 32068
rect 17192 32124 17256 32128
rect 17192 32068 17196 32124
rect 17196 32068 17252 32124
rect 17252 32068 17256 32124
rect 17192 32064 17256 32068
rect 21952 32124 22016 32128
rect 21952 32068 21956 32124
rect 21956 32068 22012 32124
rect 22012 32068 22016 32124
rect 21952 32064 22016 32068
rect 22032 32124 22096 32128
rect 22032 32068 22036 32124
rect 22036 32068 22092 32124
rect 22092 32068 22096 32124
rect 22032 32064 22096 32068
rect 22112 32124 22176 32128
rect 22112 32068 22116 32124
rect 22116 32068 22172 32124
rect 22172 32068 22176 32124
rect 22112 32064 22176 32068
rect 22192 32124 22256 32128
rect 22192 32068 22196 32124
rect 22196 32068 22252 32124
rect 22252 32068 22256 32124
rect 22192 32064 22256 32068
rect 26952 32124 27016 32128
rect 26952 32068 26956 32124
rect 26956 32068 27012 32124
rect 27012 32068 27016 32124
rect 26952 32064 27016 32068
rect 27032 32124 27096 32128
rect 27032 32068 27036 32124
rect 27036 32068 27092 32124
rect 27092 32068 27096 32124
rect 27032 32064 27096 32068
rect 27112 32124 27176 32128
rect 27112 32068 27116 32124
rect 27116 32068 27172 32124
rect 27172 32068 27176 32124
rect 27112 32064 27176 32068
rect 27192 32124 27256 32128
rect 27192 32068 27196 32124
rect 27196 32068 27252 32124
rect 27252 32068 27256 32124
rect 27192 32064 27256 32068
rect 31952 32124 32016 32128
rect 31952 32068 31956 32124
rect 31956 32068 32012 32124
rect 32012 32068 32016 32124
rect 31952 32064 32016 32068
rect 32032 32124 32096 32128
rect 32032 32068 32036 32124
rect 32036 32068 32092 32124
rect 32092 32068 32096 32124
rect 32032 32064 32096 32068
rect 32112 32124 32176 32128
rect 32112 32068 32116 32124
rect 32116 32068 32172 32124
rect 32172 32068 32176 32124
rect 32112 32064 32176 32068
rect 32192 32124 32256 32128
rect 32192 32068 32196 32124
rect 32196 32068 32252 32124
rect 32252 32068 32256 32124
rect 32192 32064 32256 32068
rect 36952 32124 37016 32128
rect 36952 32068 36956 32124
rect 36956 32068 37012 32124
rect 37012 32068 37016 32124
rect 36952 32064 37016 32068
rect 37032 32124 37096 32128
rect 37032 32068 37036 32124
rect 37036 32068 37092 32124
rect 37092 32068 37096 32124
rect 37032 32064 37096 32068
rect 37112 32124 37176 32128
rect 37112 32068 37116 32124
rect 37116 32068 37172 32124
rect 37172 32068 37176 32124
rect 37112 32064 37176 32068
rect 37192 32124 37256 32128
rect 37192 32068 37196 32124
rect 37196 32068 37252 32124
rect 37252 32068 37256 32124
rect 37192 32064 37256 32068
rect 41952 32124 42016 32128
rect 41952 32068 41956 32124
rect 41956 32068 42012 32124
rect 42012 32068 42016 32124
rect 41952 32064 42016 32068
rect 42032 32124 42096 32128
rect 42032 32068 42036 32124
rect 42036 32068 42092 32124
rect 42092 32068 42096 32124
rect 42032 32064 42096 32068
rect 42112 32124 42176 32128
rect 42112 32068 42116 32124
rect 42116 32068 42172 32124
rect 42172 32068 42176 32124
rect 42112 32064 42176 32068
rect 42192 32124 42256 32128
rect 42192 32068 42196 32124
rect 42196 32068 42252 32124
rect 42252 32068 42256 32124
rect 42192 32064 42256 32068
rect 46952 32124 47016 32128
rect 46952 32068 46956 32124
rect 46956 32068 47012 32124
rect 47012 32068 47016 32124
rect 46952 32064 47016 32068
rect 47032 32124 47096 32128
rect 47032 32068 47036 32124
rect 47036 32068 47092 32124
rect 47092 32068 47096 32124
rect 47032 32064 47096 32068
rect 47112 32124 47176 32128
rect 47112 32068 47116 32124
rect 47116 32068 47172 32124
rect 47172 32068 47176 32124
rect 47112 32064 47176 32068
rect 47192 32124 47256 32128
rect 47192 32068 47196 32124
rect 47196 32068 47252 32124
rect 47252 32068 47256 32124
rect 47192 32064 47256 32068
rect 51952 32124 52016 32128
rect 51952 32068 51956 32124
rect 51956 32068 52012 32124
rect 52012 32068 52016 32124
rect 51952 32064 52016 32068
rect 52032 32124 52096 32128
rect 52032 32068 52036 32124
rect 52036 32068 52092 32124
rect 52092 32068 52096 32124
rect 52032 32064 52096 32068
rect 52112 32124 52176 32128
rect 52112 32068 52116 32124
rect 52116 32068 52172 32124
rect 52172 32068 52176 32124
rect 52112 32064 52176 32068
rect 52192 32124 52256 32128
rect 52192 32068 52196 32124
rect 52196 32068 52252 32124
rect 52252 32068 52256 32124
rect 52192 32064 52256 32068
rect 56952 32124 57016 32128
rect 56952 32068 56956 32124
rect 56956 32068 57012 32124
rect 57012 32068 57016 32124
rect 56952 32064 57016 32068
rect 57032 32124 57096 32128
rect 57032 32068 57036 32124
rect 57036 32068 57092 32124
rect 57092 32068 57096 32124
rect 57032 32064 57096 32068
rect 57112 32124 57176 32128
rect 57112 32068 57116 32124
rect 57116 32068 57172 32124
rect 57172 32068 57176 32124
rect 57112 32064 57176 32068
rect 57192 32124 57256 32128
rect 57192 32068 57196 32124
rect 57196 32068 57252 32124
rect 57252 32068 57256 32124
rect 57192 32064 57256 32068
rect 2612 31580 2676 31584
rect 2612 31524 2616 31580
rect 2616 31524 2672 31580
rect 2672 31524 2676 31580
rect 2612 31520 2676 31524
rect 2692 31580 2756 31584
rect 2692 31524 2696 31580
rect 2696 31524 2752 31580
rect 2752 31524 2756 31580
rect 2692 31520 2756 31524
rect 2772 31580 2836 31584
rect 2772 31524 2776 31580
rect 2776 31524 2832 31580
rect 2832 31524 2836 31580
rect 2772 31520 2836 31524
rect 2852 31580 2916 31584
rect 2852 31524 2856 31580
rect 2856 31524 2912 31580
rect 2912 31524 2916 31580
rect 2852 31520 2916 31524
rect 7612 31580 7676 31584
rect 7612 31524 7616 31580
rect 7616 31524 7672 31580
rect 7672 31524 7676 31580
rect 7612 31520 7676 31524
rect 7692 31580 7756 31584
rect 7692 31524 7696 31580
rect 7696 31524 7752 31580
rect 7752 31524 7756 31580
rect 7692 31520 7756 31524
rect 7772 31580 7836 31584
rect 7772 31524 7776 31580
rect 7776 31524 7832 31580
rect 7832 31524 7836 31580
rect 7772 31520 7836 31524
rect 7852 31580 7916 31584
rect 7852 31524 7856 31580
rect 7856 31524 7912 31580
rect 7912 31524 7916 31580
rect 7852 31520 7916 31524
rect 12612 31580 12676 31584
rect 12612 31524 12616 31580
rect 12616 31524 12672 31580
rect 12672 31524 12676 31580
rect 12612 31520 12676 31524
rect 12692 31580 12756 31584
rect 12692 31524 12696 31580
rect 12696 31524 12752 31580
rect 12752 31524 12756 31580
rect 12692 31520 12756 31524
rect 12772 31580 12836 31584
rect 12772 31524 12776 31580
rect 12776 31524 12832 31580
rect 12832 31524 12836 31580
rect 12772 31520 12836 31524
rect 12852 31580 12916 31584
rect 12852 31524 12856 31580
rect 12856 31524 12912 31580
rect 12912 31524 12916 31580
rect 12852 31520 12916 31524
rect 17612 31580 17676 31584
rect 17612 31524 17616 31580
rect 17616 31524 17672 31580
rect 17672 31524 17676 31580
rect 17612 31520 17676 31524
rect 17692 31580 17756 31584
rect 17692 31524 17696 31580
rect 17696 31524 17752 31580
rect 17752 31524 17756 31580
rect 17692 31520 17756 31524
rect 17772 31580 17836 31584
rect 17772 31524 17776 31580
rect 17776 31524 17832 31580
rect 17832 31524 17836 31580
rect 17772 31520 17836 31524
rect 17852 31580 17916 31584
rect 17852 31524 17856 31580
rect 17856 31524 17912 31580
rect 17912 31524 17916 31580
rect 17852 31520 17916 31524
rect 22612 31580 22676 31584
rect 22612 31524 22616 31580
rect 22616 31524 22672 31580
rect 22672 31524 22676 31580
rect 22612 31520 22676 31524
rect 22692 31580 22756 31584
rect 22692 31524 22696 31580
rect 22696 31524 22752 31580
rect 22752 31524 22756 31580
rect 22692 31520 22756 31524
rect 22772 31580 22836 31584
rect 22772 31524 22776 31580
rect 22776 31524 22832 31580
rect 22832 31524 22836 31580
rect 22772 31520 22836 31524
rect 22852 31580 22916 31584
rect 22852 31524 22856 31580
rect 22856 31524 22912 31580
rect 22912 31524 22916 31580
rect 22852 31520 22916 31524
rect 27612 31580 27676 31584
rect 27612 31524 27616 31580
rect 27616 31524 27672 31580
rect 27672 31524 27676 31580
rect 27612 31520 27676 31524
rect 27692 31580 27756 31584
rect 27692 31524 27696 31580
rect 27696 31524 27752 31580
rect 27752 31524 27756 31580
rect 27692 31520 27756 31524
rect 27772 31580 27836 31584
rect 27772 31524 27776 31580
rect 27776 31524 27832 31580
rect 27832 31524 27836 31580
rect 27772 31520 27836 31524
rect 27852 31580 27916 31584
rect 27852 31524 27856 31580
rect 27856 31524 27912 31580
rect 27912 31524 27916 31580
rect 27852 31520 27916 31524
rect 32612 31580 32676 31584
rect 32612 31524 32616 31580
rect 32616 31524 32672 31580
rect 32672 31524 32676 31580
rect 32612 31520 32676 31524
rect 32692 31580 32756 31584
rect 32692 31524 32696 31580
rect 32696 31524 32752 31580
rect 32752 31524 32756 31580
rect 32692 31520 32756 31524
rect 32772 31580 32836 31584
rect 32772 31524 32776 31580
rect 32776 31524 32832 31580
rect 32832 31524 32836 31580
rect 32772 31520 32836 31524
rect 32852 31580 32916 31584
rect 32852 31524 32856 31580
rect 32856 31524 32912 31580
rect 32912 31524 32916 31580
rect 32852 31520 32916 31524
rect 37612 31580 37676 31584
rect 37612 31524 37616 31580
rect 37616 31524 37672 31580
rect 37672 31524 37676 31580
rect 37612 31520 37676 31524
rect 37692 31580 37756 31584
rect 37692 31524 37696 31580
rect 37696 31524 37752 31580
rect 37752 31524 37756 31580
rect 37692 31520 37756 31524
rect 37772 31580 37836 31584
rect 37772 31524 37776 31580
rect 37776 31524 37832 31580
rect 37832 31524 37836 31580
rect 37772 31520 37836 31524
rect 37852 31580 37916 31584
rect 37852 31524 37856 31580
rect 37856 31524 37912 31580
rect 37912 31524 37916 31580
rect 37852 31520 37916 31524
rect 42612 31580 42676 31584
rect 42612 31524 42616 31580
rect 42616 31524 42672 31580
rect 42672 31524 42676 31580
rect 42612 31520 42676 31524
rect 42692 31580 42756 31584
rect 42692 31524 42696 31580
rect 42696 31524 42752 31580
rect 42752 31524 42756 31580
rect 42692 31520 42756 31524
rect 42772 31580 42836 31584
rect 42772 31524 42776 31580
rect 42776 31524 42832 31580
rect 42832 31524 42836 31580
rect 42772 31520 42836 31524
rect 42852 31580 42916 31584
rect 42852 31524 42856 31580
rect 42856 31524 42912 31580
rect 42912 31524 42916 31580
rect 42852 31520 42916 31524
rect 47612 31580 47676 31584
rect 47612 31524 47616 31580
rect 47616 31524 47672 31580
rect 47672 31524 47676 31580
rect 47612 31520 47676 31524
rect 47692 31580 47756 31584
rect 47692 31524 47696 31580
rect 47696 31524 47752 31580
rect 47752 31524 47756 31580
rect 47692 31520 47756 31524
rect 47772 31580 47836 31584
rect 47772 31524 47776 31580
rect 47776 31524 47832 31580
rect 47832 31524 47836 31580
rect 47772 31520 47836 31524
rect 47852 31580 47916 31584
rect 47852 31524 47856 31580
rect 47856 31524 47912 31580
rect 47912 31524 47916 31580
rect 47852 31520 47916 31524
rect 52612 31580 52676 31584
rect 52612 31524 52616 31580
rect 52616 31524 52672 31580
rect 52672 31524 52676 31580
rect 52612 31520 52676 31524
rect 52692 31580 52756 31584
rect 52692 31524 52696 31580
rect 52696 31524 52752 31580
rect 52752 31524 52756 31580
rect 52692 31520 52756 31524
rect 52772 31580 52836 31584
rect 52772 31524 52776 31580
rect 52776 31524 52832 31580
rect 52832 31524 52836 31580
rect 52772 31520 52836 31524
rect 52852 31580 52916 31584
rect 52852 31524 52856 31580
rect 52856 31524 52912 31580
rect 52912 31524 52916 31580
rect 52852 31520 52916 31524
rect 57612 31580 57676 31584
rect 57612 31524 57616 31580
rect 57616 31524 57672 31580
rect 57672 31524 57676 31580
rect 57612 31520 57676 31524
rect 57692 31580 57756 31584
rect 57692 31524 57696 31580
rect 57696 31524 57752 31580
rect 57752 31524 57756 31580
rect 57692 31520 57756 31524
rect 57772 31580 57836 31584
rect 57772 31524 57776 31580
rect 57776 31524 57832 31580
rect 57832 31524 57836 31580
rect 57772 31520 57836 31524
rect 57852 31580 57916 31584
rect 57852 31524 57856 31580
rect 57856 31524 57912 31580
rect 57912 31524 57916 31580
rect 57852 31520 57916 31524
rect 1952 31036 2016 31040
rect 1952 30980 1956 31036
rect 1956 30980 2012 31036
rect 2012 30980 2016 31036
rect 1952 30976 2016 30980
rect 2032 31036 2096 31040
rect 2032 30980 2036 31036
rect 2036 30980 2092 31036
rect 2092 30980 2096 31036
rect 2032 30976 2096 30980
rect 2112 31036 2176 31040
rect 2112 30980 2116 31036
rect 2116 30980 2172 31036
rect 2172 30980 2176 31036
rect 2112 30976 2176 30980
rect 2192 31036 2256 31040
rect 2192 30980 2196 31036
rect 2196 30980 2252 31036
rect 2252 30980 2256 31036
rect 2192 30976 2256 30980
rect 6952 31036 7016 31040
rect 6952 30980 6956 31036
rect 6956 30980 7012 31036
rect 7012 30980 7016 31036
rect 6952 30976 7016 30980
rect 7032 31036 7096 31040
rect 7032 30980 7036 31036
rect 7036 30980 7092 31036
rect 7092 30980 7096 31036
rect 7032 30976 7096 30980
rect 7112 31036 7176 31040
rect 7112 30980 7116 31036
rect 7116 30980 7172 31036
rect 7172 30980 7176 31036
rect 7112 30976 7176 30980
rect 7192 31036 7256 31040
rect 7192 30980 7196 31036
rect 7196 30980 7252 31036
rect 7252 30980 7256 31036
rect 7192 30976 7256 30980
rect 11952 31036 12016 31040
rect 11952 30980 11956 31036
rect 11956 30980 12012 31036
rect 12012 30980 12016 31036
rect 11952 30976 12016 30980
rect 12032 31036 12096 31040
rect 12032 30980 12036 31036
rect 12036 30980 12092 31036
rect 12092 30980 12096 31036
rect 12032 30976 12096 30980
rect 12112 31036 12176 31040
rect 12112 30980 12116 31036
rect 12116 30980 12172 31036
rect 12172 30980 12176 31036
rect 12112 30976 12176 30980
rect 12192 31036 12256 31040
rect 12192 30980 12196 31036
rect 12196 30980 12252 31036
rect 12252 30980 12256 31036
rect 12192 30976 12256 30980
rect 16952 31036 17016 31040
rect 16952 30980 16956 31036
rect 16956 30980 17012 31036
rect 17012 30980 17016 31036
rect 16952 30976 17016 30980
rect 17032 31036 17096 31040
rect 17032 30980 17036 31036
rect 17036 30980 17092 31036
rect 17092 30980 17096 31036
rect 17032 30976 17096 30980
rect 17112 31036 17176 31040
rect 17112 30980 17116 31036
rect 17116 30980 17172 31036
rect 17172 30980 17176 31036
rect 17112 30976 17176 30980
rect 17192 31036 17256 31040
rect 17192 30980 17196 31036
rect 17196 30980 17252 31036
rect 17252 30980 17256 31036
rect 17192 30976 17256 30980
rect 21952 31036 22016 31040
rect 21952 30980 21956 31036
rect 21956 30980 22012 31036
rect 22012 30980 22016 31036
rect 21952 30976 22016 30980
rect 22032 31036 22096 31040
rect 22032 30980 22036 31036
rect 22036 30980 22092 31036
rect 22092 30980 22096 31036
rect 22032 30976 22096 30980
rect 22112 31036 22176 31040
rect 22112 30980 22116 31036
rect 22116 30980 22172 31036
rect 22172 30980 22176 31036
rect 22112 30976 22176 30980
rect 22192 31036 22256 31040
rect 22192 30980 22196 31036
rect 22196 30980 22252 31036
rect 22252 30980 22256 31036
rect 22192 30976 22256 30980
rect 26952 31036 27016 31040
rect 26952 30980 26956 31036
rect 26956 30980 27012 31036
rect 27012 30980 27016 31036
rect 26952 30976 27016 30980
rect 27032 31036 27096 31040
rect 27032 30980 27036 31036
rect 27036 30980 27092 31036
rect 27092 30980 27096 31036
rect 27032 30976 27096 30980
rect 27112 31036 27176 31040
rect 27112 30980 27116 31036
rect 27116 30980 27172 31036
rect 27172 30980 27176 31036
rect 27112 30976 27176 30980
rect 27192 31036 27256 31040
rect 27192 30980 27196 31036
rect 27196 30980 27252 31036
rect 27252 30980 27256 31036
rect 27192 30976 27256 30980
rect 31952 31036 32016 31040
rect 31952 30980 31956 31036
rect 31956 30980 32012 31036
rect 32012 30980 32016 31036
rect 31952 30976 32016 30980
rect 32032 31036 32096 31040
rect 32032 30980 32036 31036
rect 32036 30980 32092 31036
rect 32092 30980 32096 31036
rect 32032 30976 32096 30980
rect 32112 31036 32176 31040
rect 32112 30980 32116 31036
rect 32116 30980 32172 31036
rect 32172 30980 32176 31036
rect 32112 30976 32176 30980
rect 32192 31036 32256 31040
rect 32192 30980 32196 31036
rect 32196 30980 32252 31036
rect 32252 30980 32256 31036
rect 32192 30976 32256 30980
rect 36952 31036 37016 31040
rect 36952 30980 36956 31036
rect 36956 30980 37012 31036
rect 37012 30980 37016 31036
rect 36952 30976 37016 30980
rect 37032 31036 37096 31040
rect 37032 30980 37036 31036
rect 37036 30980 37092 31036
rect 37092 30980 37096 31036
rect 37032 30976 37096 30980
rect 37112 31036 37176 31040
rect 37112 30980 37116 31036
rect 37116 30980 37172 31036
rect 37172 30980 37176 31036
rect 37112 30976 37176 30980
rect 37192 31036 37256 31040
rect 37192 30980 37196 31036
rect 37196 30980 37252 31036
rect 37252 30980 37256 31036
rect 37192 30976 37256 30980
rect 41952 31036 42016 31040
rect 41952 30980 41956 31036
rect 41956 30980 42012 31036
rect 42012 30980 42016 31036
rect 41952 30976 42016 30980
rect 42032 31036 42096 31040
rect 42032 30980 42036 31036
rect 42036 30980 42092 31036
rect 42092 30980 42096 31036
rect 42032 30976 42096 30980
rect 42112 31036 42176 31040
rect 42112 30980 42116 31036
rect 42116 30980 42172 31036
rect 42172 30980 42176 31036
rect 42112 30976 42176 30980
rect 42192 31036 42256 31040
rect 42192 30980 42196 31036
rect 42196 30980 42252 31036
rect 42252 30980 42256 31036
rect 42192 30976 42256 30980
rect 46952 31036 47016 31040
rect 46952 30980 46956 31036
rect 46956 30980 47012 31036
rect 47012 30980 47016 31036
rect 46952 30976 47016 30980
rect 47032 31036 47096 31040
rect 47032 30980 47036 31036
rect 47036 30980 47092 31036
rect 47092 30980 47096 31036
rect 47032 30976 47096 30980
rect 47112 31036 47176 31040
rect 47112 30980 47116 31036
rect 47116 30980 47172 31036
rect 47172 30980 47176 31036
rect 47112 30976 47176 30980
rect 47192 31036 47256 31040
rect 47192 30980 47196 31036
rect 47196 30980 47252 31036
rect 47252 30980 47256 31036
rect 47192 30976 47256 30980
rect 51952 31036 52016 31040
rect 51952 30980 51956 31036
rect 51956 30980 52012 31036
rect 52012 30980 52016 31036
rect 51952 30976 52016 30980
rect 52032 31036 52096 31040
rect 52032 30980 52036 31036
rect 52036 30980 52092 31036
rect 52092 30980 52096 31036
rect 52032 30976 52096 30980
rect 52112 31036 52176 31040
rect 52112 30980 52116 31036
rect 52116 30980 52172 31036
rect 52172 30980 52176 31036
rect 52112 30976 52176 30980
rect 52192 31036 52256 31040
rect 52192 30980 52196 31036
rect 52196 30980 52252 31036
rect 52252 30980 52256 31036
rect 52192 30976 52256 30980
rect 56952 31036 57016 31040
rect 56952 30980 56956 31036
rect 56956 30980 57012 31036
rect 57012 30980 57016 31036
rect 56952 30976 57016 30980
rect 57032 31036 57096 31040
rect 57032 30980 57036 31036
rect 57036 30980 57092 31036
rect 57092 30980 57096 31036
rect 57032 30976 57096 30980
rect 57112 31036 57176 31040
rect 57112 30980 57116 31036
rect 57116 30980 57172 31036
rect 57172 30980 57176 31036
rect 57112 30976 57176 30980
rect 57192 31036 57256 31040
rect 57192 30980 57196 31036
rect 57196 30980 57252 31036
rect 57252 30980 57256 31036
rect 57192 30976 57256 30980
rect 2612 30492 2676 30496
rect 2612 30436 2616 30492
rect 2616 30436 2672 30492
rect 2672 30436 2676 30492
rect 2612 30432 2676 30436
rect 2692 30492 2756 30496
rect 2692 30436 2696 30492
rect 2696 30436 2752 30492
rect 2752 30436 2756 30492
rect 2692 30432 2756 30436
rect 2772 30492 2836 30496
rect 2772 30436 2776 30492
rect 2776 30436 2832 30492
rect 2832 30436 2836 30492
rect 2772 30432 2836 30436
rect 2852 30492 2916 30496
rect 2852 30436 2856 30492
rect 2856 30436 2912 30492
rect 2912 30436 2916 30492
rect 2852 30432 2916 30436
rect 7612 30492 7676 30496
rect 7612 30436 7616 30492
rect 7616 30436 7672 30492
rect 7672 30436 7676 30492
rect 7612 30432 7676 30436
rect 7692 30492 7756 30496
rect 7692 30436 7696 30492
rect 7696 30436 7752 30492
rect 7752 30436 7756 30492
rect 7692 30432 7756 30436
rect 7772 30492 7836 30496
rect 7772 30436 7776 30492
rect 7776 30436 7832 30492
rect 7832 30436 7836 30492
rect 7772 30432 7836 30436
rect 7852 30492 7916 30496
rect 7852 30436 7856 30492
rect 7856 30436 7912 30492
rect 7912 30436 7916 30492
rect 7852 30432 7916 30436
rect 12612 30492 12676 30496
rect 12612 30436 12616 30492
rect 12616 30436 12672 30492
rect 12672 30436 12676 30492
rect 12612 30432 12676 30436
rect 12692 30492 12756 30496
rect 12692 30436 12696 30492
rect 12696 30436 12752 30492
rect 12752 30436 12756 30492
rect 12692 30432 12756 30436
rect 12772 30492 12836 30496
rect 12772 30436 12776 30492
rect 12776 30436 12832 30492
rect 12832 30436 12836 30492
rect 12772 30432 12836 30436
rect 12852 30492 12916 30496
rect 12852 30436 12856 30492
rect 12856 30436 12912 30492
rect 12912 30436 12916 30492
rect 12852 30432 12916 30436
rect 17612 30492 17676 30496
rect 17612 30436 17616 30492
rect 17616 30436 17672 30492
rect 17672 30436 17676 30492
rect 17612 30432 17676 30436
rect 17692 30492 17756 30496
rect 17692 30436 17696 30492
rect 17696 30436 17752 30492
rect 17752 30436 17756 30492
rect 17692 30432 17756 30436
rect 17772 30492 17836 30496
rect 17772 30436 17776 30492
rect 17776 30436 17832 30492
rect 17832 30436 17836 30492
rect 17772 30432 17836 30436
rect 17852 30492 17916 30496
rect 17852 30436 17856 30492
rect 17856 30436 17912 30492
rect 17912 30436 17916 30492
rect 17852 30432 17916 30436
rect 22612 30492 22676 30496
rect 22612 30436 22616 30492
rect 22616 30436 22672 30492
rect 22672 30436 22676 30492
rect 22612 30432 22676 30436
rect 22692 30492 22756 30496
rect 22692 30436 22696 30492
rect 22696 30436 22752 30492
rect 22752 30436 22756 30492
rect 22692 30432 22756 30436
rect 22772 30492 22836 30496
rect 22772 30436 22776 30492
rect 22776 30436 22832 30492
rect 22832 30436 22836 30492
rect 22772 30432 22836 30436
rect 22852 30492 22916 30496
rect 22852 30436 22856 30492
rect 22856 30436 22912 30492
rect 22912 30436 22916 30492
rect 22852 30432 22916 30436
rect 27612 30492 27676 30496
rect 27612 30436 27616 30492
rect 27616 30436 27672 30492
rect 27672 30436 27676 30492
rect 27612 30432 27676 30436
rect 27692 30492 27756 30496
rect 27692 30436 27696 30492
rect 27696 30436 27752 30492
rect 27752 30436 27756 30492
rect 27692 30432 27756 30436
rect 27772 30492 27836 30496
rect 27772 30436 27776 30492
rect 27776 30436 27832 30492
rect 27832 30436 27836 30492
rect 27772 30432 27836 30436
rect 27852 30492 27916 30496
rect 27852 30436 27856 30492
rect 27856 30436 27912 30492
rect 27912 30436 27916 30492
rect 27852 30432 27916 30436
rect 32612 30492 32676 30496
rect 32612 30436 32616 30492
rect 32616 30436 32672 30492
rect 32672 30436 32676 30492
rect 32612 30432 32676 30436
rect 32692 30492 32756 30496
rect 32692 30436 32696 30492
rect 32696 30436 32752 30492
rect 32752 30436 32756 30492
rect 32692 30432 32756 30436
rect 32772 30492 32836 30496
rect 32772 30436 32776 30492
rect 32776 30436 32832 30492
rect 32832 30436 32836 30492
rect 32772 30432 32836 30436
rect 32852 30492 32916 30496
rect 32852 30436 32856 30492
rect 32856 30436 32912 30492
rect 32912 30436 32916 30492
rect 32852 30432 32916 30436
rect 37612 30492 37676 30496
rect 37612 30436 37616 30492
rect 37616 30436 37672 30492
rect 37672 30436 37676 30492
rect 37612 30432 37676 30436
rect 37692 30492 37756 30496
rect 37692 30436 37696 30492
rect 37696 30436 37752 30492
rect 37752 30436 37756 30492
rect 37692 30432 37756 30436
rect 37772 30492 37836 30496
rect 37772 30436 37776 30492
rect 37776 30436 37832 30492
rect 37832 30436 37836 30492
rect 37772 30432 37836 30436
rect 37852 30492 37916 30496
rect 37852 30436 37856 30492
rect 37856 30436 37912 30492
rect 37912 30436 37916 30492
rect 37852 30432 37916 30436
rect 42612 30492 42676 30496
rect 42612 30436 42616 30492
rect 42616 30436 42672 30492
rect 42672 30436 42676 30492
rect 42612 30432 42676 30436
rect 42692 30492 42756 30496
rect 42692 30436 42696 30492
rect 42696 30436 42752 30492
rect 42752 30436 42756 30492
rect 42692 30432 42756 30436
rect 42772 30492 42836 30496
rect 42772 30436 42776 30492
rect 42776 30436 42832 30492
rect 42832 30436 42836 30492
rect 42772 30432 42836 30436
rect 42852 30492 42916 30496
rect 42852 30436 42856 30492
rect 42856 30436 42912 30492
rect 42912 30436 42916 30492
rect 42852 30432 42916 30436
rect 47612 30492 47676 30496
rect 47612 30436 47616 30492
rect 47616 30436 47672 30492
rect 47672 30436 47676 30492
rect 47612 30432 47676 30436
rect 47692 30492 47756 30496
rect 47692 30436 47696 30492
rect 47696 30436 47752 30492
rect 47752 30436 47756 30492
rect 47692 30432 47756 30436
rect 47772 30492 47836 30496
rect 47772 30436 47776 30492
rect 47776 30436 47832 30492
rect 47832 30436 47836 30492
rect 47772 30432 47836 30436
rect 47852 30492 47916 30496
rect 47852 30436 47856 30492
rect 47856 30436 47912 30492
rect 47912 30436 47916 30492
rect 47852 30432 47916 30436
rect 52612 30492 52676 30496
rect 52612 30436 52616 30492
rect 52616 30436 52672 30492
rect 52672 30436 52676 30492
rect 52612 30432 52676 30436
rect 52692 30492 52756 30496
rect 52692 30436 52696 30492
rect 52696 30436 52752 30492
rect 52752 30436 52756 30492
rect 52692 30432 52756 30436
rect 52772 30492 52836 30496
rect 52772 30436 52776 30492
rect 52776 30436 52832 30492
rect 52832 30436 52836 30492
rect 52772 30432 52836 30436
rect 52852 30492 52916 30496
rect 52852 30436 52856 30492
rect 52856 30436 52912 30492
rect 52912 30436 52916 30492
rect 52852 30432 52916 30436
rect 57612 30492 57676 30496
rect 57612 30436 57616 30492
rect 57616 30436 57672 30492
rect 57672 30436 57676 30492
rect 57612 30432 57676 30436
rect 57692 30492 57756 30496
rect 57692 30436 57696 30492
rect 57696 30436 57752 30492
rect 57752 30436 57756 30492
rect 57692 30432 57756 30436
rect 57772 30492 57836 30496
rect 57772 30436 57776 30492
rect 57776 30436 57832 30492
rect 57832 30436 57836 30492
rect 57772 30432 57836 30436
rect 57852 30492 57916 30496
rect 57852 30436 57856 30492
rect 57856 30436 57912 30492
rect 57912 30436 57916 30492
rect 57852 30432 57916 30436
rect 1952 29948 2016 29952
rect 1952 29892 1956 29948
rect 1956 29892 2012 29948
rect 2012 29892 2016 29948
rect 1952 29888 2016 29892
rect 2032 29948 2096 29952
rect 2032 29892 2036 29948
rect 2036 29892 2092 29948
rect 2092 29892 2096 29948
rect 2032 29888 2096 29892
rect 2112 29948 2176 29952
rect 2112 29892 2116 29948
rect 2116 29892 2172 29948
rect 2172 29892 2176 29948
rect 2112 29888 2176 29892
rect 2192 29948 2256 29952
rect 2192 29892 2196 29948
rect 2196 29892 2252 29948
rect 2252 29892 2256 29948
rect 2192 29888 2256 29892
rect 6952 29948 7016 29952
rect 6952 29892 6956 29948
rect 6956 29892 7012 29948
rect 7012 29892 7016 29948
rect 6952 29888 7016 29892
rect 7032 29948 7096 29952
rect 7032 29892 7036 29948
rect 7036 29892 7092 29948
rect 7092 29892 7096 29948
rect 7032 29888 7096 29892
rect 7112 29948 7176 29952
rect 7112 29892 7116 29948
rect 7116 29892 7172 29948
rect 7172 29892 7176 29948
rect 7112 29888 7176 29892
rect 7192 29948 7256 29952
rect 7192 29892 7196 29948
rect 7196 29892 7252 29948
rect 7252 29892 7256 29948
rect 7192 29888 7256 29892
rect 11952 29948 12016 29952
rect 11952 29892 11956 29948
rect 11956 29892 12012 29948
rect 12012 29892 12016 29948
rect 11952 29888 12016 29892
rect 12032 29948 12096 29952
rect 12032 29892 12036 29948
rect 12036 29892 12092 29948
rect 12092 29892 12096 29948
rect 12032 29888 12096 29892
rect 12112 29948 12176 29952
rect 12112 29892 12116 29948
rect 12116 29892 12172 29948
rect 12172 29892 12176 29948
rect 12112 29888 12176 29892
rect 12192 29948 12256 29952
rect 12192 29892 12196 29948
rect 12196 29892 12252 29948
rect 12252 29892 12256 29948
rect 12192 29888 12256 29892
rect 16952 29948 17016 29952
rect 16952 29892 16956 29948
rect 16956 29892 17012 29948
rect 17012 29892 17016 29948
rect 16952 29888 17016 29892
rect 17032 29948 17096 29952
rect 17032 29892 17036 29948
rect 17036 29892 17092 29948
rect 17092 29892 17096 29948
rect 17032 29888 17096 29892
rect 17112 29948 17176 29952
rect 17112 29892 17116 29948
rect 17116 29892 17172 29948
rect 17172 29892 17176 29948
rect 17112 29888 17176 29892
rect 17192 29948 17256 29952
rect 17192 29892 17196 29948
rect 17196 29892 17252 29948
rect 17252 29892 17256 29948
rect 17192 29888 17256 29892
rect 21952 29948 22016 29952
rect 21952 29892 21956 29948
rect 21956 29892 22012 29948
rect 22012 29892 22016 29948
rect 21952 29888 22016 29892
rect 22032 29948 22096 29952
rect 22032 29892 22036 29948
rect 22036 29892 22092 29948
rect 22092 29892 22096 29948
rect 22032 29888 22096 29892
rect 22112 29948 22176 29952
rect 22112 29892 22116 29948
rect 22116 29892 22172 29948
rect 22172 29892 22176 29948
rect 22112 29888 22176 29892
rect 22192 29948 22256 29952
rect 22192 29892 22196 29948
rect 22196 29892 22252 29948
rect 22252 29892 22256 29948
rect 22192 29888 22256 29892
rect 26952 29948 27016 29952
rect 26952 29892 26956 29948
rect 26956 29892 27012 29948
rect 27012 29892 27016 29948
rect 26952 29888 27016 29892
rect 27032 29948 27096 29952
rect 27032 29892 27036 29948
rect 27036 29892 27092 29948
rect 27092 29892 27096 29948
rect 27032 29888 27096 29892
rect 27112 29948 27176 29952
rect 27112 29892 27116 29948
rect 27116 29892 27172 29948
rect 27172 29892 27176 29948
rect 27112 29888 27176 29892
rect 27192 29948 27256 29952
rect 27192 29892 27196 29948
rect 27196 29892 27252 29948
rect 27252 29892 27256 29948
rect 27192 29888 27256 29892
rect 31952 29948 32016 29952
rect 31952 29892 31956 29948
rect 31956 29892 32012 29948
rect 32012 29892 32016 29948
rect 31952 29888 32016 29892
rect 32032 29948 32096 29952
rect 32032 29892 32036 29948
rect 32036 29892 32092 29948
rect 32092 29892 32096 29948
rect 32032 29888 32096 29892
rect 32112 29948 32176 29952
rect 32112 29892 32116 29948
rect 32116 29892 32172 29948
rect 32172 29892 32176 29948
rect 32112 29888 32176 29892
rect 32192 29948 32256 29952
rect 32192 29892 32196 29948
rect 32196 29892 32252 29948
rect 32252 29892 32256 29948
rect 32192 29888 32256 29892
rect 36952 29948 37016 29952
rect 36952 29892 36956 29948
rect 36956 29892 37012 29948
rect 37012 29892 37016 29948
rect 36952 29888 37016 29892
rect 37032 29948 37096 29952
rect 37032 29892 37036 29948
rect 37036 29892 37092 29948
rect 37092 29892 37096 29948
rect 37032 29888 37096 29892
rect 37112 29948 37176 29952
rect 37112 29892 37116 29948
rect 37116 29892 37172 29948
rect 37172 29892 37176 29948
rect 37112 29888 37176 29892
rect 37192 29948 37256 29952
rect 37192 29892 37196 29948
rect 37196 29892 37252 29948
rect 37252 29892 37256 29948
rect 37192 29888 37256 29892
rect 41952 29948 42016 29952
rect 41952 29892 41956 29948
rect 41956 29892 42012 29948
rect 42012 29892 42016 29948
rect 41952 29888 42016 29892
rect 42032 29948 42096 29952
rect 42032 29892 42036 29948
rect 42036 29892 42092 29948
rect 42092 29892 42096 29948
rect 42032 29888 42096 29892
rect 42112 29948 42176 29952
rect 42112 29892 42116 29948
rect 42116 29892 42172 29948
rect 42172 29892 42176 29948
rect 42112 29888 42176 29892
rect 42192 29948 42256 29952
rect 42192 29892 42196 29948
rect 42196 29892 42252 29948
rect 42252 29892 42256 29948
rect 42192 29888 42256 29892
rect 46952 29948 47016 29952
rect 46952 29892 46956 29948
rect 46956 29892 47012 29948
rect 47012 29892 47016 29948
rect 46952 29888 47016 29892
rect 47032 29948 47096 29952
rect 47032 29892 47036 29948
rect 47036 29892 47092 29948
rect 47092 29892 47096 29948
rect 47032 29888 47096 29892
rect 47112 29948 47176 29952
rect 47112 29892 47116 29948
rect 47116 29892 47172 29948
rect 47172 29892 47176 29948
rect 47112 29888 47176 29892
rect 47192 29948 47256 29952
rect 47192 29892 47196 29948
rect 47196 29892 47252 29948
rect 47252 29892 47256 29948
rect 47192 29888 47256 29892
rect 51952 29948 52016 29952
rect 51952 29892 51956 29948
rect 51956 29892 52012 29948
rect 52012 29892 52016 29948
rect 51952 29888 52016 29892
rect 52032 29948 52096 29952
rect 52032 29892 52036 29948
rect 52036 29892 52092 29948
rect 52092 29892 52096 29948
rect 52032 29888 52096 29892
rect 52112 29948 52176 29952
rect 52112 29892 52116 29948
rect 52116 29892 52172 29948
rect 52172 29892 52176 29948
rect 52112 29888 52176 29892
rect 52192 29948 52256 29952
rect 52192 29892 52196 29948
rect 52196 29892 52252 29948
rect 52252 29892 52256 29948
rect 52192 29888 52256 29892
rect 56952 29948 57016 29952
rect 56952 29892 56956 29948
rect 56956 29892 57012 29948
rect 57012 29892 57016 29948
rect 56952 29888 57016 29892
rect 57032 29948 57096 29952
rect 57032 29892 57036 29948
rect 57036 29892 57092 29948
rect 57092 29892 57096 29948
rect 57032 29888 57096 29892
rect 57112 29948 57176 29952
rect 57112 29892 57116 29948
rect 57116 29892 57172 29948
rect 57172 29892 57176 29948
rect 57112 29888 57176 29892
rect 57192 29948 57256 29952
rect 57192 29892 57196 29948
rect 57196 29892 57252 29948
rect 57252 29892 57256 29948
rect 57192 29888 57256 29892
rect 2612 29404 2676 29408
rect 2612 29348 2616 29404
rect 2616 29348 2672 29404
rect 2672 29348 2676 29404
rect 2612 29344 2676 29348
rect 2692 29404 2756 29408
rect 2692 29348 2696 29404
rect 2696 29348 2752 29404
rect 2752 29348 2756 29404
rect 2692 29344 2756 29348
rect 2772 29404 2836 29408
rect 2772 29348 2776 29404
rect 2776 29348 2832 29404
rect 2832 29348 2836 29404
rect 2772 29344 2836 29348
rect 2852 29404 2916 29408
rect 2852 29348 2856 29404
rect 2856 29348 2912 29404
rect 2912 29348 2916 29404
rect 2852 29344 2916 29348
rect 7612 29404 7676 29408
rect 7612 29348 7616 29404
rect 7616 29348 7672 29404
rect 7672 29348 7676 29404
rect 7612 29344 7676 29348
rect 7692 29404 7756 29408
rect 7692 29348 7696 29404
rect 7696 29348 7752 29404
rect 7752 29348 7756 29404
rect 7692 29344 7756 29348
rect 7772 29404 7836 29408
rect 7772 29348 7776 29404
rect 7776 29348 7832 29404
rect 7832 29348 7836 29404
rect 7772 29344 7836 29348
rect 7852 29404 7916 29408
rect 7852 29348 7856 29404
rect 7856 29348 7912 29404
rect 7912 29348 7916 29404
rect 7852 29344 7916 29348
rect 12612 29404 12676 29408
rect 12612 29348 12616 29404
rect 12616 29348 12672 29404
rect 12672 29348 12676 29404
rect 12612 29344 12676 29348
rect 12692 29404 12756 29408
rect 12692 29348 12696 29404
rect 12696 29348 12752 29404
rect 12752 29348 12756 29404
rect 12692 29344 12756 29348
rect 12772 29404 12836 29408
rect 12772 29348 12776 29404
rect 12776 29348 12832 29404
rect 12832 29348 12836 29404
rect 12772 29344 12836 29348
rect 12852 29404 12916 29408
rect 12852 29348 12856 29404
rect 12856 29348 12912 29404
rect 12912 29348 12916 29404
rect 12852 29344 12916 29348
rect 17612 29404 17676 29408
rect 17612 29348 17616 29404
rect 17616 29348 17672 29404
rect 17672 29348 17676 29404
rect 17612 29344 17676 29348
rect 17692 29404 17756 29408
rect 17692 29348 17696 29404
rect 17696 29348 17752 29404
rect 17752 29348 17756 29404
rect 17692 29344 17756 29348
rect 17772 29404 17836 29408
rect 17772 29348 17776 29404
rect 17776 29348 17832 29404
rect 17832 29348 17836 29404
rect 17772 29344 17836 29348
rect 17852 29404 17916 29408
rect 17852 29348 17856 29404
rect 17856 29348 17912 29404
rect 17912 29348 17916 29404
rect 17852 29344 17916 29348
rect 22612 29404 22676 29408
rect 22612 29348 22616 29404
rect 22616 29348 22672 29404
rect 22672 29348 22676 29404
rect 22612 29344 22676 29348
rect 22692 29404 22756 29408
rect 22692 29348 22696 29404
rect 22696 29348 22752 29404
rect 22752 29348 22756 29404
rect 22692 29344 22756 29348
rect 22772 29404 22836 29408
rect 22772 29348 22776 29404
rect 22776 29348 22832 29404
rect 22832 29348 22836 29404
rect 22772 29344 22836 29348
rect 22852 29404 22916 29408
rect 22852 29348 22856 29404
rect 22856 29348 22912 29404
rect 22912 29348 22916 29404
rect 22852 29344 22916 29348
rect 27612 29404 27676 29408
rect 27612 29348 27616 29404
rect 27616 29348 27672 29404
rect 27672 29348 27676 29404
rect 27612 29344 27676 29348
rect 27692 29404 27756 29408
rect 27692 29348 27696 29404
rect 27696 29348 27752 29404
rect 27752 29348 27756 29404
rect 27692 29344 27756 29348
rect 27772 29404 27836 29408
rect 27772 29348 27776 29404
rect 27776 29348 27832 29404
rect 27832 29348 27836 29404
rect 27772 29344 27836 29348
rect 27852 29404 27916 29408
rect 27852 29348 27856 29404
rect 27856 29348 27912 29404
rect 27912 29348 27916 29404
rect 27852 29344 27916 29348
rect 32612 29404 32676 29408
rect 32612 29348 32616 29404
rect 32616 29348 32672 29404
rect 32672 29348 32676 29404
rect 32612 29344 32676 29348
rect 32692 29404 32756 29408
rect 32692 29348 32696 29404
rect 32696 29348 32752 29404
rect 32752 29348 32756 29404
rect 32692 29344 32756 29348
rect 32772 29404 32836 29408
rect 32772 29348 32776 29404
rect 32776 29348 32832 29404
rect 32832 29348 32836 29404
rect 32772 29344 32836 29348
rect 32852 29404 32916 29408
rect 32852 29348 32856 29404
rect 32856 29348 32912 29404
rect 32912 29348 32916 29404
rect 32852 29344 32916 29348
rect 37612 29404 37676 29408
rect 37612 29348 37616 29404
rect 37616 29348 37672 29404
rect 37672 29348 37676 29404
rect 37612 29344 37676 29348
rect 37692 29404 37756 29408
rect 37692 29348 37696 29404
rect 37696 29348 37752 29404
rect 37752 29348 37756 29404
rect 37692 29344 37756 29348
rect 37772 29404 37836 29408
rect 37772 29348 37776 29404
rect 37776 29348 37832 29404
rect 37832 29348 37836 29404
rect 37772 29344 37836 29348
rect 37852 29404 37916 29408
rect 37852 29348 37856 29404
rect 37856 29348 37912 29404
rect 37912 29348 37916 29404
rect 37852 29344 37916 29348
rect 42612 29404 42676 29408
rect 42612 29348 42616 29404
rect 42616 29348 42672 29404
rect 42672 29348 42676 29404
rect 42612 29344 42676 29348
rect 42692 29404 42756 29408
rect 42692 29348 42696 29404
rect 42696 29348 42752 29404
rect 42752 29348 42756 29404
rect 42692 29344 42756 29348
rect 42772 29404 42836 29408
rect 42772 29348 42776 29404
rect 42776 29348 42832 29404
rect 42832 29348 42836 29404
rect 42772 29344 42836 29348
rect 42852 29404 42916 29408
rect 42852 29348 42856 29404
rect 42856 29348 42912 29404
rect 42912 29348 42916 29404
rect 42852 29344 42916 29348
rect 47612 29404 47676 29408
rect 47612 29348 47616 29404
rect 47616 29348 47672 29404
rect 47672 29348 47676 29404
rect 47612 29344 47676 29348
rect 47692 29404 47756 29408
rect 47692 29348 47696 29404
rect 47696 29348 47752 29404
rect 47752 29348 47756 29404
rect 47692 29344 47756 29348
rect 47772 29404 47836 29408
rect 47772 29348 47776 29404
rect 47776 29348 47832 29404
rect 47832 29348 47836 29404
rect 47772 29344 47836 29348
rect 47852 29404 47916 29408
rect 47852 29348 47856 29404
rect 47856 29348 47912 29404
rect 47912 29348 47916 29404
rect 47852 29344 47916 29348
rect 52612 29404 52676 29408
rect 52612 29348 52616 29404
rect 52616 29348 52672 29404
rect 52672 29348 52676 29404
rect 52612 29344 52676 29348
rect 52692 29404 52756 29408
rect 52692 29348 52696 29404
rect 52696 29348 52752 29404
rect 52752 29348 52756 29404
rect 52692 29344 52756 29348
rect 52772 29404 52836 29408
rect 52772 29348 52776 29404
rect 52776 29348 52832 29404
rect 52832 29348 52836 29404
rect 52772 29344 52836 29348
rect 52852 29404 52916 29408
rect 52852 29348 52856 29404
rect 52856 29348 52912 29404
rect 52912 29348 52916 29404
rect 52852 29344 52916 29348
rect 57612 29404 57676 29408
rect 57612 29348 57616 29404
rect 57616 29348 57672 29404
rect 57672 29348 57676 29404
rect 57612 29344 57676 29348
rect 57692 29404 57756 29408
rect 57692 29348 57696 29404
rect 57696 29348 57752 29404
rect 57752 29348 57756 29404
rect 57692 29344 57756 29348
rect 57772 29404 57836 29408
rect 57772 29348 57776 29404
rect 57776 29348 57832 29404
rect 57832 29348 57836 29404
rect 57772 29344 57836 29348
rect 57852 29404 57916 29408
rect 57852 29348 57856 29404
rect 57856 29348 57912 29404
rect 57912 29348 57916 29404
rect 57852 29344 57916 29348
rect 1952 28860 2016 28864
rect 1952 28804 1956 28860
rect 1956 28804 2012 28860
rect 2012 28804 2016 28860
rect 1952 28800 2016 28804
rect 2032 28860 2096 28864
rect 2032 28804 2036 28860
rect 2036 28804 2092 28860
rect 2092 28804 2096 28860
rect 2032 28800 2096 28804
rect 2112 28860 2176 28864
rect 2112 28804 2116 28860
rect 2116 28804 2172 28860
rect 2172 28804 2176 28860
rect 2112 28800 2176 28804
rect 2192 28860 2256 28864
rect 2192 28804 2196 28860
rect 2196 28804 2252 28860
rect 2252 28804 2256 28860
rect 2192 28800 2256 28804
rect 6952 28860 7016 28864
rect 6952 28804 6956 28860
rect 6956 28804 7012 28860
rect 7012 28804 7016 28860
rect 6952 28800 7016 28804
rect 7032 28860 7096 28864
rect 7032 28804 7036 28860
rect 7036 28804 7092 28860
rect 7092 28804 7096 28860
rect 7032 28800 7096 28804
rect 7112 28860 7176 28864
rect 7112 28804 7116 28860
rect 7116 28804 7172 28860
rect 7172 28804 7176 28860
rect 7112 28800 7176 28804
rect 7192 28860 7256 28864
rect 7192 28804 7196 28860
rect 7196 28804 7252 28860
rect 7252 28804 7256 28860
rect 7192 28800 7256 28804
rect 11952 28860 12016 28864
rect 11952 28804 11956 28860
rect 11956 28804 12012 28860
rect 12012 28804 12016 28860
rect 11952 28800 12016 28804
rect 12032 28860 12096 28864
rect 12032 28804 12036 28860
rect 12036 28804 12092 28860
rect 12092 28804 12096 28860
rect 12032 28800 12096 28804
rect 12112 28860 12176 28864
rect 12112 28804 12116 28860
rect 12116 28804 12172 28860
rect 12172 28804 12176 28860
rect 12112 28800 12176 28804
rect 12192 28860 12256 28864
rect 12192 28804 12196 28860
rect 12196 28804 12252 28860
rect 12252 28804 12256 28860
rect 12192 28800 12256 28804
rect 16952 28860 17016 28864
rect 16952 28804 16956 28860
rect 16956 28804 17012 28860
rect 17012 28804 17016 28860
rect 16952 28800 17016 28804
rect 17032 28860 17096 28864
rect 17032 28804 17036 28860
rect 17036 28804 17092 28860
rect 17092 28804 17096 28860
rect 17032 28800 17096 28804
rect 17112 28860 17176 28864
rect 17112 28804 17116 28860
rect 17116 28804 17172 28860
rect 17172 28804 17176 28860
rect 17112 28800 17176 28804
rect 17192 28860 17256 28864
rect 17192 28804 17196 28860
rect 17196 28804 17252 28860
rect 17252 28804 17256 28860
rect 17192 28800 17256 28804
rect 21952 28860 22016 28864
rect 21952 28804 21956 28860
rect 21956 28804 22012 28860
rect 22012 28804 22016 28860
rect 21952 28800 22016 28804
rect 22032 28860 22096 28864
rect 22032 28804 22036 28860
rect 22036 28804 22092 28860
rect 22092 28804 22096 28860
rect 22032 28800 22096 28804
rect 22112 28860 22176 28864
rect 22112 28804 22116 28860
rect 22116 28804 22172 28860
rect 22172 28804 22176 28860
rect 22112 28800 22176 28804
rect 22192 28860 22256 28864
rect 22192 28804 22196 28860
rect 22196 28804 22252 28860
rect 22252 28804 22256 28860
rect 22192 28800 22256 28804
rect 26952 28860 27016 28864
rect 26952 28804 26956 28860
rect 26956 28804 27012 28860
rect 27012 28804 27016 28860
rect 26952 28800 27016 28804
rect 27032 28860 27096 28864
rect 27032 28804 27036 28860
rect 27036 28804 27092 28860
rect 27092 28804 27096 28860
rect 27032 28800 27096 28804
rect 27112 28860 27176 28864
rect 27112 28804 27116 28860
rect 27116 28804 27172 28860
rect 27172 28804 27176 28860
rect 27112 28800 27176 28804
rect 27192 28860 27256 28864
rect 27192 28804 27196 28860
rect 27196 28804 27252 28860
rect 27252 28804 27256 28860
rect 27192 28800 27256 28804
rect 31952 28860 32016 28864
rect 31952 28804 31956 28860
rect 31956 28804 32012 28860
rect 32012 28804 32016 28860
rect 31952 28800 32016 28804
rect 32032 28860 32096 28864
rect 32032 28804 32036 28860
rect 32036 28804 32092 28860
rect 32092 28804 32096 28860
rect 32032 28800 32096 28804
rect 32112 28860 32176 28864
rect 32112 28804 32116 28860
rect 32116 28804 32172 28860
rect 32172 28804 32176 28860
rect 32112 28800 32176 28804
rect 32192 28860 32256 28864
rect 32192 28804 32196 28860
rect 32196 28804 32252 28860
rect 32252 28804 32256 28860
rect 32192 28800 32256 28804
rect 36952 28860 37016 28864
rect 36952 28804 36956 28860
rect 36956 28804 37012 28860
rect 37012 28804 37016 28860
rect 36952 28800 37016 28804
rect 37032 28860 37096 28864
rect 37032 28804 37036 28860
rect 37036 28804 37092 28860
rect 37092 28804 37096 28860
rect 37032 28800 37096 28804
rect 37112 28860 37176 28864
rect 37112 28804 37116 28860
rect 37116 28804 37172 28860
rect 37172 28804 37176 28860
rect 37112 28800 37176 28804
rect 37192 28860 37256 28864
rect 37192 28804 37196 28860
rect 37196 28804 37252 28860
rect 37252 28804 37256 28860
rect 37192 28800 37256 28804
rect 41952 28860 42016 28864
rect 41952 28804 41956 28860
rect 41956 28804 42012 28860
rect 42012 28804 42016 28860
rect 41952 28800 42016 28804
rect 42032 28860 42096 28864
rect 42032 28804 42036 28860
rect 42036 28804 42092 28860
rect 42092 28804 42096 28860
rect 42032 28800 42096 28804
rect 42112 28860 42176 28864
rect 42112 28804 42116 28860
rect 42116 28804 42172 28860
rect 42172 28804 42176 28860
rect 42112 28800 42176 28804
rect 42192 28860 42256 28864
rect 42192 28804 42196 28860
rect 42196 28804 42252 28860
rect 42252 28804 42256 28860
rect 42192 28800 42256 28804
rect 46952 28860 47016 28864
rect 46952 28804 46956 28860
rect 46956 28804 47012 28860
rect 47012 28804 47016 28860
rect 46952 28800 47016 28804
rect 47032 28860 47096 28864
rect 47032 28804 47036 28860
rect 47036 28804 47092 28860
rect 47092 28804 47096 28860
rect 47032 28800 47096 28804
rect 47112 28860 47176 28864
rect 47112 28804 47116 28860
rect 47116 28804 47172 28860
rect 47172 28804 47176 28860
rect 47112 28800 47176 28804
rect 47192 28860 47256 28864
rect 47192 28804 47196 28860
rect 47196 28804 47252 28860
rect 47252 28804 47256 28860
rect 47192 28800 47256 28804
rect 51952 28860 52016 28864
rect 51952 28804 51956 28860
rect 51956 28804 52012 28860
rect 52012 28804 52016 28860
rect 51952 28800 52016 28804
rect 52032 28860 52096 28864
rect 52032 28804 52036 28860
rect 52036 28804 52092 28860
rect 52092 28804 52096 28860
rect 52032 28800 52096 28804
rect 52112 28860 52176 28864
rect 52112 28804 52116 28860
rect 52116 28804 52172 28860
rect 52172 28804 52176 28860
rect 52112 28800 52176 28804
rect 52192 28860 52256 28864
rect 52192 28804 52196 28860
rect 52196 28804 52252 28860
rect 52252 28804 52256 28860
rect 52192 28800 52256 28804
rect 56952 28860 57016 28864
rect 56952 28804 56956 28860
rect 56956 28804 57012 28860
rect 57012 28804 57016 28860
rect 56952 28800 57016 28804
rect 57032 28860 57096 28864
rect 57032 28804 57036 28860
rect 57036 28804 57092 28860
rect 57092 28804 57096 28860
rect 57032 28800 57096 28804
rect 57112 28860 57176 28864
rect 57112 28804 57116 28860
rect 57116 28804 57172 28860
rect 57172 28804 57176 28860
rect 57112 28800 57176 28804
rect 57192 28860 57256 28864
rect 57192 28804 57196 28860
rect 57196 28804 57252 28860
rect 57252 28804 57256 28860
rect 57192 28800 57256 28804
rect 2612 28316 2676 28320
rect 2612 28260 2616 28316
rect 2616 28260 2672 28316
rect 2672 28260 2676 28316
rect 2612 28256 2676 28260
rect 2692 28316 2756 28320
rect 2692 28260 2696 28316
rect 2696 28260 2752 28316
rect 2752 28260 2756 28316
rect 2692 28256 2756 28260
rect 2772 28316 2836 28320
rect 2772 28260 2776 28316
rect 2776 28260 2832 28316
rect 2832 28260 2836 28316
rect 2772 28256 2836 28260
rect 2852 28316 2916 28320
rect 2852 28260 2856 28316
rect 2856 28260 2912 28316
rect 2912 28260 2916 28316
rect 2852 28256 2916 28260
rect 7612 28316 7676 28320
rect 7612 28260 7616 28316
rect 7616 28260 7672 28316
rect 7672 28260 7676 28316
rect 7612 28256 7676 28260
rect 7692 28316 7756 28320
rect 7692 28260 7696 28316
rect 7696 28260 7752 28316
rect 7752 28260 7756 28316
rect 7692 28256 7756 28260
rect 7772 28316 7836 28320
rect 7772 28260 7776 28316
rect 7776 28260 7832 28316
rect 7832 28260 7836 28316
rect 7772 28256 7836 28260
rect 7852 28316 7916 28320
rect 7852 28260 7856 28316
rect 7856 28260 7912 28316
rect 7912 28260 7916 28316
rect 7852 28256 7916 28260
rect 12612 28316 12676 28320
rect 12612 28260 12616 28316
rect 12616 28260 12672 28316
rect 12672 28260 12676 28316
rect 12612 28256 12676 28260
rect 12692 28316 12756 28320
rect 12692 28260 12696 28316
rect 12696 28260 12752 28316
rect 12752 28260 12756 28316
rect 12692 28256 12756 28260
rect 12772 28316 12836 28320
rect 12772 28260 12776 28316
rect 12776 28260 12832 28316
rect 12832 28260 12836 28316
rect 12772 28256 12836 28260
rect 12852 28316 12916 28320
rect 12852 28260 12856 28316
rect 12856 28260 12912 28316
rect 12912 28260 12916 28316
rect 12852 28256 12916 28260
rect 17612 28316 17676 28320
rect 17612 28260 17616 28316
rect 17616 28260 17672 28316
rect 17672 28260 17676 28316
rect 17612 28256 17676 28260
rect 17692 28316 17756 28320
rect 17692 28260 17696 28316
rect 17696 28260 17752 28316
rect 17752 28260 17756 28316
rect 17692 28256 17756 28260
rect 17772 28316 17836 28320
rect 17772 28260 17776 28316
rect 17776 28260 17832 28316
rect 17832 28260 17836 28316
rect 17772 28256 17836 28260
rect 17852 28316 17916 28320
rect 17852 28260 17856 28316
rect 17856 28260 17912 28316
rect 17912 28260 17916 28316
rect 17852 28256 17916 28260
rect 22612 28316 22676 28320
rect 22612 28260 22616 28316
rect 22616 28260 22672 28316
rect 22672 28260 22676 28316
rect 22612 28256 22676 28260
rect 22692 28316 22756 28320
rect 22692 28260 22696 28316
rect 22696 28260 22752 28316
rect 22752 28260 22756 28316
rect 22692 28256 22756 28260
rect 22772 28316 22836 28320
rect 22772 28260 22776 28316
rect 22776 28260 22832 28316
rect 22832 28260 22836 28316
rect 22772 28256 22836 28260
rect 22852 28316 22916 28320
rect 22852 28260 22856 28316
rect 22856 28260 22912 28316
rect 22912 28260 22916 28316
rect 22852 28256 22916 28260
rect 27612 28316 27676 28320
rect 27612 28260 27616 28316
rect 27616 28260 27672 28316
rect 27672 28260 27676 28316
rect 27612 28256 27676 28260
rect 27692 28316 27756 28320
rect 27692 28260 27696 28316
rect 27696 28260 27752 28316
rect 27752 28260 27756 28316
rect 27692 28256 27756 28260
rect 27772 28316 27836 28320
rect 27772 28260 27776 28316
rect 27776 28260 27832 28316
rect 27832 28260 27836 28316
rect 27772 28256 27836 28260
rect 27852 28316 27916 28320
rect 27852 28260 27856 28316
rect 27856 28260 27912 28316
rect 27912 28260 27916 28316
rect 27852 28256 27916 28260
rect 32612 28316 32676 28320
rect 32612 28260 32616 28316
rect 32616 28260 32672 28316
rect 32672 28260 32676 28316
rect 32612 28256 32676 28260
rect 32692 28316 32756 28320
rect 32692 28260 32696 28316
rect 32696 28260 32752 28316
rect 32752 28260 32756 28316
rect 32692 28256 32756 28260
rect 32772 28316 32836 28320
rect 32772 28260 32776 28316
rect 32776 28260 32832 28316
rect 32832 28260 32836 28316
rect 32772 28256 32836 28260
rect 32852 28316 32916 28320
rect 32852 28260 32856 28316
rect 32856 28260 32912 28316
rect 32912 28260 32916 28316
rect 32852 28256 32916 28260
rect 37612 28316 37676 28320
rect 37612 28260 37616 28316
rect 37616 28260 37672 28316
rect 37672 28260 37676 28316
rect 37612 28256 37676 28260
rect 37692 28316 37756 28320
rect 37692 28260 37696 28316
rect 37696 28260 37752 28316
rect 37752 28260 37756 28316
rect 37692 28256 37756 28260
rect 37772 28316 37836 28320
rect 37772 28260 37776 28316
rect 37776 28260 37832 28316
rect 37832 28260 37836 28316
rect 37772 28256 37836 28260
rect 37852 28316 37916 28320
rect 37852 28260 37856 28316
rect 37856 28260 37912 28316
rect 37912 28260 37916 28316
rect 37852 28256 37916 28260
rect 42612 28316 42676 28320
rect 42612 28260 42616 28316
rect 42616 28260 42672 28316
rect 42672 28260 42676 28316
rect 42612 28256 42676 28260
rect 42692 28316 42756 28320
rect 42692 28260 42696 28316
rect 42696 28260 42752 28316
rect 42752 28260 42756 28316
rect 42692 28256 42756 28260
rect 42772 28316 42836 28320
rect 42772 28260 42776 28316
rect 42776 28260 42832 28316
rect 42832 28260 42836 28316
rect 42772 28256 42836 28260
rect 42852 28316 42916 28320
rect 42852 28260 42856 28316
rect 42856 28260 42912 28316
rect 42912 28260 42916 28316
rect 42852 28256 42916 28260
rect 47612 28316 47676 28320
rect 47612 28260 47616 28316
rect 47616 28260 47672 28316
rect 47672 28260 47676 28316
rect 47612 28256 47676 28260
rect 47692 28316 47756 28320
rect 47692 28260 47696 28316
rect 47696 28260 47752 28316
rect 47752 28260 47756 28316
rect 47692 28256 47756 28260
rect 47772 28316 47836 28320
rect 47772 28260 47776 28316
rect 47776 28260 47832 28316
rect 47832 28260 47836 28316
rect 47772 28256 47836 28260
rect 47852 28316 47916 28320
rect 47852 28260 47856 28316
rect 47856 28260 47912 28316
rect 47912 28260 47916 28316
rect 47852 28256 47916 28260
rect 52612 28316 52676 28320
rect 52612 28260 52616 28316
rect 52616 28260 52672 28316
rect 52672 28260 52676 28316
rect 52612 28256 52676 28260
rect 52692 28316 52756 28320
rect 52692 28260 52696 28316
rect 52696 28260 52752 28316
rect 52752 28260 52756 28316
rect 52692 28256 52756 28260
rect 52772 28316 52836 28320
rect 52772 28260 52776 28316
rect 52776 28260 52832 28316
rect 52832 28260 52836 28316
rect 52772 28256 52836 28260
rect 52852 28316 52916 28320
rect 52852 28260 52856 28316
rect 52856 28260 52912 28316
rect 52912 28260 52916 28316
rect 52852 28256 52916 28260
rect 57612 28316 57676 28320
rect 57612 28260 57616 28316
rect 57616 28260 57672 28316
rect 57672 28260 57676 28316
rect 57612 28256 57676 28260
rect 57692 28316 57756 28320
rect 57692 28260 57696 28316
rect 57696 28260 57752 28316
rect 57752 28260 57756 28316
rect 57692 28256 57756 28260
rect 57772 28316 57836 28320
rect 57772 28260 57776 28316
rect 57776 28260 57832 28316
rect 57832 28260 57836 28316
rect 57772 28256 57836 28260
rect 57852 28316 57916 28320
rect 57852 28260 57856 28316
rect 57856 28260 57912 28316
rect 57912 28260 57916 28316
rect 57852 28256 57916 28260
rect 1952 27772 2016 27776
rect 1952 27716 1956 27772
rect 1956 27716 2012 27772
rect 2012 27716 2016 27772
rect 1952 27712 2016 27716
rect 2032 27772 2096 27776
rect 2032 27716 2036 27772
rect 2036 27716 2092 27772
rect 2092 27716 2096 27772
rect 2032 27712 2096 27716
rect 2112 27772 2176 27776
rect 2112 27716 2116 27772
rect 2116 27716 2172 27772
rect 2172 27716 2176 27772
rect 2112 27712 2176 27716
rect 2192 27772 2256 27776
rect 2192 27716 2196 27772
rect 2196 27716 2252 27772
rect 2252 27716 2256 27772
rect 2192 27712 2256 27716
rect 6952 27772 7016 27776
rect 6952 27716 6956 27772
rect 6956 27716 7012 27772
rect 7012 27716 7016 27772
rect 6952 27712 7016 27716
rect 7032 27772 7096 27776
rect 7032 27716 7036 27772
rect 7036 27716 7092 27772
rect 7092 27716 7096 27772
rect 7032 27712 7096 27716
rect 7112 27772 7176 27776
rect 7112 27716 7116 27772
rect 7116 27716 7172 27772
rect 7172 27716 7176 27772
rect 7112 27712 7176 27716
rect 7192 27772 7256 27776
rect 7192 27716 7196 27772
rect 7196 27716 7252 27772
rect 7252 27716 7256 27772
rect 7192 27712 7256 27716
rect 11952 27772 12016 27776
rect 11952 27716 11956 27772
rect 11956 27716 12012 27772
rect 12012 27716 12016 27772
rect 11952 27712 12016 27716
rect 12032 27772 12096 27776
rect 12032 27716 12036 27772
rect 12036 27716 12092 27772
rect 12092 27716 12096 27772
rect 12032 27712 12096 27716
rect 12112 27772 12176 27776
rect 12112 27716 12116 27772
rect 12116 27716 12172 27772
rect 12172 27716 12176 27772
rect 12112 27712 12176 27716
rect 12192 27772 12256 27776
rect 12192 27716 12196 27772
rect 12196 27716 12252 27772
rect 12252 27716 12256 27772
rect 12192 27712 12256 27716
rect 16952 27772 17016 27776
rect 16952 27716 16956 27772
rect 16956 27716 17012 27772
rect 17012 27716 17016 27772
rect 16952 27712 17016 27716
rect 17032 27772 17096 27776
rect 17032 27716 17036 27772
rect 17036 27716 17092 27772
rect 17092 27716 17096 27772
rect 17032 27712 17096 27716
rect 17112 27772 17176 27776
rect 17112 27716 17116 27772
rect 17116 27716 17172 27772
rect 17172 27716 17176 27772
rect 17112 27712 17176 27716
rect 17192 27772 17256 27776
rect 17192 27716 17196 27772
rect 17196 27716 17252 27772
rect 17252 27716 17256 27772
rect 17192 27712 17256 27716
rect 21952 27772 22016 27776
rect 21952 27716 21956 27772
rect 21956 27716 22012 27772
rect 22012 27716 22016 27772
rect 21952 27712 22016 27716
rect 22032 27772 22096 27776
rect 22032 27716 22036 27772
rect 22036 27716 22092 27772
rect 22092 27716 22096 27772
rect 22032 27712 22096 27716
rect 22112 27772 22176 27776
rect 22112 27716 22116 27772
rect 22116 27716 22172 27772
rect 22172 27716 22176 27772
rect 22112 27712 22176 27716
rect 22192 27772 22256 27776
rect 22192 27716 22196 27772
rect 22196 27716 22252 27772
rect 22252 27716 22256 27772
rect 22192 27712 22256 27716
rect 26952 27772 27016 27776
rect 26952 27716 26956 27772
rect 26956 27716 27012 27772
rect 27012 27716 27016 27772
rect 26952 27712 27016 27716
rect 27032 27772 27096 27776
rect 27032 27716 27036 27772
rect 27036 27716 27092 27772
rect 27092 27716 27096 27772
rect 27032 27712 27096 27716
rect 27112 27772 27176 27776
rect 27112 27716 27116 27772
rect 27116 27716 27172 27772
rect 27172 27716 27176 27772
rect 27112 27712 27176 27716
rect 27192 27772 27256 27776
rect 27192 27716 27196 27772
rect 27196 27716 27252 27772
rect 27252 27716 27256 27772
rect 27192 27712 27256 27716
rect 31952 27772 32016 27776
rect 31952 27716 31956 27772
rect 31956 27716 32012 27772
rect 32012 27716 32016 27772
rect 31952 27712 32016 27716
rect 32032 27772 32096 27776
rect 32032 27716 32036 27772
rect 32036 27716 32092 27772
rect 32092 27716 32096 27772
rect 32032 27712 32096 27716
rect 32112 27772 32176 27776
rect 32112 27716 32116 27772
rect 32116 27716 32172 27772
rect 32172 27716 32176 27772
rect 32112 27712 32176 27716
rect 32192 27772 32256 27776
rect 32192 27716 32196 27772
rect 32196 27716 32252 27772
rect 32252 27716 32256 27772
rect 32192 27712 32256 27716
rect 36952 27772 37016 27776
rect 36952 27716 36956 27772
rect 36956 27716 37012 27772
rect 37012 27716 37016 27772
rect 36952 27712 37016 27716
rect 37032 27772 37096 27776
rect 37032 27716 37036 27772
rect 37036 27716 37092 27772
rect 37092 27716 37096 27772
rect 37032 27712 37096 27716
rect 37112 27772 37176 27776
rect 37112 27716 37116 27772
rect 37116 27716 37172 27772
rect 37172 27716 37176 27772
rect 37112 27712 37176 27716
rect 37192 27772 37256 27776
rect 37192 27716 37196 27772
rect 37196 27716 37252 27772
rect 37252 27716 37256 27772
rect 37192 27712 37256 27716
rect 41952 27772 42016 27776
rect 41952 27716 41956 27772
rect 41956 27716 42012 27772
rect 42012 27716 42016 27772
rect 41952 27712 42016 27716
rect 42032 27772 42096 27776
rect 42032 27716 42036 27772
rect 42036 27716 42092 27772
rect 42092 27716 42096 27772
rect 42032 27712 42096 27716
rect 42112 27772 42176 27776
rect 42112 27716 42116 27772
rect 42116 27716 42172 27772
rect 42172 27716 42176 27772
rect 42112 27712 42176 27716
rect 42192 27772 42256 27776
rect 42192 27716 42196 27772
rect 42196 27716 42252 27772
rect 42252 27716 42256 27772
rect 42192 27712 42256 27716
rect 46952 27772 47016 27776
rect 46952 27716 46956 27772
rect 46956 27716 47012 27772
rect 47012 27716 47016 27772
rect 46952 27712 47016 27716
rect 47032 27772 47096 27776
rect 47032 27716 47036 27772
rect 47036 27716 47092 27772
rect 47092 27716 47096 27772
rect 47032 27712 47096 27716
rect 47112 27772 47176 27776
rect 47112 27716 47116 27772
rect 47116 27716 47172 27772
rect 47172 27716 47176 27772
rect 47112 27712 47176 27716
rect 47192 27772 47256 27776
rect 47192 27716 47196 27772
rect 47196 27716 47252 27772
rect 47252 27716 47256 27772
rect 47192 27712 47256 27716
rect 51952 27772 52016 27776
rect 51952 27716 51956 27772
rect 51956 27716 52012 27772
rect 52012 27716 52016 27772
rect 51952 27712 52016 27716
rect 52032 27772 52096 27776
rect 52032 27716 52036 27772
rect 52036 27716 52092 27772
rect 52092 27716 52096 27772
rect 52032 27712 52096 27716
rect 52112 27772 52176 27776
rect 52112 27716 52116 27772
rect 52116 27716 52172 27772
rect 52172 27716 52176 27772
rect 52112 27712 52176 27716
rect 52192 27772 52256 27776
rect 52192 27716 52196 27772
rect 52196 27716 52252 27772
rect 52252 27716 52256 27772
rect 52192 27712 52256 27716
rect 56952 27772 57016 27776
rect 56952 27716 56956 27772
rect 56956 27716 57012 27772
rect 57012 27716 57016 27772
rect 56952 27712 57016 27716
rect 57032 27772 57096 27776
rect 57032 27716 57036 27772
rect 57036 27716 57092 27772
rect 57092 27716 57096 27772
rect 57032 27712 57096 27716
rect 57112 27772 57176 27776
rect 57112 27716 57116 27772
rect 57116 27716 57172 27772
rect 57172 27716 57176 27772
rect 57112 27712 57176 27716
rect 57192 27772 57256 27776
rect 57192 27716 57196 27772
rect 57196 27716 57252 27772
rect 57252 27716 57256 27772
rect 57192 27712 57256 27716
rect 2612 27228 2676 27232
rect 2612 27172 2616 27228
rect 2616 27172 2672 27228
rect 2672 27172 2676 27228
rect 2612 27168 2676 27172
rect 2692 27228 2756 27232
rect 2692 27172 2696 27228
rect 2696 27172 2752 27228
rect 2752 27172 2756 27228
rect 2692 27168 2756 27172
rect 2772 27228 2836 27232
rect 2772 27172 2776 27228
rect 2776 27172 2832 27228
rect 2832 27172 2836 27228
rect 2772 27168 2836 27172
rect 2852 27228 2916 27232
rect 2852 27172 2856 27228
rect 2856 27172 2912 27228
rect 2912 27172 2916 27228
rect 2852 27168 2916 27172
rect 7612 27228 7676 27232
rect 7612 27172 7616 27228
rect 7616 27172 7672 27228
rect 7672 27172 7676 27228
rect 7612 27168 7676 27172
rect 7692 27228 7756 27232
rect 7692 27172 7696 27228
rect 7696 27172 7752 27228
rect 7752 27172 7756 27228
rect 7692 27168 7756 27172
rect 7772 27228 7836 27232
rect 7772 27172 7776 27228
rect 7776 27172 7832 27228
rect 7832 27172 7836 27228
rect 7772 27168 7836 27172
rect 7852 27228 7916 27232
rect 7852 27172 7856 27228
rect 7856 27172 7912 27228
rect 7912 27172 7916 27228
rect 7852 27168 7916 27172
rect 12612 27228 12676 27232
rect 12612 27172 12616 27228
rect 12616 27172 12672 27228
rect 12672 27172 12676 27228
rect 12612 27168 12676 27172
rect 12692 27228 12756 27232
rect 12692 27172 12696 27228
rect 12696 27172 12752 27228
rect 12752 27172 12756 27228
rect 12692 27168 12756 27172
rect 12772 27228 12836 27232
rect 12772 27172 12776 27228
rect 12776 27172 12832 27228
rect 12832 27172 12836 27228
rect 12772 27168 12836 27172
rect 12852 27228 12916 27232
rect 12852 27172 12856 27228
rect 12856 27172 12912 27228
rect 12912 27172 12916 27228
rect 12852 27168 12916 27172
rect 17612 27228 17676 27232
rect 17612 27172 17616 27228
rect 17616 27172 17672 27228
rect 17672 27172 17676 27228
rect 17612 27168 17676 27172
rect 17692 27228 17756 27232
rect 17692 27172 17696 27228
rect 17696 27172 17752 27228
rect 17752 27172 17756 27228
rect 17692 27168 17756 27172
rect 17772 27228 17836 27232
rect 17772 27172 17776 27228
rect 17776 27172 17832 27228
rect 17832 27172 17836 27228
rect 17772 27168 17836 27172
rect 17852 27228 17916 27232
rect 17852 27172 17856 27228
rect 17856 27172 17912 27228
rect 17912 27172 17916 27228
rect 17852 27168 17916 27172
rect 22612 27228 22676 27232
rect 22612 27172 22616 27228
rect 22616 27172 22672 27228
rect 22672 27172 22676 27228
rect 22612 27168 22676 27172
rect 22692 27228 22756 27232
rect 22692 27172 22696 27228
rect 22696 27172 22752 27228
rect 22752 27172 22756 27228
rect 22692 27168 22756 27172
rect 22772 27228 22836 27232
rect 22772 27172 22776 27228
rect 22776 27172 22832 27228
rect 22832 27172 22836 27228
rect 22772 27168 22836 27172
rect 22852 27228 22916 27232
rect 22852 27172 22856 27228
rect 22856 27172 22912 27228
rect 22912 27172 22916 27228
rect 22852 27168 22916 27172
rect 27612 27228 27676 27232
rect 27612 27172 27616 27228
rect 27616 27172 27672 27228
rect 27672 27172 27676 27228
rect 27612 27168 27676 27172
rect 27692 27228 27756 27232
rect 27692 27172 27696 27228
rect 27696 27172 27752 27228
rect 27752 27172 27756 27228
rect 27692 27168 27756 27172
rect 27772 27228 27836 27232
rect 27772 27172 27776 27228
rect 27776 27172 27832 27228
rect 27832 27172 27836 27228
rect 27772 27168 27836 27172
rect 27852 27228 27916 27232
rect 27852 27172 27856 27228
rect 27856 27172 27912 27228
rect 27912 27172 27916 27228
rect 27852 27168 27916 27172
rect 32612 27228 32676 27232
rect 32612 27172 32616 27228
rect 32616 27172 32672 27228
rect 32672 27172 32676 27228
rect 32612 27168 32676 27172
rect 32692 27228 32756 27232
rect 32692 27172 32696 27228
rect 32696 27172 32752 27228
rect 32752 27172 32756 27228
rect 32692 27168 32756 27172
rect 32772 27228 32836 27232
rect 32772 27172 32776 27228
rect 32776 27172 32832 27228
rect 32832 27172 32836 27228
rect 32772 27168 32836 27172
rect 32852 27228 32916 27232
rect 32852 27172 32856 27228
rect 32856 27172 32912 27228
rect 32912 27172 32916 27228
rect 32852 27168 32916 27172
rect 37612 27228 37676 27232
rect 37612 27172 37616 27228
rect 37616 27172 37672 27228
rect 37672 27172 37676 27228
rect 37612 27168 37676 27172
rect 37692 27228 37756 27232
rect 37692 27172 37696 27228
rect 37696 27172 37752 27228
rect 37752 27172 37756 27228
rect 37692 27168 37756 27172
rect 37772 27228 37836 27232
rect 37772 27172 37776 27228
rect 37776 27172 37832 27228
rect 37832 27172 37836 27228
rect 37772 27168 37836 27172
rect 37852 27228 37916 27232
rect 37852 27172 37856 27228
rect 37856 27172 37912 27228
rect 37912 27172 37916 27228
rect 37852 27168 37916 27172
rect 42612 27228 42676 27232
rect 42612 27172 42616 27228
rect 42616 27172 42672 27228
rect 42672 27172 42676 27228
rect 42612 27168 42676 27172
rect 42692 27228 42756 27232
rect 42692 27172 42696 27228
rect 42696 27172 42752 27228
rect 42752 27172 42756 27228
rect 42692 27168 42756 27172
rect 42772 27228 42836 27232
rect 42772 27172 42776 27228
rect 42776 27172 42832 27228
rect 42832 27172 42836 27228
rect 42772 27168 42836 27172
rect 42852 27228 42916 27232
rect 42852 27172 42856 27228
rect 42856 27172 42912 27228
rect 42912 27172 42916 27228
rect 42852 27168 42916 27172
rect 47612 27228 47676 27232
rect 47612 27172 47616 27228
rect 47616 27172 47672 27228
rect 47672 27172 47676 27228
rect 47612 27168 47676 27172
rect 47692 27228 47756 27232
rect 47692 27172 47696 27228
rect 47696 27172 47752 27228
rect 47752 27172 47756 27228
rect 47692 27168 47756 27172
rect 47772 27228 47836 27232
rect 47772 27172 47776 27228
rect 47776 27172 47832 27228
rect 47832 27172 47836 27228
rect 47772 27168 47836 27172
rect 47852 27228 47916 27232
rect 47852 27172 47856 27228
rect 47856 27172 47912 27228
rect 47912 27172 47916 27228
rect 47852 27168 47916 27172
rect 52612 27228 52676 27232
rect 52612 27172 52616 27228
rect 52616 27172 52672 27228
rect 52672 27172 52676 27228
rect 52612 27168 52676 27172
rect 52692 27228 52756 27232
rect 52692 27172 52696 27228
rect 52696 27172 52752 27228
rect 52752 27172 52756 27228
rect 52692 27168 52756 27172
rect 52772 27228 52836 27232
rect 52772 27172 52776 27228
rect 52776 27172 52832 27228
rect 52832 27172 52836 27228
rect 52772 27168 52836 27172
rect 52852 27228 52916 27232
rect 52852 27172 52856 27228
rect 52856 27172 52912 27228
rect 52912 27172 52916 27228
rect 52852 27168 52916 27172
rect 57612 27228 57676 27232
rect 57612 27172 57616 27228
rect 57616 27172 57672 27228
rect 57672 27172 57676 27228
rect 57612 27168 57676 27172
rect 57692 27228 57756 27232
rect 57692 27172 57696 27228
rect 57696 27172 57752 27228
rect 57752 27172 57756 27228
rect 57692 27168 57756 27172
rect 57772 27228 57836 27232
rect 57772 27172 57776 27228
rect 57776 27172 57832 27228
rect 57832 27172 57836 27228
rect 57772 27168 57836 27172
rect 57852 27228 57916 27232
rect 57852 27172 57856 27228
rect 57856 27172 57912 27228
rect 57912 27172 57916 27228
rect 57852 27168 57916 27172
rect 1952 26684 2016 26688
rect 1952 26628 1956 26684
rect 1956 26628 2012 26684
rect 2012 26628 2016 26684
rect 1952 26624 2016 26628
rect 2032 26684 2096 26688
rect 2032 26628 2036 26684
rect 2036 26628 2092 26684
rect 2092 26628 2096 26684
rect 2032 26624 2096 26628
rect 2112 26684 2176 26688
rect 2112 26628 2116 26684
rect 2116 26628 2172 26684
rect 2172 26628 2176 26684
rect 2112 26624 2176 26628
rect 2192 26684 2256 26688
rect 2192 26628 2196 26684
rect 2196 26628 2252 26684
rect 2252 26628 2256 26684
rect 2192 26624 2256 26628
rect 6952 26684 7016 26688
rect 6952 26628 6956 26684
rect 6956 26628 7012 26684
rect 7012 26628 7016 26684
rect 6952 26624 7016 26628
rect 7032 26684 7096 26688
rect 7032 26628 7036 26684
rect 7036 26628 7092 26684
rect 7092 26628 7096 26684
rect 7032 26624 7096 26628
rect 7112 26684 7176 26688
rect 7112 26628 7116 26684
rect 7116 26628 7172 26684
rect 7172 26628 7176 26684
rect 7112 26624 7176 26628
rect 7192 26684 7256 26688
rect 7192 26628 7196 26684
rect 7196 26628 7252 26684
rect 7252 26628 7256 26684
rect 7192 26624 7256 26628
rect 11952 26684 12016 26688
rect 11952 26628 11956 26684
rect 11956 26628 12012 26684
rect 12012 26628 12016 26684
rect 11952 26624 12016 26628
rect 12032 26684 12096 26688
rect 12032 26628 12036 26684
rect 12036 26628 12092 26684
rect 12092 26628 12096 26684
rect 12032 26624 12096 26628
rect 12112 26684 12176 26688
rect 12112 26628 12116 26684
rect 12116 26628 12172 26684
rect 12172 26628 12176 26684
rect 12112 26624 12176 26628
rect 12192 26684 12256 26688
rect 12192 26628 12196 26684
rect 12196 26628 12252 26684
rect 12252 26628 12256 26684
rect 12192 26624 12256 26628
rect 16952 26684 17016 26688
rect 16952 26628 16956 26684
rect 16956 26628 17012 26684
rect 17012 26628 17016 26684
rect 16952 26624 17016 26628
rect 17032 26684 17096 26688
rect 17032 26628 17036 26684
rect 17036 26628 17092 26684
rect 17092 26628 17096 26684
rect 17032 26624 17096 26628
rect 17112 26684 17176 26688
rect 17112 26628 17116 26684
rect 17116 26628 17172 26684
rect 17172 26628 17176 26684
rect 17112 26624 17176 26628
rect 17192 26684 17256 26688
rect 17192 26628 17196 26684
rect 17196 26628 17252 26684
rect 17252 26628 17256 26684
rect 17192 26624 17256 26628
rect 21952 26684 22016 26688
rect 21952 26628 21956 26684
rect 21956 26628 22012 26684
rect 22012 26628 22016 26684
rect 21952 26624 22016 26628
rect 22032 26684 22096 26688
rect 22032 26628 22036 26684
rect 22036 26628 22092 26684
rect 22092 26628 22096 26684
rect 22032 26624 22096 26628
rect 22112 26684 22176 26688
rect 22112 26628 22116 26684
rect 22116 26628 22172 26684
rect 22172 26628 22176 26684
rect 22112 26624 22176 26628
rect 22192 26684 22256 26688
rect 22192 26628 22196 26684
rect 22196 26628 22252 26684
rect 22252 26628 22256 26684
rect 22192 26624 22256 26628
rect 26952 26684 27016 26688
rect 26952 26628 26956 26684
rect 26956 26628 27012 26684
rect 27012 26628 27016 26684
rect 26952 26624 27016 26628
rect 27032 26684 27096 26688
rect 27032 26628 27036 26684
rect 27036 26628 27092 26684
rect 27092 26628 27096 26684
rect 27032 26624 27096 26628
rect 27112 26684 27176 26688
rect 27112 26628 27116 26684
rect 27116 26628 27172 26684
rect 27172 26628 27176 26684
rect 27112 26624 27176 26628
rect 27192 26684 27256 26688
rect 27192 26628 27196 26684
rect 27196 26628 27252 26684
rect 27252 26628 27256 26684
rect 27192 26624 27256 26628
rect 31952 26684 32016 26688
rect 31952 26628 31956 26684
rect 31956 26628 32012 26684
rect 32012 26628 32016 26684
rect 31952 26624 32016 26628
rect 32032 26684 32096 26688
rect 32032 26628 32036 26684
rect 32036 26628 32092 26684
rect 32092 26628 32096 26684
rect 32032 26624 32096 26628
rect 32112 26684 32176 26688
rect 32112 26628 32116 26684
rect 32116 26628 32172 26684
rect 32172 26628 32176 26684
rect 32112 26624 32176 26628
rect 32192 26684 32256 26688
rect 32192 26628 32196 26684
rect 32196 26628 32252 26684
rect 32252 26628 32256 26684
rect 32192 26624 32256 26628
rect 36952 26684 37016 26688
rect 36952 26628 36956 26684
rect 36956 26628 37012 26684
rect 37012 26628 37016 26684
rect 36952 26624 37016 26628
rect 37032 26684 37096 26688
rect 37032 26628 37036 26684
rect 37036 26628 37092 26684
rect 37092 26628 37096 26684
rect 37032 26624 37096 26628
rect 37112 26684 37176 26688
rect 37112 26628 37116 26684
rect 37116 26628 37172 26684
rect 37172 26628 37176 26684
rect 37112 26624 37176 26628
rect 37192 26684 37256 26688
rect 37192 26628 37196 26684
rect 37196 26628 37252 26684
rect 37252 26628 37256 26684
rect 37192 26624 37256 26628
rect 41952 26684 42016 26688
rect 41952 26628 41956 26684
rect 41956 26628 42012 26684
rect 42012 26628 42016 26684
rect 41952 26624 42016 26628
rect 42032 26684 42096 26688
rect 42032 26628 42036 26684
rect 42036 26628 42092 26684
rect 42092 26628 42096 26684
rect 42032 26624 42096 26628
rect 42112 26684 42176 26688
rect 42112 26628 42116 26684
rect 42116 26628 42172 26684
rect 42172 26628 42176 26684
rect 42112 26624 42176 26628
rect 42192 26684 42256 26688
rect 42192 26628 42196 26684
rect 42196 26628 42252 26684
rect 42252 26628 42256 26684
rect 42192 26624 42256 26628
rect 46952 26684 47016 26688
rect 46952 26628 46956 26684
rect 46956 26628 47012 26684
rect 47012 26628 47016 26684
rect 46952 26624 47016 26628
rect 47032 26684 47096 26688
rect 47032 26628 47036 26684
rect 47036 26628 47092 26684
rect 47092 26628 47096 26684
rect 47032 26624 47096 26628
rect 47112 26684 47176 26688
rect 47112 26628 47116 26684
rect 47116 26628 47172 26684
rect 47172 26628 47176 26684
rect 47112 26624 47176 26628
rect 47192 26684 47256 26688
rect 47192 26628 47196 26684
rect 47196 26628 47252 26684
rect 47252 26628 47256 26684
rect 47192 26624 47256 26628
rect 51952 26684 52016 26688
rect 51952 26628 51956 26684
rect 51956 26628 52012 26684
rect 52012 26628 52016 26684
rect 51952 26624 52016 26628
rect 52032 26684 52096 26688
rect 52032 26628 52036 26684
rect 52036 26628 52092 26684
rect 52092 26628 52096 26684
rect 52032 26624 52096 26628
rect 52112 26684 52176 26688
rect 52112 26628 52116 26684
rect 52116 26628 52172 26684
rect 52172 26628 52176 26684
rect 52112 26624 52176 26628
rect 52192 26684 52256 26688
rect 52192 26628 52196 26684
rect 52196 26628 52252 26684
rect 52252 26628 52256 26684
rect 52192 26624 52256 26628
rect 56952 26684 57016 26688
rect 56952 26628 56956 26684
rect 56956 26628 57012 26684
rect 57012 26628 57016 26684
rect 56952 26624 57016 26628
rect 57032 26684 57096 26688
rect 57032 26628 57036 26684
rect 57036 26628 57092 26684
rect 57092 26628 57096 26684
rect 57032 26624 57096 26628
rect 57112 26684 57176 26688
rect 57112 26628 57116 26684
rect 57116 26628 57172 26684
rect 57172 26628 57176 26684
rect 57112 26624 57176 26628
rect 57192 26684 57256 26688
rect 57192 26628 57196 26684
rect 57196 26628 57252 26684
rect 57252 26628 57256 26684
rect 57192 26624 57256 26628
rect 2612 26140 2676 26144
rect 2612 26084 2616 26140
rect 2616 26084 2672 26140
rect 2672 26084 2676 26140
rect 2612 26080 2676 26084
rect 2692 26140 2756 26144
rect 2692 26084 2696 26140
rect 2696 26084 2752 26140
rect 2752 26084 2756 26140
rect 2692 26080 2756 26084
rect 2772 26140 2836 26144
rect 2772 26084 2776 26140
rect 2776 26084 2832 26140
rect 2832 26084 2836 26140
rect 2772 26080 2836 26084
rect 2852 26140 2916 26144
rect 2852 26084 2856 26140
rect 2856 26084 2912 26140
rect 2912 26084 2916 26140
rect 2852 26080 2916 26084
rect 7612 26140 7676 26144
rect 7612 26084 7616 26140
rect 7616 26084 7672 26140
rect 7672 26084 7676 26140
rect 7612 26080 7676 26084
rect 7692 26140 7756 26144
rect 7692 26084 7696 26140
rect 7696 26084 7752 26140
rect 7752 26084 7756 26140
rect 7692 26080 7756 26084
rect 7772 26140 7836 26144
rect 7772 26084 7776 26140
rect 7776 26084 7832 26140
rect 7832 26084 7836 26140
rect 7772 26080 7836 26084
rect 7852 26140 7916 26144
rect 7852 26084 7856 26140
rect 7856 26084 7912 26140
rect 7912 26084 7916 26140
rect 7852 26080 7916 26084
rect 12612 26140 12676 26144
rect 12612 26084 12616 26140
rect 12616 26084 12672 26140
rect 12672 26084 12676 26140
rect 12612 26080 12676 26084
rect 12692 26140 12756 26144
rect 12692 26084 12696 26140
rect 12696 26084 12752 26140
rect 12752 26084 12756 26140
rect 12692 26080 12756 26084
rect 12772 26140 12836 26144
rect 12772 26084 12776 26140
rect 12776 26084 12832 26140
rect 12832 26084 12836 26140
rect 12772 26080 12836 26084
rect 12852 26140 12916 26144
rect 12852 26084 12856 26140
rect 12856 26084 12912 26140
rect 12912 26084 12916 26140
rect 12852 26080 12916 26084
rect 17612 26140 17676 26144
rect 17612 26084 17616 26140
rect 17616 26084 17672 26140
rect 17672 26084 17676 26140
rect 17612 26080 17676 26084
rect 17692 26140 17756 26144
rect 17692 26084 17696 26140
rect 17696 26084 17752 26140
rect 17752 26084 17756 26140
rect 17692 26080 17756 26084
rect 17772 26140 17836 26144
rect 17772 26084 17776 26140
rect 17776 26084 17832 26140
rect 17832 26084 17836 26140
rect 17772 26080 17836 26084
rect 17852 26140 17916 26144
rect 17852 26084 17856 26140
rect 17856 26084 17912 26140
rect 17912 26084 17916 26140
rect 17852 26080 17916 26084
rect 22612 26140 22676 26144
rect 22612 26084 22616 26140
rect 22616 26084 22672 26140
rect 22672 26084 22676 26140
rect 22612 26080 22676 26084
rect 22692 26140 22756 26144
rect 22692 26084 22696 26140
rect 22696 26084 22752 26140
rect 22752 26084 22756 26140
rect 22692 26080 22756 26084
rect 22772 26140 22836 26144
rect 22772 26084 22776 26140
rect 22776 26084 22832 26140
rect 22832 26084 22836 26140
rect 22772 26080 22836 26084
rect 22852 26140 22916 26144
rect 22852 26084 22856 26140
rect 22856 26084 22912 26140
rect 22912 26084 22916 26140
rect 22852 26080 22916 26084
rect 27612 26140 27676 26144
rect 27612 26084 27616 26140
rect 27616 26084 27672 26140
rect 27672 26084 27676 26140
rect 27612 26080 27676 26084
rect 27692 26140 27756 26144
rect 27692 26084 27696 26140
rect 27696 26084 27752 26140
rect 27752 26084 27756 26140
rect 27692 26080 27756 26084
rect 27772 26140 27836 26144
rect 27772 26084 27776 26140
rect 27776 26084 27832 26140
rect 27832 26084 27836 26140
rect 27772 26080 27836 26084
rect 27852 26140 27916 26144
rect 27852 26084 27856 26140
rect 27856 26084 27912 26140
rect 27912 26084 27916 26140
rect 27852 26080 27916 26084
rect 32612 26140 32676 26144
rect 32612 26084 32616 26140
rect 32616 26084 32672 26140
rect 32672 26084 32676 26140
rect 32612 26080 32676 26084
rect 32692 26140 32756 26144
rect 32692 26084 32696 26140
rect 32696 26084 32752 26140
rect 32752 26084 32756 26140
rect 32692 26080 32756 26084
rect 32772 26140 32836 26144
rect 32772 26084 32776 26140
rect 32776 26084 32832 26140
rect 32832 26084 32836 26140
rect 32772 26080 32836 26084
rect 32852 26140 32916 26144
rect 32852 26084 32856 26140
rect 32856 26084 32912 26140
rect 32912 26084 32916 26140
rect 32852 26080 32916 26084
rect 37612 26140 37676 26144
rect 37612 26084 37616 26140
rect 37616 26084 37672 26140
rect 37672 26084 37676 26140
rect 37612 26080 37676 26084
rect 37692 26140 37756 26144
rect 37692 26084 37696 26140
rect 37696 26084 37752 26140
rect 37752 26084 37756 26140
rect 37692 26080 37756 26084
rect 37772 26140 37836 26144
rect 37772 26084 37776 26140
rect 37776 26084 37832 26140
rect 37832 26084 37836 26140
rect 37772 26080 37836 26084
rect 37852 26140 37916 26144
rect 37852 26084 37856 26140
rect 37856 26084 37912 26140
rect 37912 26084 37916 26140
rect 37852 26080 37916 26084
rect 42612 26140 42676 26144
rect 42612 26084 42616 26140
rect 42616 26084 42672 26140
rect 42672 26084 42676 26140
rect 42612 26080 42676 26084
rect 42692 26140 42756 26144
rect 42692 26084 42696 26140
rect 42696 26084 42752 26140
rect 42752 26084 42756 26140
rect 42692 26080 42756 26084
rect 42772 26140 42836 26144
rect 42772 26084 42776 26140
rect 42776 26084 42832 26140
rect 42832 26084 42836 26140
rect 42772 26080 42836 26084
rect 42852 26140 42916 26144
rect 42852 26084 42856 26140
rect 42856 26084 42912 26140
rect 42912 26084 42916 26140
rect 42852 26080 42916 26084
rect 47612 26140 47676 26144
rect 47612 26084 47616 26140
rect 47616 26084 47672 26140
rect 47672 26084 47676 26140
rect 47612 26080 47676 26084
rect 47692 26140 47756 26144
rect 47692 26084 47696 26140
rect 47696 26084 47752 26140
rect 47752 26084 47756 26140
rect 47692 26080 47756 26084
rect 47772 26140 47836 26144
rect 47772 26084 47776 26140
rect 47776 26084 47832 26140
rect 47832 26084 47836 26140
rect 47772 26080 47836 26084
rect 47852 26140 47916 26144
rect 47852 26084 47856 26140
rect 47856 26084 47912 26140
rect 47912 26084 47916 26140
rect 47852 26080 47916 26084
rect 52612 26140 52676 26144
rect 52612 26084 52616 26140
rect 52616 26084 52672 26140
rect 52672 26084 52676 26140
rect 52612 26080 52676 26084
rect 52692 26140 52756 26144
rect 52692 26084 52696 26140
rect 52696 26084 52752 26140
rect 52752 26084 52756 26140
rect 52692 26080 52756 26084
rect 52772 26140 52836 26144
rect 52772 26084 52776 26140
rect 52776 26084 52832 26140
rect 52832 26084 52836 26140
rect 52772 26080 52836 26084
rect 52852 26140 52916 26144
rect 52852 26084 52856 26140
rect 52856 26084 52912 26140
rect 52912 26084 52916 26140
rect 52852 26080 52916 26084
rect 57612 26140 57676 26144
rect 57612 26084 57616 26140
rect 57616 26084 57672 26140
rect 57672 26084 57676 26140
rect 57612 26080 57676 26084
rect 57692 26140 57756 26144
rect 57692 26084 57696 26140
rect 57696 26084 57752 26140
rect 57752 26084 57756 26140
rect 57692 26080 57756 26084
rect 57772 26140 57836 26144
rect 57772 26084 57776 26140
rect 57776 26084 57832 26140
rect 57832 26084 57836 26140
rect 57772 26080 57836 26084
rect 57852 26140 57916 26144
rect 57852 26084 57856 26140
rect 57856 26084 57912 26140
rect 57912 26084 57916 26140
rect 57852 26080 57916 26084
rect 1952 25596 2016 25600
rect 1952 25540 1956 25596
rect 1956 25540 2012 25596
rect 2012 25540 2016 25596
rect 1952 25536 2016 25540
rect 2032 25596 2096 25600
rect 2032 25540 2036 25596
rect 2036 25540 2092 25596
rect 2092 25540 2096 25596
rect 2032 25536 2096 25540
rect 2112 25596 2176 25600
rect 2112 25540 2116 25596
rect 2116 25540 2172 25596
rect 2172 25540 2176 25596
rect 2112 25536 2176 25540
rect 2192 25596 2256 25600
rect 2192 25540 2196 25596
rect 2196 25540 2252 25596
rect 2252 25540 2256 25596
rect 2192 25536 2256 25540
rect 6952 25596 7016 25600
rect 6952 25540 6956 25596
rect 6956 25540 7012 25596
rect 7012 25540 7016 25596
rect 6952 25536 7016 25540
rect 7032 25596 7096 25600
rect 7032 25540 7036 25596
rect 7036 25540 7092 25596
rect 7092 25540 7096 25596
rect 7032 25536 7096 25540
rect 7112 25596 7176 25600
rect 7112 25540 7116 25596
rect 7116 25540 7172 25596
rect 7172 25540 7176 25596
rect 7112 25536 7176 25540
rect 7192 25596 7256 25600
rect 7192 25540 7196 25596
rect 7196 25540 7252 25596
rect 7252 25540 7256 25596
rect 7192 25536 7256 25540
rect 11952 25596 12016 25600
rect 11952 25540 11956 25596
rect 11956 25540 12012 25596
rect 12012 25540 12016 25596
rect 11952 25536 12016 25540
rect 12032 25596 12096 25600
rect 12032 25540 12036 25596
rect 12036 25540 12092 25596
rect 12092 25540 12096 25596
rect 12032 25536 12096 25540
rect 12112 25596 12176 25600
rect 12112 25540 12116 25596
rect 12116 25540 12172 25596
rect 12172 25540 12176 25596
rect 12112 25536 12176 25540
rect 12192 25596 12256 25600
rect 12192 25540 12196 25596
rect 12196 25540 12252 25596
rect 12252 25540 12256 25596
rect 12192 25536 12256 25540
rect 16952 25596 17016 25600
rect 16952 25540 16956 25596
rect 16956 25540 17012 25596
rect 17012 25540 17016 25596
rect 16952 25536 17016 25540
rect 17032 25596 17096 25600
rect 17032 25540 17036 25596
rect 17036 25540 17092 25596
rect 17092 25540 17096 25596
rect 17032 25536 17096 25540
rect 17112 25596 17176 25600
rect 17112 25540 17116 25596
rect 17116 25540 17172 25596
rect 17172 25540 17176 25596
rect 17112 25536 17176 25540
rect 17192 25596 17256 25600
rect 17192 25540 17196 25596
rect 17196 25540 17252 25596
rect 17252 25540 17256 25596
rect 17192 25536 17256 25540
rect 21952 25596 22016 25600
rect 21952 25540 21956 25596
rect 21956 25540 22012 25596
rect 22012 25540 22016 25596
rect 21952 25536 22016 25540
rect 22032 25596 22096 25600
rect 22032 25540 22036 25596
rect 22036 25540 22092 25596
rect 22092 25540 22096 25596
rect 22032 25536 22096 25540
rect 22112 25596 22176 25600
rect 22112 25540 22116 25596
rect 22116 25540 22172 25596
rect 22172 25540 22176 25596
rect 22112 25536 22176 25540
rect 22192 25596 22256 25600
rect 22192 25540 22196 25596
rect 22196 25540 22252 25596
rect 22252 25540 22256 25596
rect 22192 25536 22256 25540
rect 26952 25596 27016 25600
rect 26952 25540 26956 25596
rect 26956 25540 27012 25596
rect 27012 25540 27016 25596
rect 26952 25536 27016 25540
rect 27032 25596 27096 25600
rect 27032 25540 27036 25596
rect 27036 25540 27092 25596
rect 27092 25540 27096 25596
rect 27032 25536 27096 25540
rect 27112 25596 27176 25600
rect 27112 25540 27116 25596
rect 27116 25540 27172 25596
rect 27172 25540 27176 25596
rect 27112 25536 27176 25540
rect 27192 25596 27256 25600
rect 27192 25540 27196 25596
rect 27196 25540 27252 25596
rect 27252 25540 27256 25596
rect 27192 25536 27256 25540
rect 31952 25596 32016 25600
rect 31952 25540 31956 25596
rect 31956 25540 32012 25596
rect 32012 25540 32016 25596
rect 31952 25536 32016 25540
rect 32032 25596 32096 25600
rect 32032 25540 32036 25596
rect 32036 25540 32092 25596
rect 32092 25540 32096 25596
rect 32032 25536 32096 25540
rect 32112 25596 32176 25600
rect 32112 25540 32116 25596
rect 32116 25540 32172 25596
rect 32172 25540 32176 25596
rect 32112 25536 32176 25540
rect 32192 25596 32256 25600
rect 32192 25540 32196 25596
rect 32196 25540 32252 25596
rect 32252 25540 32256 25596
rect 32192 25536 32256 25540
rect 36952 25596 37016 25600
rect 36952 25540 36956 25596
rect 36956 25540 37012 25596
rect 37012 25540 37016 25596
rect 36952 25536 37016 25540
rect 37032 25596 37096 25600
rect 37032 25540 37036 25596
rect 37036 25540 37092 25596
rect 37092 25540 37096 25596
rect 37032 25536 37096 25540
rect 37112 25596 37176 25600
rect 37112 25540 37116 25596
rect 37116 25540 37172 25596
rect 37172 25540 37176 25596
rect 37112 25536 37176 25540
rect 37192 25596 37256 25600
rect 37192 25540 37196 25596
rect 37196 25540 37252 25596
rect 37252 25540 37256 25596
rect 37192 25536 37256 25540
rect 41952 25596 42016 25600
rect 41952 25540 41956 25596
rect 41956 25540 42012 25596
rect 42012 25540 42016 25596
rect 41952 25536 42016 25540
rect 42032 25596 42096 25600
rect 42032 25540 42036 25596
rect 42036 25540 42092 25596
rect 42092 25540 42096 25596
rect 42032 25536 42096 25540
rect 42112 25596 42176 25600
rect 42112 25540 42116 25596
rect 42116 25540 42172 25596
rect 42172 25540 42176 25596
rect 42112 25536 42176 25540
rect 42192 25596 42256 25600
rect 42192 25540 42196 25596
rect 42196 25540 42252 25596
rect 42252 25540 42256 25596
rect 42192 25536 42256 25540
rect 46952 25596 47016 25600
rect 46952 25540 46956 25596
rect 46956 25540 47012 25596
rect 47012 25540 47016 25596
rect 46952 25536 47016 25540
rect 47032 25596 47096 25600
rect 47032 25540 47036 25596
rect 47036 25540 47092 25596
rect 47092 25540 47096 25596
rect 47032 25536 47096 25540
rect 47112 25596 47176 25600
rect 47112 25540 47116 25596
rect 47116 25540 47172 25596
rect 47172 25540 47176 25596
rect 47112 25536 47176 25540
rect 47192 25596 47256 25600
rect 47192 25540 47196 25596
rect 47196 25540 47252 25596
rect 47252 25540 47256 25596
rect 47192 25536 47256 25540
rect 51952 25596 52016 25600
rect 51952 25540 51956 25596
rect 51956 25540 52012 25596
rect 52012 25540 52016 25596
rect 51952 25536 52016 25540
rect 52032 25596 52096 25600
rect 52032 25540 52036 25596
rect 52036 25540 52092 25596
rect 52092 25540 52096 25596
rect 52032 25536 52096 25540
rect 52112 25596 52176 25600
rect 52112 25540 52116 25596
rect 52116 25540 52172 25596
rect 52172 25540 52176 25596
rect 52112 25536 52176 25540
rect 52192 25596 52256 25600
rect 52192 25540 52196 25596
rect 52196 25540 52252 25596
rect 52252 25540 52256 25596
rect 52192 25536 52256 25540
rect 56952 25596 57016 25600
rect 56952 25540 56956 25596
rect 56956 25540 57012 25596
rect 57012 25540 57016 25596
rect 56952 25536 57016 25540
rect 57032 25596 57096 25600
rect 57032 25540 57036 25596
rect 57036 25540 57092 25596
rect 57092 25540 57096 25596
rect 57032 25536 57096 25540
rect 57112 25596 57176 25600
rect 57112 25540 57116 25596
rect 57116 25540 57172 25596
rect 57172 25540 57176 25596
rect 57112 25536 57176 25540
rect 57192 25596 57256 25600
rect 57192 25540 57196 25596
rect 57196 25540 57252 25596
rect 57252 25540 57256 25596
rect 57192 25536 57256 25540
rect 2612 25052 2676 25056
rect 2612 24996 2616 25052
rect 2616 24996 2672 25052
rect 2672 24996 2676 25052
rect 2612 24992 2676 24996
rect 2692 25052 2756 25056
rect 2692 24996 2696 25052
rect 2696 24996 2752 25052
rect 2752 24996 2756 25052
rect 2692 24992 2756 24996
rect 2772 25052 2836 25056
rect 2772 24996 2776 25052
rect 2776 24996 2832 25052
rect 2832 24996 2836 25052
rect 2772 24992 2836 24996
rect 2852 25052 2916 25056
rect 2852 24996 2856 25052
rect 2856 24996 2912 25052
rect 2912 24996 2916 25052
rect 2852 24992 2916 24996
rect 7612 25052 7676 25056
rect 7612 24996 7616 25052
rect 7616 24996 7672 25052
rect 7672 24996 7676 25052
rect 7612 24992 7676 24996
rect 7692 25052 7756 25056
rect 7692 24996 7696 25052
rect 7696 24996 7752 25052
rect 7752 24996 7756 25052
rect 7692 24992 7756 24996
rect 7772 25052 7836 25056
rect 7772 24996 7776 25052
rect 7776 24996 7832 25052
rect 7832 24996 7836 25052
rect 7772 24992 7836 24996
rect 7852 25052 7916 25056
rect 7852 24996 7856 25052
rect 7856 24996 7912 25052
rect 7912 24996 7916 25052
rect 7852 24992 7916 24996
rect 12612 25052 12676 25056
rect 12612 24996 12616 25052
rect 12616 24996 12672 25052
rect 12672 24996 12676 25052
rect 12612 24992 12676 24996
rect 12692 25052 12756 25056
rect 12692 24996 12696 25052
rect 12696 24996 12752 25052
rect 12752 24996 12756 25052
rect 12692 24992 12756 24996
rect 12772 25052 12836 25056
rect 12772 24996 12776 25052
rect 12776 24996 12832 25052
rect 12832 24996 12836 25052
rect 12772 24992 12836 24996
rect 12852 25052 12916 25056
rect 12852 24996 12856 25052
rect 12856 24996 12912 25052
rect 12912 24996 12916 25052
rect 12852 24992 12916 24996
rect 17612 25052 17676 25056
rect 17612 24996 17616 25052
rect 17616 24996 17672 25052
rect 17672 24996 17676 25052
rect 17612 24992 17676 24996
rect 17692 25052 17756 25056
rect 17692 24996 17696 25052
rect 17696 24996 17752 25052
rect 17752 24996 17756 25052
rect 17692 24992 17756 24996
rect 17772 25052 17836 25056
rect 17772 24996 17776 25052
rect 17776 24996 17832 25052
rect 17832 24996 17836 25052
rect 17772 24992 17836 24996
rect 17852 25052 17916 25056
rect 17852 24996 17856 25052
rect 17856 24996 17912 25052
rect 17912 24996 17916 25052
rect 17852 24992 17916 24996
rect 22612 25052 22676 25056
rect 22612 24996 22616 25052
rect 22616 24996 22672 25052
rect 22672 24996 22676 25052
rect 22612 24992 22676 24996
rect 22692 25052 22756 25056
rect 22692 24996 22696 25052
rect 22696 24996 22752 25052
rect 22752 24996 22756 25052
rect 22692 24992 22756 24996
rect 22772 25052 22836 25056
rect 22772 24996 22776 25052
rect 22776 24996 22832 25052
rect 22832 24996 22836 25052
rect 22772 24992 22836 24996
rect 22852 25052 22916 25056
rect 22852 24996 22856 25052
rect 22856 24996 22912 25052
rect 22912 24996 22916 25052
rect 22852 24992 22916 24996
rect 27612 25052 27676 25056
rect 27612 24996 27616 25052
rect 27616 24996 27672 25052
rect 27672 24996 27676 25052
rect 27612 24992 27676 24996
rect 27692 25052 27756 25056
rect 27692 24996 27696 25052
rect 27696 24996 27752 25052
rect 27752 24996 27756 25052
rect 27692 24992 27756 24996
rect 27772 25052 27836 25056
rect 27772 24996 27776 25052
rect 27776 24996 27832 25052
rect 27832 24996 27836 25052
rect 27772 24992 27836 24996
rect 27852 25052 27916 25056
rect 27852 24996 27856 25052
rect 27856 24996 27912 25052
rect 27912 24996 27916 25052
rect 27852 24992 27916 24996
rect 32612 25052 32676 25056
rect 32612 24996 32616 25052
rect 32616 24996 32672 25052
rect 32672 24996 32676 25052
rect 32612 24992 32676 24996
rect 32692 25052 32756 25056
rect 32692 24996 32696 25052
rect 32696 24996 32752 25052
rect 32752 24996 32756 25052
rect 32692 24992 32756 24996
rect 32772 25052 32836 25056
rect 32772 24996 32776 25052
rect 32776 24996 32832 25052
rect 32832 24996 32836 25052
rect 32772 24992 32836 24996
rect 32852 25052 32916 25056
rect 32852 24996 32856 25052
rect 32856 24996 32912 25052
rect 32912 24996 32916 25052
rect 32852 24992 32916 24996
rect 37612 25052 37676 25056
rect 37612 24996 37616 25052
rect 37616 24996 37672 25052
rect 37672 24996 37676 25052
rect 37612 24992 37676 24996
rect 37692 25052 37756 25056
rect 37692 24996 37696 25052
rect 37696 24996 37752 25052
rect 37752 24996 37756 25052
rect 37692 24992 37756 24996
rect 37772 25052 37836 25056
rect 37772 24996 37776 25052
rect 37776 24996 37832 25052
rect 37832 24996 37836 25052
rect 37772 24992 37836 24996
rect 37852 25052 37916 25056
rect 37852 24996 37856 25052
rect 37856 24996 37912 25052
rect 37912 24996 37916 25052
rect 37852 24992 37916 24996
rect 42612 25052 42676 25056
rect 42612 24996 42616 25052
rect 42616 24996 42672 25052
rect 42672 24996 42676 25052
rect 42612 24992 42676 24996
rect 42692 25052 42756 25056
rect 42692 24996 42696 25052
rect 42696 24996 42752 25052
rect 42752 24996 42756 25052
rect 42692 24992 42756 24996
rect 42772 25052 42836 25056
rect 42772 24996 42776 25052
rect 42776 24996 42832 25052
rect 42832 24996 42836 25052
rect 42772 24992 42836 24996
rect 42852 25052 42916 25056
rect 42852 24996 42856 25052
rect 42856 24996 42912 25052
rect 42912 24996 42916 25052
rect 42852 24992 42916 24996
rect 47612 25052 47676 25056
rect 47612 24996 47616 25052
rect 47616 24996 47672 25052
rect 47672 24996 47676 25052
rect 47612 24992 47676 24996
rect 47692 25052 47756 25056
rect 47692 24996 47696 25052
rect 47696 24996 47752 25052
rect 47752 24996 47756 25052
rect 47692 24992 47756 24996
rect 47772 25052 47836 25056
rect 47772 24996 47776 25052
rect 47776 24996 47832 25052
rect 47832 24996 47836 25052
rect 47772 24992 47836 24996
rect 47852 25052 47916 25056
rect 47852 24996 47856 25052
rect 47856 24996 47912 25052
rect 47912 24996 47916 25052
rect 47852 24992 47916 24996
rect 52612 25052 52676 25056
rect 52612 24996 52616 25052
rect 52616 24996 52672 25052
rect 52672 24996 52676 25052
rect 52612 24992 52676 24996
rect 52692 25052 52756 25056
rect 52692 24996 52696 25052
rect 52696 24996 52752 25052
rect 52752 24996 52756 25052
rect 52692 24992 52756 24996
rect 52772 25052 52836 25056
rect 52772 24996 52776 25052
rect 52776 24996 52832 25052
rect 52832 24996 52836 25052
rect 52772 24992 52836 24996
rect 52852 25052 52916 25056
rect 52852 24996 52856 25052
rect 52856 24996 52912 25052
rect 52912 24996 52916 25052
rect 52852 24992 52916 24996
rect 57612 25052 57676 25056
rect 57612 24996 57616 25052
rect 57616 24996 57672 25052
rect 57672 24996 57676 25052
rect 57612 24992 57676 24996
rect 57692 25052 57756 25056
rect 57692 24996 57696 25052
rect 57696 24996 57752 25052
rect 57752 24996 57756 25052
rect 57692 24992 57756 24996
rect 57772 25052 57836 25056
rect 57772 24996 57776 25052
rect 57776 24996 57832 25052
rect 57832 24996 57836 25052
rect 57772 24992 57836 24996
rect 57852 25052 57916 25056
rect 57852 24996 57856 25052
rect 57856 24996 57912 25052
rect 57912 24996 57916 25052
rect 57852 24992 57916 24996
rect 1952 24508 2016 24512
rect 1952 24452 1956 24508
rect 1956 24452 2012 24508
rect 2012 24452 2016 24508
rect 1952 24448 2016 24452
rect 2032 24508 2096 24512
rect 2032 24452 2036 24508
rect 2036 24452 2092 24508
rect 2092 24452 2096 24508
rect 2032 24448 2096 24452
rect 2112 24508 2176 24512
rect 2112 24452 2116 24508
rect 2116 24452 2172 24508
rect 2172 24452 2176 24508
rect 2112 24448 2176 24452
rect 2192 24508 2256 24512
rect 2192 24452 2196 24508
rect 2196 24452 2252 24508
rect 2252 24452 2256 24508
rect 2192 24448 2256 24452
rect 6952 24508 7016 24512
rect 6952 24452 6956 24508
rect 6956 24452 7012 24508
rect 7012 24452 7016 24508
rect 6952 24448 7016 24452
rect 7032 24508 7096 24512
rect 7032 24452 7036 24508
rect 7036 24452 7092 24508
rect 7092 24452 7096 24508
rect 7032 24448 7096 24452
rect 7112 24508 7176 24512
rect 7112 24452 7116 24508
rect 7116 24452 7172 24508
rect 7172 24452 7176 24508
rect 7112 24448 7176 24452
rect 7192 24508 7256 24512
rect 7192 24452 7196 24508
rect 7196 24452 7252 24508
rect 7252 24452 7256 24508
rect 7192 24448 7256 24452
rect 11952 24508 12016 24512
rect 11952 24452 11956 24508
rect 11956 24452 12012 24508
rect 12012 24452 12016 24508
rect 11952 24448 12016 24452
rect 12032 24508 12096 24512
rect 12032 24452 12036 24508
rect 12036 24452 12092 24508
rect 12092 24452 12096 24508
rect 12032 24448 12096 24452
rect 12112 24508 12176 24512
rect 12112 24452 12116 24508
rect 12116 24452 12172 24508
rect 12172 24452 12176 24508
rect 12112 24448 12176 24452
rect 12192 24508 12256 24512
rect 12192 24452 12196 24508
rect 12196 24452 12252 24508
rect 12252 24452 12256 24508
rect 12192 24448 12256 24452
rect 16952 24508 17016 24512
rect 16952 24452 16956 24508
rect 16956 24452 17012 24508
rect 17012 24452 17016 24508
rect 16952 24448 17016 24452
rect 17032 24508 17096 24512
rect 17032 24452 17036 24508
rect 17036 24452 17092 24508
rect 17092 24452 17096 24508
rect 17032 24448 17096 24452
rect 17112 24508 17176 24512
rect 17112 24452 17116 24508
rect 17116 24452 17172 24508
rect 17172 24452 17176 24508
rect 17112 24448 17176 24452
rect 17192 24508 17256 24512
rect 17192 24452 17196 24508
rect 17196 24452 17252 24508
rect 17252 24452 17256 24508
rect 17192 24448 17256 24452
rect 21952 24508 22016 24512
rect 21952 24452 21956 24508
rect 21956 24452 22012 24508
rect 22012 24452 22016 24508
rect 21952 24448 22016 24452
rect 22032 24508 22096 24512
rect 22032 24452 22036 24508
rect 22036 24452 22092 24508
rect 22092 24452 22096 24508
rect 22032 24448 22096 24452
rect 22112 24508 22176 24512
rect 22112 24452 22116 24508
rect 22116 24452 22172 24508
rect 22172 24452 22176 24508
rect 22112 24448 22176 24452
rect 22192 24508 22256 24512
rect 22192 24452 22196 24508
rect 22196 24452 22252 24508
rect 22252 24452 22256 24508
rect 22192 24448 22256 24452
rect 26952 24508 27016 24512
rect 26952 24452 26956 24508
rect 26956 24452 27012 24508
rect 27012 24452 27016 24508
rect 26952 24448 27016 24452
rect 27032 24508 27096 24512
rect 27032 24452 27036 24508
rect 27036 24452 27092 24508
rect 27092 24452 27096 24508
rect 27032 24448 27096 24452
rect 27112 24508 27176 24512
rect 27112 24452 27116 24508
rect 27116 24452 27172 24508
rect 27172 24452 27176 24508
rect 27112 24448 27176 24452
rect 27192 24508 27256 24512
rect 27192 24452 27196 24508
rect 27196 24452 27252 24508
rect 27252 24452 27256 24508
rect 27192 24448 27256 24452
rect 31952 24508 32016 24512
rect 31952 24452 31956 24508
rect 31956 24452 32012 24508
rect 32012 24452 32016 24508
rect 31952 24448 32016 24452
rect 32032 24508 32096 24512
rect 32032 24452 32036 24508
rect 32036 24452 32092 24508
rect 32092 24452 32096 24508
rect 32032 24448 32096 24452
rect 32112 24508 32176 24512
rect 32112 24452 32116 24508
rect 32116 24452 32172 24508
rect 32172 24452 32176 24508
rect 32112 24448 32176 24452
rect 32192 24508 32256 24512
rect 32192 24452 32196 24508
rect 32196 24452 32252 24508
rect 32252 24452 32256 24508
rect 32192 24448 32256 24452
rect 36952 24508 37016 24512
rect 36952 24452 36956 24508
rect 36956 24452 37012 24508
rect 37012 24452 37016 24508
rect 36952 24448 37016 24452
rect 37032 24508 37096 24512
rect 37032 24452 37036 24508
rect 37036 24452 37092 24508
rect 37092 24452 37096 24508
rect 37032 24448 37096 24452
rect 37112 24508 37176 24512
rect 37112 24452 37116 24508
rect 37116 24452 37172 24508
rect 37172 24452 37176 24508
rect 37112 24448 37176 24452
rect 37192 24508 37256 24512
rect 37192 24452 37196 24508
rect 37196 24452 37252 24508
rect 37252 24452 37256 24508
rect 37192 24448 37256 24452
rect 41952 24508 42016 24512
rect 41952 24452 41956 24508
rect 41956 24452 42012 24508
rect 42012 24452 42016 24508
rect 41952 24448 42016 24452
rect 42032 24508 42096 24512
rect 42032 24452 42036 24508
rect 42036 24452 42092 24508
rect 42092 24452 42096 24508
rect 42032 24448 42096 24452
rect 42112 24508 42176 24512
rect 42112 24452 42116 24508
rect 42116 24452 42172 24508
rect 42172 24452 42176 24508
rect 42112 24448 42176 24452
rect 42192 24508 42256 24512
rect 42192 24452 42196 24508
rect 42196 24452 42252 24508
rect 42252 24452 42256 24508
rect 42192 24448 42256 24452
rect 46952 24508 47016 24512
rect 46952 24452 46956 24508
rect 46956 24452 47012 24508
rect 47012 24452 47016 24508
rect 46952 24448 47016 24452
rect 47032 24508 47096 24512
rect 47032 24452 47036 24508
rect 47036 24452 47092 24508
rect 47092 24452 47096 24508
rect 47032 24448 47096 24452
rect 47112 24508 47176 24512
rect 47112 24452 47116 24508
rect 47116 24452 47172 24508
rect 47172 24452 47176 24508
rect 47112 24448 47176 24452
rect 47192 24508 47256 24512
rect 47192 24452 47196 24508
rect 47196 24452 47252 24508
rect 47252 24452 47256 24508
rect 47192 24448 47256 24452
rect 51952 24508 52016 24512
rect 51952 24452 51956 24508
rect 51956 24452 52012 24508
rect 52012 24452 52016 24508
rect 51952 24448 52016 24452
rect 52032 24508 52096 24512
rect 52032 24452 52036 24508
rect 52036 24452 52092 24508
rect 52092 24452 52096 24508
rect 52032 24448 52096 24452
rect 52112 24508 52176 24512
rect 52112 24452 52116 24508
rect 52116 24452 52172 24508
rect 52172 24452 52176 24508
rect 52112 24448 52176 24452
rect 52192 24508 52256 24512
rect 52192 24452 52196 24508
rect 52196 24452 52252 24508
rect 52252 24452 52256 24508
rect 52192 24448 52256 24452
rect 56952 24508 57016 24512
rect 56952 24452 56956 24508
rect 56956 24452 57012 24508
rect 57012 24452 57016 24508
rect 56952 24448 57016 24452
rect 57032 24508 57096 24512
rect 57032 24452 57036 24508
rect 57036 24452 57092 24508
rect 57092 24452 57096 24508
rect 57032 24448 57096 24452
rect 57112 24508 57176 24512
rect 57112 24452 57116 24508
rect 57116 24452 57172 24508
rect 57172 24452 57176 24508
rect 57112 24448 57176 24452
rect 57192 24508 57256 24512
rect 57192 24452 57196 24508
rect 57196 24452 57252 24508
rect 57252 24452 57256 24508
rect 57192 24448 57256 24452
rect 2612 23964 2676 23968
rect 2612 23908 2616 23964
rect 2616 23908 2672 23964
rect 2672 23908 2676 23964
rect 2612 23904 2676 23908
rect 2692 23964 2756 23968
rect 2692 23908 2696 23964
rect 2696 23908 2752 23964
rect 2752 23908 2756 23964
rect 2692 23904 2756 23908
rect 2772 23964 2836 23968
rect 2772 23908 2776 23964
rect 2776 23908 2832 23964
rect 2832 23908 2836 23964
rect 2772 23904 2836 23908
rect 2852 23964 2916 23968
rect 2852 23908 2856 23964
rect 2856 23908 2912 23964
rect 2912 23908 2916 23964
rect 2852 23904 2916 23908
rect 7612 23964 7676 23968
rect 7612 23908 7616 23964
rect 7616 23908 7672 23964
rect 7672 23908 7676 23964
rect 7612 23904 7676 23908
rect 7692 23964 7756 23968
rect 7692 23908 7696 23964
rect 7696 23908 7752 23964
rect 7752 23908 7756 23964
rect 7692 23904 7756 23908
rect 7772 23964 7836 23968
rect 7772 23908 7776 23964
rect 7776 23908 7832 23964
rect 7832 23908 7836 23964
rect 7772 23904 7836 23908
rect 7852 23964 7916 23968
rect 7852 23908 7856 23964
rect 7856 23908 7912 23964
rect 7912 23908 7916 23964
rect 7852 23904 7916 23908
rect 12612 23964 12676 23968
rect 12612 23908 12616 23964
rect 12616 23908 12672 23964
rect 12672 23908 12676 23964
rect 12612 23904 12676 23908
rect 12692 23964 12756 23968
rect 12692 23908 12696 23964
rect 12696 23908 12752 23964
rect 12752 23908 12756 23964
rect 12692 23904 12756 23908
rect 12772 23964 12836 23968
rect 12772 23908 12776 23964
rect 12776 23908 12832 23964
rect 12832 23908 12836 23964
rect 12772 23904 12836 23908
rect 12852 23964 12916 23968
rect 12852 23908 12856 23964
rect 12856 23908 12912 23964
rect 12912 23908 12916 23964
rect 12852 23904 12916 23908
rect 17612 23964 17676 23968
rect 17612 23908 17616 23964
rect 17616 23908 17672 23964
rect 17672 23908 17676 23964
rect 17612 23904 17676 23908
rect 17692 23964 17756 23968
rect 17692 23908 17696 23964
rect 17696 23908 17752 23964
rect 17752 23908 17756 23964
rect 17692 23904 17756 23908
rect 17772 23964 17836 23968
rect 17772 23908 17776 23964
rect 17776 23908 17832 23964
rect 17832 23908 17836 23964
rect 17772 23904 17836 23908
rect 17852 23964 17916 23968
rect 17852 23908 17856 23964
rect 17856 23908 17912 23964
rect 17912 23908 17916 23964
rect 17852 23904 17916 23908
rect 22612 23964 22676 23968
rect 22612 23908 22616 23964
rect 22616 23908 22672 23964
rect 22672 23908 22676 23964
rect 22612 23904 22676 23908
rect 22692 23964 22756 23968
rect 22692 23908 22696 23964
rect 22696 23908 22752 23964
rect 22752 23908 22756 23964
rect 22692 23904 22756 23908
rect 22772 23964 22836 23968
rect 22772 23908 22776 23964
rect 22776 23908 22832 23964
rect 22832 23908 22836 23964
rect 22772 23904 22836 23908
rect 22852 23964 22916 23968
rect 22852 23908 22856 23964
rect 22856 23908 22912 23964
rect 22912 23908 22916 23964
rect 22852 23904 22916 23908
rect 27612 23964 27676 23968
rect 27612 23908 27616 23964
rect 27616 23908 27672 23964
rect 27672 23908 27676 23964
rect 27612 23904 27676 23908
rect 27692 23964 27756 23968
rect 27692 23908 27696 23964
rect 27696 23908 27752 23964
rect 27752 23908 27756 23964
rect 27692 23904 27756 23908
rect 27772 23964 27836 23968
rect 27772 23908 27776 23964
rect 27776 23908 27832 23964
rect 27832 23908 27836 23964
rect 27772 23904 27836 23908
rect 27852 23964 27916 23968
rect 27852 23908 27856 23964
rect 27856 23908 27912 23964
rect 27912 23908 27916 23964
rect 27852 23904 27916 23908
rect 32612 23964 32676 23968
rect 32612 23908 32616 23964
rect 32616 23908 32672 23964
rect 32672 23908 32676 23964
rect 32612 23904 32676 23908
rect 32692 23964 32756 23968
rect 32692 23908 32696 23964
rect 32696 23908 32752 23964
rect 32752 23908 32756 23964
rect 32692 23904 32756 23908
rect 32772 23964 32836 23968
rect 32772 23908 32776 23964
rect 32776 23908 32832 23964
rect 32832 23908 32836 23964
rect 32772 23904 32836 23908
rect 32852 23964 32916 23968
rect 32852 23908 32856 23964
rect 32856 23908 32912 23964
rect 32912 23908 32916 23964
rect 32852 23904 32916 23908
rect 37612 23964 37676 23968
rect 37612 23908 37616 23964
rect 37616 23908 37672 23964
rect 37672 23908 37676 23964
rect 37612 23904 37676 23908
rect 37692 23964 37756 23968
rect 37692 23908 37696 23964
rect 37696 23908 37752 23964
rect 37752 23908 37756 23964
rect 37692 23904 37756 23908
rect 37772 23964 37836 23968
rect 37772 23908 37776 23964
rect 37776 23908 37832 23964
rect 37832 23908 37836 23964
rect 37772 23904 37836 23908
rect 37852 23964 37916 23968
rect 37852 23908 37856 23964
rect 37856 23908 37912 23964
rect 37912 23908 37916 23964
rect 37852 23904 37916 23908
rect 42612 23964 42676 23968
rect 42612 23908 42616 23964
rect 42616 23908 42672 23964
rect 42672 23908 42676 23964
rect 42612 23904 42676 23908
rect 42692 23964 42756 23968
rect 42692 23908 42696 23964
rect 42696 23908 42752 23964
rect 42752 23908 42756 23964
rect 42692 23904 42756 23908
rect 42772 23964 42836 23968
rect 42772 23908 42776 23964
rect 42776 23908 42832 23964
rect 42832 23908 42836 23964
rect 42772 23904 42836 23908
rect 42852 23964 42916 23968
rect 42852 23908 42856 23964
rect 42856 23908 42912 23964
rect 42912 23908 42916 23964
rect 42852 23904 42916 23908
rect 47612 23964 47676 23968
rect 47612 23908 47616 23964
rect 47616 23908 47672 23964
rect 47672 23908 47676 23964
rect 47612 23904 47676 23908
rect 47692 23964 47756 23968
rect 47692 23908 47696 23964
rect 47696 23908 47752 23964
rect 47752 23908 47756 23964
rect 47692 23904 47756 23908
rect 47772 23964 47836 23968
rect 47772 23908 47776 23964
rect 47776 23908 47832 23964
rect 47832 23908 47836 23964
rect 47772 23904 47836 23908
rect 47852 23964 47916 23968
rect 47852 23908 47856 23964
rect 47856 23908 47912 23964
rect 47912 23908 47916 23964
rect 47852 23904 47916 23908
rect 52612 23964 52676 23968
rect 52612 23908 52616 23964
rect 52616 23908 52672 23964
rect 52672 23908 52676 23964
rect 52612 23904 52676 23908
rect 52692 23964 52756 23968
rect 52692 23908 52696 23964
rect 52696 23908 52752 23964
rect 52752 23908 52756 23964
rect 52692 23904 52756 23908
rect 52772 23964 52836 23968
rect 52772 23908 52776 23964
rect 52776 23908 52832 23964
rect 52832 23908 52836 23964
rect 52772 23904 52836 23908
rect 52852 23964 52916 23968
rect 52852 23908 52856 23964
rect 52856 23908 52912 23964
rect 52912 23908 52916 23964
rect 52852 23904 52916 23908
rect 57612 23964 57676 23968
rect 57612 23908 57616 23964
rect 57616 23908 57672 23964
rect 57672 23908 57676 23964
rect 57612 23904 57676 23908
rect 57692 23964 57756 23968
rect 57692 23908 57696 23964
rect 57696 23908 57752 23964
rect 57752 23908 57756 23964
rect 57692 23904 57756 23908
rect 57772 23964 57836 23968
rect 57772 23908 57776 23964
rect 57776 23908 57832 23964
rect 57832 23908 57836 23964
rect 57772 23904 57836 23908
rect 57852 23964 57916 23968
rect 57852 23908 57856 23964
rect 57856 23908 57912 23964
rect 57912 23908 57916 23964
rect 57852 23904 57916 23908
rect 1952 23420 2016 23424
rect 1952 23364 1956 23420
rect 1956 23364 2012 23420
rect 2012 23364 2016 23420
rect 1952 23360 2016 23364
rect 2032 23420 2096 23424
rect 2032 23364 2036 23420
rect 2036 23364 2092 23420
rect 2092 23364 2096 23420
rect 2032 23360 2096 23364
rect 2112 23420 2176 23424
rect 2112 23364 2116 23420
rect 2116 23364 2172 23420
rect 2172 23364 2176 23420
rect 2112 23360 2176 23364
rect 2192 23420 2256 23424
rect 2192 23364 2196 23420
rect 2196 23364 2252 23420
rect 2252 23364 2256 23420
rect 2192 23360 2256 23364
rect 6952 23420 7016 23424
rect 6952 23364 6956 23420
rect 6956 23364 7012 23420
rect 7012 23364 7016 23420
rect 6952 23360 7016 23364
rect 7032 23420 7096 23424
rect 7032 23364 7036 23420
rect 7036 23364 7092 23420
rect 7092 23364 7096 23420
rect 7032 23360 7096 23364
rect 7112 23420 7176 23424
rect 7112 23364 7116 23420
rect 7116 23364 7172 23420
rect 7172 23364 7176 23420
rect 7112 23360 7176 23364
rect 7192 23420 7256 23424
rect 7192 23364 7196 23420
rect 7196 23364 7252 23420
rect 7252 23364 7256 23420
rect 7192 23360 7256 23364
rect 11952 23420 12016 23424
rect 11952 23364 11956 23420
rect 11956 23364 12012 23420
rect 12012 23364 12016 23420
rect 11952 23360 12016 23364
rect 12032 23420 12096 23424
rect 12032 23364 12036 23420
rect 12036 23364 12092 23420
rect 12092 23364 12096 23420
rect 12032 23360 12096 23364
rect 12112 23420 12176 23424
rect 12112 23364 12116 23420
rect 12116 23364 12172 23420
rect 12172 23364 12176 23420
rect 12112 23360 12176 23364
rect 12192 23420 12256 23424
rect 12192 23364 12196 23420
rect 12196 23364 12252 23420
rect 12252 23364 12256 23420
rect 12192 23360 12256 23364
rect 16952 23420 17016 23424
rect 16952 23364 16956 23420
rect 16956 23364 17012 23420
rect 17012 23364 17016 23420
rect 16952 23360 17016 23364
rect 17032 23420 17096 23424
rect 17032 23364 17036 23420
rect 17036 23364 17092 23420
rect 17092 23364 17096 23420
rect 17032 23360 17096 23364
rect 17112 23420 17176 23424
rect 17112 23364 17116 23420
rect 17116 23364 17172 23420
rect 17172 23364 17176 23420
rect 17112 23360 17176 23364
rect 17192 23420 17256 23424
rect 17192 23364 17196 23420
rect 17196 23364 17252 23420
rect 17252 23364 17256 23420
rect 17192 23360 17256 23364
rect 21952 23420 22016 23424
rect 21952 23364 21956 23420
rect 21956 23364 22012 23420
rect 22012 23364 22016 23420
rect 21952 23360 22016 23364
rect 22032 23420 22096 23424
rect 22032 23364 22036 23420
rect 22036 23364 22092 23420
rect 22092 23364 22096 23420
rect 22032 23360 22096 23364
rect 22112 23420 22176 23424
rect 22112 23364 22116 23420
rect 22116 23364 22172 23420
rect 22172 23364 22176 23420
rect 22112 23360 22176 23364
rect 22192 23420 22256 23424
rect 22192 23364 22196 23420
rect 22196 23364 22252 23420
rect 22252 23364 22256 23420
rect 22192 23360 22256 23364
rect 26952 23420 27016 23424
rect 26952 23364 26956 23420
rect 26956 23364 27012 23420
rect 27012 23364 27016 23420
rect 26952 23360 27016 23364
rect 27032 23420 27096 23424
rect 27032 23364 27036 23420
rect 27036 23364 27092 23420
rect 27092 23364 27096 23420
rect 27032 23360 27096 23364
rect 27112 23420 27176 23424
rect 27112 23364 27116 23420
rect 27116 23364 27172 23420
rect 27172 23364 27176 23420
rect 27112 23360 27176 23364
rect 27192 23420 27256 23424
rect 27192 23364 27196 23420
rect 27196 23364 27252 23420
rect 27252 23364 27256 23420
rect 27192 23360 27256 23364
rect 31952 23420 32016 23424
rect 31952 23364 31956 23420
rect 31956 23364 32012 23420
rect 32012 23364 32016 23420
rect 31952 23360 32016 23364
rect 32032 23420 32096 23424
rect 32032 23364 32036 23420
rect 32036 23364 32092 23420
rect 32092 23364 32096 23420
rect 32032 23360 32096 23364
rect 32112 23420 32176 23424
rect 32112 23364 32116 23420
rect 32116 23364 32172 23420
rect 32172 23364 32176 23420
rect 32112 23360 32176 23364
rect 32192 23420 32256 23424
rect 32192 23364 32196 23420
rect 32196 23364 32252 23420
rect 32252 23364 32256 23420
rect 32192 23360 32256 23364
rect 36952 23420 37016 23424
rect 36952 23364 36956 23420
rect 36956 23364 37012 23420
rect 37012 23364 37016 23420
rect 36952 23360 37016 23364
rect 37032 23420 37096 23424
rect 37032 23364 37036 23420
rect 37036 23364 37092 23420
rect 37092 23364 37096 23420
rect 37032 23360 37096 23364
rect 37112 23420 37176 23424
rect 37112 23364 37116 23420
rect 37116 23364 37172 23420
rect 37172 23364 37176 23420
rect 37112 23360 37176 23364
rect 37192 23420 37256 23424
rect 37192 23364 37196 23420
rect 37196 23364 37252 23420
rect 37252 23364 37256 23420
rect 37192 23360 37256 23364
rect 41952 23420 42016 23424
rect 41952 23364 41956 23420
rect 41956 23364 42012 23420
rect 42012 23364 42016 23420
rect 41952 23360 42016 23364
rect 42032 23420 42096 23424
rect 42032 23364 42036 23420
rect 42036 23364 42092 23420
rect 42092 23364 42096 23420
rect 42032 23360 42096 23364
rect 42112 23420 42176 23424
rect 42112 23364 42116 23420
rect 42116 23364 42172 23420
rect 42172 23364 42176 23420
rect 42112 23360 42176 23364
rect 42192 23420 42256 23424
rect 42192 23364 42196 23420
rect 42196 23364 42252 23420
rect 42252 23364 42256 23420
rect 42192 23360 42256 23364
rect 46952 23420 47016 23424
rect 46952 23364 46956 23420
rect 46956 23364 47012 23420
rect 47012 23364 47016 23420
rect 46952 23360 47016 23364
rect 47032 23420 47096 23424
rect 47032 23364 47036 23420
rect 47036 23364 47092 23420
rect 47092 23364 47096 23420
rect 47032 23360 47096 23364
rect 47112 23420 47176 23424
rect 47112 23364 47116 23420
rect 47116 23364 47172 23420
rect 47172 23364 47176 23420
rect 47112 23360 47176 23364
rect 47192 23420 47256 23424
rect 47192 23364 47196 23420
rect 47196 23364 47252 23420
rect 47252 23364 47256 23420
rect 47192 23360 47256 23364
rect 51952 23420 52016 23424
rect 51952 23364 51956 23420
rect 51956 23364 52012 23420
rect 52012 23364 52016 23420
rect 51952 23360 52016 23364
rect 52032 23420 52096 23424
rect 52032 23364 52036 23420
rect 52036 23364 52092 23420
rect 52092 23364 52096 23420
rect 52032 23360 52096 23364
rect 52112 23420 52176 23424
rect 52112 23364 52116 23420
rect 52116 23364 52172 23420
rect 52172 23364 52176 23420
rect 52112 23360 52176 23364
rect 52192 23420 52256 23424
rect 52192 23364 52196 23420
rect 52196 23364 52252 23420
rect 52252 23364 52256 23420
rect 52192 23360 52256 23364
rect 56952 23420 57016 23424
rect 56952 23364 56956 23420
rect 56956 23364 57012 23420
rect 57012 23364 57016 23420
rect 56952 23360 57016 23364
rect 57032 23420 57096 23424
rect 57032 23364 57036 23420
rect 57036 23364 57092 23420
rect 57092 23364 57096 23420
rect 57032 23360 57096 23364
rect 57112 23420 57176 23424
rect 57112 23364 57116 23420
rect 57116 23364 57172 23420
rect 57172 23364 57176 23420
rect 57112 23360 57176 23364
rect 57192 23420 57256 23424
rect 57192 23364 57196 23420
rect 57196 23364 57252 23420
rect 57252 23364 57256 23420
rect 57192 23360 57256 23364
rect 2612 22876 2676 22880
rect 2612 22820 2616 22876
rect 2616 22820 2672 22876
rect 2672 22820 2676 22876
rect 2612 22816 2676 22820
rect 2692 22876 2756 22880
rect 2692 22820 2696 22876
rect 2696 22820 2752 22876
rect 2752 22820 2756 22876
rect 2692 22816 2756 22820
rect 2772 22876 2836 22880
rect 2772 22820 2776 22876
rect 2776 22820 2832 22876
rect 2832 22820 2836 22876
rect 2772 22816 2836 22820
rect 2852 22876 2916 22880
rect 2852 22820 2856 22876
rect 2856 22820 2912 22876
rect 2912 22820 2916 22876
rect 2852 22816 2916 22820
rect 7612 22876 7676 22880
rect 7612 22820 7616 22876
rect 7616 22820 7672 22876
rect 7672 22820 7676 22876
rect 7612 22816 7676 22820
rect 7692 22876 7756 22880
rect 7692 22820 7696 22876
rect 7696 22820 7752 22876
rect 7752 22820 7756 22876
rect 7692 22816 7756 22820
rect 7772 22876 7836 22880
rect 7772 22820 7776 22876
rect 7776 22820 7832 22876
rect 7832 22820 7836 22876
rect 7772 22816 7836 22820
rect 7852 22876 7916 22880
rect 7852 22820 7856 22876
rect 7856 22820 7912 22876
rect 7912 22820 7916 22876
rect 7852 22816 7916 22820
rect 12612 22876 12676 22880
rect 12612 22820 12616 22876
rect 12616 22820 12672 22876
rect 12672 22820 12676 22876
rect 12612 22816 12676 22820
rect 12692 22876 12756 22880
rect 12692 22820 12696 22876
rect 12696 22820 12752 22876
rect 12752 22820 12756 22876
rect 12692 22816 12756 22820
rect 12772 22876 12836 22880
rect 12772 22820 12776 22876
rect 12776 22820 12832 22876
rect 12832 22820 12836 22876
rect 12772 22816 12836 22820
rect 12852 22876 12916 22880
rect 12852 22820 12856 22876
rect 12856 22820 12912 22876
rect 12912 22820 12916 22876
rect 12852 22816 12916 22820
rect 17612 22876 17676 22880
rect 17612 22820 17616 22876
rect 17616 22820 17672 22876
rect 17672 22820 17676 22876
rect 17612 22816 17676 22820
rect 17692 22876 17756 22880
rect 17692 22820 17696 22876
rect 17696 22820 17752 22876
rect 17752 22820 17756 22876
rect 17692 22816 17756 22820
rect 17772 22876 17836 22880
rect 17772 22820 17776 22876
rect 17776 22820 17832 22876
rect 17832 22820 17836 22876
rect 17772 22816 17836 22820
rect 17852 22876 17916 22880
rect 17852 22820 17856 22876
rect 17856 22820 17912 22876
rect 17912 22820 17916 22876
rect 17852 22816 17916 22820
rect 22612 22876 22676 22880
rect 22612 22820 22616 22876
rect 22616 22820 22672 22876
rect 22672 22820 22676 22876
rect 22612 22816 22676 22820
rect 22692 22876 22756 22880
rect 22692 22820 22696 22876
rect 22696 22820 22752 22876
rect 22752 22820 22756 22876
rect 22692 22816 22756 22820
rect 22772 22876 22836 22880
rect 22772 22820 22776 22876
rect 22776 22820 22832 22876
rect 22832 22820 22836 22876
rect 22772 22816 22836 22820
rect 22852 22876 22916 22880
rect 22852 22820 22856 22876
rect 22856 22820 22912 22876
rect 22912 22820 22916 22876
rect 22852 22816 22916 22820
rect 27612 22876 27676 22880
rect 27612 22820 27616 22876
rect 27616 22820 27672 22876
rect 27672 22820 27676 22876
rect 27612 22816 27676 22820
rect 27692 22876 27756 22880
rect 27692 22820 27696 22876
rect 27696 22820 27752 22876
rect 27752 22820 27756 22876
rect 27692 22816 27756 22820
rect 27772 22876 27836 22880
rect 27772 22820 27776 22876
rect 27776 22820 27832 22876
rect 27832 22820 27836 22876
rect 27772 22816 27836 22820
rect 27852 22876 27916 22880
rect 27852 22820 27856 22876
rect 27856 22820 27912 22876
rect 27912 22820 27916 22876
rect 27852 22816 27916 22820
rect 32612 22876 32676 22880
rect 32612 22820 32616 22876
rect 32616 22820 32672 22876
rect 32672 22820 32676 22876
rect 32612 22816 32676 22820
rect 32692 22876 32756 22880
rect 32692 22820 32696 22876
rect 32696 22820 32752 22876
rect 32752 22820 32756 22876
rect 32692 22816 32756 22820
rect 32772 22876 32836 22880
rect 32772 22820 32776 22876
rect 32776 22820 32832 22876
rect 32832 22820 32836 22876
rect 32772 22816 32836 22820
rect 32852 22876 32916 22880
rect 32852 22820 32856 22876
rect 32856 22820 32912 22876
rect 32912 22820 32916 22876
rect 32852 22816 32916 22820
rect 37612 22876 37676 22880
rect 37612 22820 37616 22876
rect 37616 22820 37672 22876
rect 37672 22820 37676 22876
rect 37612 22816 37676 22820
rect 37692 22876 37756 22880
rect 37692 22820 37696 22876
rect 37696 22820 37752 22876
rect 37752 22820 37756 22876
rect 37692 22816 37756 22820
rect 37772 22876 37836 22880
rect 37772 22820 37776 22876
rect 37776 22820 37832 22876
rect 37832 22820 37836 22876
rect 37772 22816 37836 22820
rect 37852 22876 37916 22880
rect 37852 22820 37856 22876
rect 37856 22820 37912 22876
rect 37912 22820 37916 22876
rect 37852 22816 37916 22820
rect 42612 22876 42676 22880
rect 42612 22820 42616 22876
rect 42616 22820 42672 22876
rect 42672 22820 42676 22876
rect 42612 22816 42676 22820
rect 42692 22876 42756 22880
rect 42692 22820 42696 22876
rect 42696 22820 42752 22876
rect 42752 22820 42756 22876
rect 42692 22816 42756 22820
rect 42772 22876 42836 22880
rect 42772 22820 42776 22876
rect 42776 22820 42832 22876
rect 42832 22820 42836 22876
rect 42772 22816 42836 22820
rect 42852 22876 42916 22880
rect 42852 22820 42856 22876
rect 42856 22820 42912 22876
rect 42912 22820 42916 22876
rect 42852 22816 42916 22820
rect 47612 22876 47676 22880
rect 47612 22820 47616 22876
rect 47616 22820 47672 22876
rect 47672 22820 47676 22876
rect 47612 22816 47676 22820
rect 47692 22876 47756 22880
rect 47692 22820 47696 22876
rect 47696 22820 47752 22876
rect 47752 22820 47756 22876
rect 47692 22816 47756 22820
rect 47772 22876 47836 22880
rect 47772 22820 47776 22876
rect 47776 22820 47832 22876
rect 47832 22820 47836 22876
rect 47772 22816 47836 22820
rect 47852 22876 47916 22880
rect 47852 22820 47856 22876
rect 47856 22820 47912 22876
rect 47912 22820 47916 22876
rect 47852 22816 47916 22820
rect 52612 22876 52676 22880
rect 52612 22820 52616 22876
rect 52616 22820 52672 22876
rect 52672 22820 52676 22876
rect 52612 22816 52676 22820
rect 52692 22876 52756 22880
rect 52692 22820 52696 22876
rect 52696 22820 52752 22876
rect 52752 22820 52756 22876
rect 52692 22816 52756 22820
rect 52772 22876 52836 22880
rect 52772 22820 52776 22876
rect 52776 22820 52832 22876
rect 52832 22820 52836 22876
rect 52772 22816 52836 22820
rect 52852 22876 52916 22880
rect 52852 22820 52856 22876
rect 52856 22820 52912 22876
rect 52912 22820 52916 22876
rect 52852 22816 52916 22820
rect 57612 22876 57676 22880
rect 57612 22820 57616 22876
rect 57616 22820 57672 22876
rect 57672 22820 57676 22876
rect 57612 22816 57676 22820
rect 57692 22876 57756 22880
rect 57692 22820 57696 22876
rect 57696 22820 57752 22876
rect 57752 22820 57756 22876
rect 57692 22816 57756 22820
rect 57772 22876 57836 22880
rect 57772 22820 57776 22876
rect 57776 22820 57832 22876
rect 57832 22820 57836 22876
rect 57772 22816 57836 22820
rect 57852 22876 57916 22880
rect 57852 22820 57856 22876
rect 57856 22820 57912 22876
rect 57912 22820 57916 22876
rect 57852 22816 57916 22820
rect 1952 22332 2016 22336
rect 1952 22276 1956 22332
rect 1956 22276 2012 22332
rect 2012 22276 2016 22332
rect 1952 22272 2016 22276
rect 2032 22332 2096 22336
rect 2032 22276 2036 22332
rect 2036 22276 2092 22332
rect 2092 22276 2096 22332
rect 2032 22272 2096 22276
rect 2112 22332 2176 22336
rect 2112 22276 2116 22332
rect 2116 22276 2172 22332
rect 2172 22276 2176 22332
rect 2112 22272 2176 22276
rect 2192 22332 2256 22336
rect 2192 22276 2196 22332
rect 2196 22276 2252 22332
rect 2252 22276 2256 22332
rect 2192 22272 2256 22276
rect 6952 22332 7016 22336
rect 6952 22276 6956 22332
rect 6956 22276 7012 22332
rect 7012 22276 7016 22332
rect 6952 22272 7016 22276
rect 7032 22332 7096 22336
rect 7032 22276 7036 22332
rect 7036 22276 7092 22332
rect 7092 22276 7096 22332
rect 7032 22272 7096 22276
rect 7112 22332 7176 22336
rect 7112 22276 7116 22332
rect 7116 22276 7172 22332
rect 7172 22276 7176 22332
rect 7112 22272 7176 22276
rect 7192 22332 7256 22336
rect 7192 22276 7196 22332
rect 7196 22276 7252 22332
rect 7252 22276 7256 22332
rect 7192 22272 7256 22276
rect 11952 22332 12016 22336
rect 11952 22276 11956 22332
rect 11956 22276 12012 22332
rect 12012 22276 12016 22332
rect 11952 22272 12016 22276
rect 12032 22332 12096 22336
rect 12032 22276 12036 22332
rect 12036 22276 12092 22332
rect 12092 22276 12096 22332
rect 12032 22272 12096 22276
rect 12112 22332 12176 22336
rect 12112 22276 12116 22332
rect 12116 22276 12172 22332
rect 12172 22276 12176 22332
rect 12112 22272 12176 22276
rect 12192 22332 12256 22336
rect 12192 22276 12196 22332
rect 12196 22276 12252 22332
rect 12252 22276 12256 22332
rect 12192 22272 12256 22276
rect 16952 22332 17016 22336
rect 16952 22276 16956 22332
rect 16956 22276 17012 22332
rect 17012 22276 17016 22332
rect 16952 22272 17016 22276
rect 17032 22332 17096 22336
rect 17032 22276 17036 22332
rect 17036 22276 17092 22332
rect 17092 22276 17096 22332
rect 17032 22272 17096 22276
rect 17112 22332 17176 22336
rect 17112 22276 17116 22332
rect 17116 22276 17172 22332
rect 17172 22276 17176 22332
rect 17112 22272 17176 22276
rect 17192 22332 17256 22336
rect 17192 22276 17196 22332
rect 17196 22276 17252 22332
rect 17252 22276 17256 22332
rect 17192 22272 17256 22276
rect 21952 22332 22016 22336
rect 21952 22276 21956 22332
rect 21956 22276 22012 22332
rect 22012 22276 22016 22332
rect 21952 22272 22016 22276
rect 22032 22332 22096 22336
rect 22032 22276 22036 22332
rect 22036 22276 22092 22332
rect 22092 22276 22096 22332
rect 22032 22272 22096 22276
rect 22112 22332 22176 22336
rect 22112 22276 22116 22332
rect 22116 22276 22172 22332
rect 22172 22276 22176 22332
rect 22112 22272 22176 22276
rect 22192 22332 22256 22336
rect 22192 22276 22196 22332
rect 22196 22276 22252 22332
rect 22252 22276 22256 22332
rect 22192 22272 22256 22276
rect 26952 22332 27016 22336
rect 26952 22276 26956 22332
rect 26956 22276 27012 22332
rect 27012 22276 27016 22332
rect 26952 22272 27016 22276
rect 27032 22332 27096 22336
rect 27032 22276 27036 22332
rect 27036 22276 27092 22332
rect 27092 22276 27096 22332
rect 27032 22272 27096 22276
rect 27112 22332 27176 22336
rect 27112 22276 27116 22332
rect 27116 22276 27172 22332
rect 27172 22276 27176 22332
rect 27112 22272 27176 22276
rect 27192 22332 27256 22336
rect 27192 22276 27196 22332
rect 27196 22276 27252 22332
rect 27252 22276 27256 22332
rect 27192 22272 27256 22276
rect 31952 22332 32016 22336
rect 31952 22276 31956 22332
rect 31956 22276 32012 22332
rect 32012 22276 32016 22332
rect 31952 22272 32016 22276
rect 32032 22332 32096 22336
rect 32032 22276 32036 22332
rect 32036 22276 32092 22332
rect 32092 22276 32096 22332
rect 32032 22272 32096 22276
rect 32112 22332 32176 22336
rect 32112 22276 32116 22332
rect 32116 22276 32172 22332
rect 32172 22276 32176 22332
rect 32112 22272 32176 22276
rect 32192 22332 32256 22336
rect 32192 22276 32196 22332
rect 32196 22276 32252 22332
rect 32252 22276 32256 22332
rect 32192 22272 32256 22276
rect 36952 22332 37016 22336
rect 36952 22276 36956 22332
rect 36956 22276 37012 22332
rect 37012 22276 37016 22332
rect 36952 22272 37016 22276
rect 37032 22332 37096 22336
rect 37032 22276 37036 22332
rect 37036 22276 37092 22332
rect 37092 22276 37096 22332
rect 37032 22272 37096 22276
rect 37112 22332 37176 22336
rect 37112 22276 37116 22332
rect 37116 22276 37172 22332
rect 37172 22276 37176 22332
rect 37112 22272 37176 22276
rect 37192 22332 37256 22336
rect 37192 22276 37196 22332
rect 37196 22276 37252 22332
rect 37252 22276 37256 22332
rect 37192 22272 37256 22276
rect 41952 22332 42016 22336
rect 41952 22276 41956 22332
rect 41956 22276 42012 22332
rect 42012 22276 42016 22332
rect 41952 22272 42016 22276
rect 42032 22332 42096 22336
rect 42032 22276 42036 22332
rect 42036 22276 42092 22332
rect 42092 22276 42096 22332
rect 42032 22272 42096 22276
rect 42112 22332 42176 22336
rect 42112 22276 42116 22332
rect 42116 22276 42172 22332
rect 42172 22276 42176 22332
rect 42112 22272 42176 22276
rect 42192 22332 42256 22336
rect 42192 22276 42196 22332
rect 42196 22276 42252 22332
rect 42252 22276 42256 22332
rect 42192 22272 42256 22276
rect 46952 22332 47016 22336
rect 46952 22276 46956 22332
rect 46956 22276 47012 22332
rect 47012 22276 47016 22332
rect 46952 22272 47016 22276
rect 47032 22332 47096 22336
rect 47032 22276 47036 22332
rect 47036 22276 47092 22332
rect 47092 22276 47096 22332
rect 47032 22272 47096 22276
rect 47112 22332 47176 22336
rect 47112 22276 47116 22332
rect 47116 22276 47172 22332
rect 47172 22276 47176 22332
rect 47112 22272 47176 22276
rect 47192 22332 47256 22336
rect 47192 22276 47196 22332
rect 47196 22276 47252 22332
rect 47252 22276 47256 22332
rect 47192 22272 47256 22276
rect 51952 22332 52016 22336
rect 51952 22276 51956 22332
rect 51956 22276 52012 22332
rect 52012 22276 52016 22332
rect 51952 22272 52016 22276
rect 52032 22332 52096 22336
rect 52032 22276 52036 22332
rect 52036 22276 52092 22332
rect 52092 22276 52096 22332
rect 52032 22272 52096 22276
rect 52112 22332 52176 22336
rect 52112 22276 52116 22332
rect 52116 22276 52172 22332
rect 52172 22276 52176 22332
rect 52112 22272 52176 22276
rect 52192 22332 52256 22336
rect 52192 22276 52196 22332
rect 52196 22276 52252 22332
rect 52252 22276 52256 22332
rect 52192 22272 52256 22276
rect 56952 22332 57016 22336
rect 56952 22276 56956 22332
rect 56956 22276 57012 22332
rect 57012 22276 57016 22332
rect 56952 22272 57016 22276
rect 57032 22332 57096 22336
rect 57032 22276 57036 22332
rect 57036 22276 57092 22332
rect 57092 22276 57096 22332
rect 57032 22272 57096 22276
rect 57112 22332 57176 22336
rect 57112 22276 57116 22332
rect 57116 22276 57172 22332
rect 57172 22276 57176 22332
rect 57112 22272 57176 22276
rect 57192 22332 57256 22336
rect 57192 22276 57196 22332
rect 57196 22276 57252 22332
rect 57252 22276 57256 22332
rect 57192 22272 57256 22276
rect 2612 21788 2676 21792
rect 2612 21732 2616 21788
rect 2616 21732 2672 21788
rect 2672 21732 2676 21788
rect 2612 21728 2676 21732
rect 2692 21788 2756 21792
rect 2692 21732 2696 21788
rect 2696 21732 2752 21788
rect 2752 21732 2756 21788
rect 2692 21728 2756 21732
rect 2772 21788 2836 21792
rect 2772 21732 2776 21788
rect 2776 21732 2832 21788
rect 2832 21732 2836 21788
rect 2772 21728 2836 21732
rect 2852 21788 2916 21792
rect 2852 21732 2856 21788
rect 2856 21732 2912 21788
rect 2912 21732 2916 21788
rect 2852 21728 2916 21732
rect 7612 21788 7676 21792
rect 7612 21732 7616 21788
rect 7616 21732 7672 21788
rect 7672 21732 7676 21788
rect 7612 21728 7676 21732
rect 7692 21788 7756 21792
rect 7692 21732 7696 21788
rect 7696 21732 7752 21788
rect 7752 21732 7756 21788
rect 7692 21728 7756 21732
rect 7772 21788 7836 21792
rect 7772 21732 7776 21788
rect 7776 21732 7832 21788
rect 7832 21732 7836 21788
rect 7772 21728 7836 21732
rect 7852 21788 7916 21792
rect 7852 21732 7856 21788
rect 7856 21732 7912 21788
rect 7912 21732 7916 21788
rect 7852 21728 7916 21732
rect 12612 21788 12676 21792
rect 12612 21732 12616 21788
rect 12616 21732 12672 21788
rect 12672 21732 12676 21788
rect 12612 21728 12676 21732
rect 12692 21788 12756 21792
rect 12692 21732 12696 21788
rect 12696 21732 12752 21788
rect 12752 21732 12756 21788
rect 12692 21728 12756 21732
rect 12772 21788 12836 21792
rect 12772 21732 12776 21788
rect 12776 21732 12832 21788
rect 12832 21732 12836 21788
rect 12772 21728 12836 21732
rect 12852 21788 12916 21792
rect 12852 21732 12856 21788
rect 12856 21732 12912 21788
rect 12912 21732 12916 21788
rect 12852 21728 12916 21732
rect 17612 21788 17676 21792
rect 17612 21732 17616 21788
rect 17616 21732 17672 21788
rect 17672 21732 17676 21788
rect 17612 21728 17676 21732
rect 17692 21788 17756 21792
rect 17692 21732 17696 21788
rect 17696 21732 17752 21788
rect 17752 21732 17756 21788
rect 17692 21728 17756 21732
rect 17772 21788 17836 21792
rect 17772 21732 17776 21788
rect 17776 21732 17832 21788
rect 17832 21732 17836 21788
rect 17772 21728 17836 21732
rect 17852 21788 17916 21792
rect 17852 21732 17856 21788
rect 17856 21732 17912 21788
rect 17912 21732 17916 21788
rect 17852 21728 17916 21732
rect 22612 21788 22676 21792
rect 22612 21732 22616 21788
rect 22616 21732 22672 21788
rect 22672 21732 22676 21788
rect 22612 21728 22676 21732
rect 22692 21788 22756 21792
rect 22692 21732 22696 21788
rect 22696 21732 22752 21788
rect 22752 21732 22756 21788
rect 22692 21728 22756 21732
rect 22772 21788 22836 21792
rect 22772 21732 22776 21788
rect 22776 21732 22832 21788
rect 22832 21732 22836 21788
rect 22772 21728 22836 21732
rect 22852 21788 22916 21792
rect 22852 21732 22856 21788
rect 22856 21732 22912 21788
rect 22912 21732 22916 21788
rect 22852 21728 22916 21732
rect 27612 21788 27676 21792
rect 27612 21732 27616 21788
rect 27616 21732 27672 21788
rect 27672 21732 27676 21788
rect 27612 21728 27676 21732
rect 27692 21788 27756 21792
rect 27692 21732 27696 21788
rect 27696 21732 27752 21788
rect 27752 21732 27756 21788
rect 27692 21728 27756 21732
rect 27772 21788 27836 21792
rect 27772 21732 27776 21788
rect 27776 21732 27832 21788
rect 27832 21732 27836 21788
rect 27772 21728 27836 21732
rect 27852 21788 27916 21792
rect 27852 21732 27856 21788
rect 27856 21732 27912 21788
rect 27912 21732 27916 21788
rect 27852 21728 27916 21732
rect 32612 21788 32676 21792
rect 32612 21732 32616 21788
rect 32616 21732 32672 21788
rect 32672 21732 32676 21788
rect 32612 21728 32676 21732
rect 32692 21788 32756 21792
rect 32692 21732 32696 21788
rect 32696 21732 32752 21788
rect 32752 21732 32756 21788
rect 32692 21728 32756 21732
rect 32772 21788 32836 21792
rect 32772 21732 32776 21788
rect 32776 21732 32832 21788
rect 32832 21732 32836 21788
rect 32772 21728 32836 21732
rect 32852 21788 32916 21792
rect 32852 21732 32856 21788
rect 32856 21732 32912 21788
rect 32912 21732 32916 21788
rect 32852 21728 32916 21732
rect 37612 21788 37676 21792
rect 37612 21732 37616 21788
rect 37616 21732 37672 21788
rect 37672 21732 37676 21788
rect 37612 21728 37676 21732
rect 37692 21788 37756 21792
rect 37692 21732 37696 21788
rect 37696 21732 37752 21788
rect 37752 21732 37756 21788
rect 37692 21728 37756 21732
rect 37772 21788 37836 21792
rect 37772 21732 37776 21788
rect 37776 21732 37832 21788
rect 37832 21732 37836 21788
rect 37772 21728 37836 21732
rect 37852 21788 37916 21792
rect 37852 21732 37856 21788
rect 37856 21732 37912 21788
rect 37912 21732 37916 21788
rect 37852 21728 37916 21732
rect 42612 21788 42676 21792
rect 42612 21732 42616 21788
rect 42616 21732 42672 21788
rect 42672 21732 42676 21788
rect 42612 21728 42676 21732
rect 42692 21788 42756 21792
rect 42692 21732 42696 21788
rect 42696 21732 42752 21788
rect 42752 21732 42756 21788
rect 42692 21728 42756 21732
rect 42772 21788 42836 21792
rect 42772 21732 42776 21788
rect 42776 21732 42832 21788
rect 42832 21732 42836 21788
rect 42772 21728 42836 21732
rect 42852 21788 42916 21792
rect 42852 21732 42856 21788
rect 42856 21732 42912 21788
rect 42912 21732 42916 21788
rect 42852 21728 42916 21732
rect 47612 21788 47676 21792
rect 47612 21732 47616 21788
rect 47616 21732 47672 21788
rect 47672 21732 47676 21788
rect 47612 21728 47676 21732
rect 47692 21788 47756 21792
rect 47692 21732 47696 21788
rect 47696 21732 47752 21788
rect 47752 21732 47756 21788
rect 47692 21728 47756 21732
rect 47772 21788 47836 21792
rect 47772 21732 47776 21788
rect 47776 21732 47832 21788
rect 47832 21732 47836 21788
rect 47772 21728 47836 21732
rect 47852 21788 47916 21792
rect 47852 21732 47856 21788
rect 47856 21732 47912 21788
rect 47912 21732 47916 21788
rect 47852 21728 47916 21732
rect 52612 21788 52676 21792
rect 52612 21732 52616 21788
rect 52616 21732 52672 21788
rect 52672 21732 52676 21788
rect 52612 21728 52676 21732
rect 52692 21788 52756 21792
rect 52692 21732 52696 21788
rect 52696 21732 52752 21788
rect 52752 21732 52756 21788
rect 52692 21728 52756 21732
rect 52772 21788 52836 21792
rect 52772 21732 52776 21788
rect 52776 21732 52832 21788
rect 52832 21732 52836 21788
rect 52772 21728 52836 21732
rect 52852 21788 52916 21792
rect 52852 21732 52856 21788
rect 52856 21732 52912 21788
rect 52912 21732 52916 21788
rect 52852 21728 52916 21732
rect 57612 21788 57676 21792
rect 57612 21732 57616 21788
rect 57616 21732 57672 21788
rect 57672 21732 57676 21788
rect 57612 21728 57676 21732
rect 57692 21788 57756 21792
rect 57692 21732 57696 21788
rect 57696 21732 57752 21788
rect 57752 21732 57756 21788
rect 57692 21728 57756 21732
rect 57772 21788 57836 21792
rect 57772 21732 57776 21788
rect 57776 21732 57832 21788
rect 57832 21732 57836 21788
rect 57772 21728 57836 21732
rect 57852 21788 57916 21792
rect 57852 21732 57856 21788
rect 57856 21732 57912 21788
rect 57912 21732 57916 21788
rect 57852 21728 57916 21732
rect 1952 21244 2016 21248
rect 1952 21188 1956 21244
rect 1956 21188 2012 21244
rect 2012 21188 2016 21244
rect 1952 21184 2016 21188
rect 2032 21244 2096 21248
rect 2032 21188 2036 21244
rect 2036 21188 2092 21244
rect 2092 21188 2096 21244
rect 2032 21184 2096 21188
rect 2112 21244 2176 21248
rect 2112 21188 2116 21244
rect 2116 21188 2172 21244
rect 2172 21188 2176 21244
rect 2112 21184 2176 21188
rect 2192 21244 2256 21248
rect 2192 21188 2196 21244
rect 2196 21188 2252 21244
rect 2252 21188 2256 21244
rect 2192 21184 2256 21188
rect 6952 21244 7016 21248
rect 6952 21188 6956 21244
rect 6956 21188 7012 21244
rect 7012 21188 7016 21244
rect 6952 21184 7016 21188
rect 7032 21244 7096 21248
rect 7032 21188 7036 21244
rect 7036 21188 7092 21244
rect 7092 21188 7096 21244
rect 7032 21184 7096 21188
rect 7112 21244 7176 21248
rect 7112 21188 7116 21244
rect 7116 21188 7172 21244
rect 7172 21188 7176 21244
rect 7112 21184 7176 21188
rect 7192 21244 7256 21248
rect 7192 21188 7196 21244
rect 7196 21188 7252 21244
rect 7252 21188 7256 21244
rect 7192 21184 7256 21188
rect 11952 21244 12016 21248
rect 11952 21188 11956 21244
rect 11956 21188 12012 21244
rect 12012 21188 12016 21244
rect 11952 21184 12016 21188
rect 12032 21244 12096 21248
rect 12032 21188 12036 21244
rect 12036 21188 12092 21244
rect 12092 21188 12096 21244
rect 12032 21184 12096 21188
rect 12112 21244 12176 21248
rect 12112 21188 12116 21244
rect 12116 21188 12172 21244
rect 12172 21188 12176 21244
rect 12112 21184 12176 21188
rect 12192 21244 12256 21248
rect 12192 21188 12196 21244
rect 12196 21188 12252 21244
rect 12252 21188 12256 21244
rect 12192 21184 12256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 21952 21244 22016 21248
rect 21952 21188 21956 21244
rect 21956 21188 22012 21244
rect 22012 21188 22016 21244
rect 21952 21184 22016 21188
rect 22032 21244 22096 21248
rect 22032 21188 22036 21244
rect 22036 21188 22092 21244
rect 22092 21188 22096 21244
rect 22032 21184 22096 21188
rect 22112 21244 22176 21248
rect 22112 21188 22116 21244
rect 22116 21188 22172 21244
rect 22172 21188 22176 21244
rect 22112 21184 22176 21188
rect 22192 21244 22256 21248
rect 22192 21188 22196 21244
rect 22196 21188 22252 21244
rect 22252 21188 22256 21244
rect 22192 21184 22256 21188
rect 26952 21244 27016 21248
rect 26952 21188 26956 21244
rect 26956 21188 27012 21244
rect 27012 21188 27016 21244
rect 26952 21184 27016 21188
rect 27032 21244 27096 21248
rect 27032 21188 27036 21244
rect 27036 21188 27092 21244
rect 27092 21188 27096 21244
rect 27032 21184 27096 21188
rect 27112 21244 27176 21248
rect 27112 21188 27116 21244
rect 27116 21188 27172 21244
rect 27172 21188 27176 21244
rect 27112 21184 27176 21188
rect 27192 21244 27256 21248
rect 27192 21188 27196 21244
rect 27196 21188 27252 21244
rect 27252 21188 27256 21244
rect 27192 21184 27256 21188
rect 31952 21244 32016 21248
rect 31952 21188 31956 21244
rect 31956 21188 32012 21244
rect 32012 21188 32016 21244
rect 31952 21184 32016 21188
rect 32032 21244 32096 21248
rect 32032 21188 32036 21244
rect 32036 21188 32092 21244
rect 32092 21188 32096 21244
rect 32032 21184 32096 21188
rect 32112 21244 32176 21248
rect 32112 21188 32116 21244
rect 32116 21188 32172 21244
rect 32172 21188 32176 21244
rect 32112 21184 32176 21188
rect 32192 21244 32256 21248
rect 32192 21188 32196 21244
rect 32196 21188 32252 21244
rect 32252 21188 32256 21244
rect 32192 21184 32256 21188
rect 36952 21244 37016 21248
rect 36952 21188 36956 21244
rect 36956 21188 37012 21244
rect 37012 21188 37016 21244
rect 36952 21184 37016 21188
rect 37032 21244 37096 21248
rect 37032 21188 37036 21244
rect 37036 21188 37092 21244
rect 37092 21188 37096 21244
rect 37032 21184 37096 21188
rect 37112 21244 37176 21248
rect 37112 21188 37116 21244
rect 37116 21188 37172 21244
rect 37172 21188 37176 21244
rect 37112 21184 37176 21188
rect 37192 21244 37256 21248
rect 37192 21188 37196 21244
rect 37196 21188 37252 21244
rect 37252 21188 37256 21244
rect 37192 21184 37256 21188
rect 41952 21244 42016 21248
rect 41952 21188 41956 21244
rect 41956 21188 42012 21244
rect 42012 21188 42016 21244
rect 41952 21184 42016 21188
rect 42032 21244 42096 21248
rect 42032 21188 42036 21244
rect 42036 21188 42092 21244
rect 42092 21188 42096 21244
rect 42032 21184 42096 21188
rect 42112 21244 42176 21248
rect 42112 21188 42116 21244
rect 42116 21188 42172 21244
rect 42172 21188 42176 21244
rect 42112 21184 42176 21188
rect 42192 21244 42256 21248
rect 42192 21188 42196 21244
rect 42196 21188 42252 21244
rect 42252 21188 42256 21244
rect 42192 21184 42256 21188
rect 46952 21244 47016 21248
rect 46952 21188 46956 21244
rect 46956 21188 47012 21244
rect 47012 21188 47016 21244
rect 46952 21184 47016 21188
rect 47032 21244 47096 21248
rect 47032 21188 47036 21244
rect 47036 21188 47092 21244
rect 47092 21188 47096 21244
rect 47032 21184 47096 21188
rect 47112 21244 47176 21248
rect 47112 21188 47116 21244
rect 47116 21188 47172 21244
rect 47172 21188 47176 21244
rect 47112 21184 47176 21188
rect 47192 21244 47256 21248
rect 47192 21188 47196 21244
rect 47196 21188 47252 21244
rect 47252 21188 47256 21244
rect 47192 21184 47256 21188
rect 51952 21244 52016 21248
rect 51952 21188 51956 21244
rect 51956 21188 52012 21244
rect 52012 21188 52016 21244
rect 51952 21184 52016 21188
rect 52032 21244 52096 21248
rect 52032 21188 52036 21244
rect 52036 21188 52092 21244
rect 52092 21188 52096 21244
rect 52032 21184 52096 21188
rect 52112 21244 52176 21248
rect 52112 21188 52116 21244
rect 52116 21188 52172 21244
rect 52172 21188 52176 21244
rect 52112 21184 52176 21188
rect 52192 21244 52256 21248
rect 52192 21188 52196 21244
rect 52196 21188 52252 21244
rect 52252 21188 52256 21244
rect 52192 21184 52256 21188
rect 56952 21244 57016 21248
rect 56952 21188 56956 21244
rect 56956 21188 57012 21244
rect 57012 21188 57016 21244
rect 56952 21184 57016 21188
rect 57032 21244 57096 21248
rect 57032 21188 57036 21244
rect 57036 21188 57092 21244
rect 57092 21188 57096 21244
rect 57032 21184 57096 21188
rect 57112 21244 57176 21248
rect 57112 21188 57116 21244
rect 57116 21188 57172 21244
rect 57172 21188 57176 21244
rect 57112 21184 57176 21188
rect 57192 21244 57256 21248
rect 57192 21188 57196 21244
rect 57196 21188 57252 21244
rect 57252 21188 57256 21244
rect 57192 21184 57256 21188
rect 2612 20700 2676 20704
rect 2612 20644 2616 20700
rect 2616 20644 2672 20700
rect 2672 20644 2676 20700
rect 2612 20640 2676 20644
rect 2692 20700 2756 20704
rect 2692 20644 2696 20700
rect 2696 20644 2752 20700
rect 2752 20644 2756 20700
rect 2692 20640 2756 20644
rect 2772 20700 2836 20704
rect 2772 20644 2776 20700
rect 2776 20644 2832 20700
rect 2832 20644 2836 20700
rect 2772 20640 2836 20644
rect 2852 20700 2916 20704
rect 2852 20644 2856 20700
rect 2856 20644 2912 20700
rect 2912 20644 2916 20700
rect 2852 20640 2916 20644
rect 7612 20700 7676 20704
rect 7612 20644 7616 20700
rect 7616 20644 7672 20700
rect 7672 20644 7676 20700
rect 7612 20640 7676 20644
rect 7692 20700 7756 20704
rect 7692 20644 7696 20700
rect 7696 20644 7752 20700
rect 7752 20644 7756 20700
rect 7692 20640 7756 20644
rect 7772 20700 7836 20704
rect 7772 20644 7776 20700
rect 7776 20644 7832 20700
rect 7832 20644 7836 20700
rect 7772 20640 7836 20644
rect 7852 20700 7916 20704
rect 7852 20644 7856 20700
rect 7856 20644 7912 20700
rect 7912 20644 7916 20700
rect 7852 20640 7916 20644
rect 12612 20700 12676 20704
rect 12612 20644 12616 20700
rect 12616 20644 12672 20700
rect 12672 20644 12676 20700
rect 12612 20640 12676 20644
rect 12692 20700 12756 20704
rect 12692 20644 12696 20700
rect 12696 20644 12752 20700
rect 12752 20644 12756 20700
rect 12692 20640 12756 20644
rect 12772 20700 12836 20704
rect 12772 20644 12776 20700
rect 12776 20644 12832 20700
rect 12832 20644 12836 20700
rect 12772 20640 12836 20644
rect 12852 20700 12916 20704
rect 12852 20644 12856 20700
rect 12856 20644 12912 20700
rect 12912 20644 12916 20700
rect 12852 20640 12916 20644
rect 17612 20700 17676 20704
rect 17612 20644 17616 20700
rect 17616 20644 17672 20700
rect 17672 20644 17676 20700
rect 17612 20640 17676 20644
rect 17692 20700 17756 20704
rect 17692 20644 17696 20700
rect 17696 20644 17752 20700
rect 17752 20644 17756 20700
rect 17692 20640 17756 20644
rect 17772 20700 17836 20704
rect 17772 20644 17776 20700
rect 17776 20644 17832 20700
rect 17832 20644 17836 20700
rect 17772 20640 17836 20644
rect 17852 20700 17916 20704
rect 17852 20644 17856 20700
rect 17856 20644 17912 20700
rect 17912 20644 17916 20700
rect 17852 20640 17916 20644
rect 22612 20700 22676 20704
rect 22612 20644 22616 20700
rect 22616 20644 22672 20700
rect 22672 20644 22676 20700
rect 22612 20640 22676 20644
rect 22692 20700 22756 20704
rect 22692 20644 22696 20700
rect 22696 20644 22752 20700
rect 22752 20644 22756 20700
rect 22692 20640 22756 20644
rect 22772 20700 22836 20704
rect 22772 20644 22776 20700
rect 22776 20644 22832 20700
rect 22832 20644 22836 20700
rect 22772 20640 22836 20644
rect 22852 20700 22916 20704
rect 22852 20644 22856 20700
rect 22856 20644 22912 20700
rect 22912 20644 22916 20700
rect 22852 20640 22916 20644
rect 27612 20700 27676 20704
rect 27612 20644 27616 20700
rect 27616 20644 27672 20700
rect 27672 20644 27676 20700
rect 27612 20640 27676 20644
rect 27692 20700 27756 20704
rect 27692 20644 27696 20700
rect 27696 20644 27752 20700
rect 27752 20644 27756 20700
rect 27692 20640 27756 20644
rect 27772 20700 27836 20704
rect 27772 20644 27776 20700
rect 27776 20644 27832 20700
rect 27832 20644 27836 20700
rect 27772 20640 27836 20644
rect 27852 20700 27916 20704
rect 27852 20644 27856 20700
rect 27856 20644 27912 20700
rect 27912 20644 27916 20700
rect 27852 20640 27916 20644
rect 32612 20700 32676 20704
rect 32612 20644 32616 20700
rect 32616 20644 32672 20700
rect 32672 20644 32676 20700
rect 32612 20640 32676 20644
rect 32692 20700 32756 20704
rect 32692 20644 32696 20700
rect 32696 20644 32752 20700
rect 32752 20644 32756 20700
rect 32692 20640 32756 20644
rect 32772 20700 32836 20704
rect 32772 20644 32776 20700
rect 32776 20644 32832 20700
rect 32832 20644 32836 20700
rect 32772 20640 32836 20644
rect 32852 20700 32916 20704
rect 32852 20644 32856 20700
rect 32856 20644 32912 20700
rect 32912 20644 32916 20700
rect 32852 20640 32916 20644
rect 37612 20700 37676 20704
rect 37612 20644 37616 20700
rect 37616 20644 37672 20700
rect 37672 20644 37676 20700
rect 37612 20640 37676 20644
rect 37692 20700 37756 20704
rect 37692 20644 37696 20700
rect 37696 20644 37752 20700
rect 37752 20644 37756 20700
rect 37692 20640 37756 20644
rect 37772 20700 37836 20704
rect 37772 20644 37776 20700
rect 37776 20644 37832 20700
rect 37832 20644 37836 20700
rect 37772 20640 37836 20644
rect 37852 20700 37916 20704
rect 37852 20644 37856 20700
rect 37856 20644 37912 20700
rect 37912 20644 37916 20700
rect 37852 20640 37916 20644
rect 42612 20700 42676 20704
rect 42612 20644 42616 20700
rect 42616 20644 42672 20700
rect 42672 20644 42676 20700
rect 42612 20640 42676 20644
rect 42692 20700 42756 20704
rect 42692 20644 42696 20700
rect 42696 20644 42752 20700
rect 42752 20644 42756 20700
rect 42692 20640 42756 20644
rect 42772 20700 42836 20704
rect 42772 20644 42776 20700
rect 42776 20644 42832 20700
rect 42832 20644 42836 20700
rect 42772 20640 42836 20644
rect 42852 20700 42916 20704
rect 42852 20644 42856 20700
rect 42856 20644 42912 20700
rect 42912 20644 42916 20700
rect 42852 20640 42916 20644
rect 47612 20700 47676 20704
rect 47612 20644 47616 20700
rect 47616 20644 47672 20700
rect 47672 20644 47676 20700
rect 47612 20640 47676 20644
rect 47692 20700 47756 20704
rect 47692 20644 47696 20700
rect 47696 20644 47752 20700
rect 47752 20644 47756 20700
rect 47692 20640 47756 20644
rect 47772 20700 47836 20704
rect 47772 20644 47776 20700
rect 47776 20644 47832 20700
rect 47832 20644 47836 20700
rect 47772 20640 47836 20644
rect 47852 20700 47916 20704
rect 47852 20644 47856 20700
rect 47856 20644 47912 20700
rect 47912 20644 47916 20700
rect 47852 20640 47916 20644
rect 52612 20700 52676 20704
rect 52612 20644 52616 20700
rect 52616 20644 52672 20700
rect 52672 20644 52676 20700
rect 52612 20640 52676 20644
rect 52692 20700 52756 20704
rect 52692 20644 52696 20700
rect 52696 20644 52752 20700
rect 52752 20644 52756 20700
rect 52692 20640 52756 20644
rect 52772 20700 52836 20704
rect 52772 20644 52776 20700
rect 52776 20644 52832 20700
rect 52832 20644 52836 20700
rect 52772 20640 52836 20644
rect 52852 20700 52916 20704
rect 52852 20644 52856 20700
rect 52856 20644 52912 20700
rect 52912 20644 52916 20700
rect 52852 20640 52916 20644
rect 57612 20700 57676 20704
rect 57612 20644 57616 20700
rect 57616 20644 57672 20700
rect 57672 20644 57676 20700
rect 57612 20640 57676 20644
rect 57692 20700 57756 20704
rect 57692 20644 57696 20700
rect 57696 20644 57752 20700
rect 57752 20644 57756 20700
rect 57692 20640 57756 20644
rect 57772 20700 57836 20704
rect 57772 20644 57776 20700
rect 57776 20644 57832 20700
rect 57832 20644 57836 20700
rect 57772 20640 57836 20644
rect 57852 20700 57916 20704
rect 57852 20644 57856 20700
rect 57856 20644 57912 20700
rect 57912 20644 57916 20700
rect 57852 20640 57916 20644
rect 1952 20156 2016 20160
rect 1952 20100 1956 20156
rect 1956 20100 2012 20156
rect 2012 20100 2016 20156
rect 1952 20096 2016 20100
rect 2032 20156 2096 20160
rect 2032 20100 2036 20156
rect 2036 20100 2092 20156
rect 2092 20100 2096 20156
rect 2032 20096 2096 20100
rect 2112 20156 2176 20160
rect 2112 20100 2116 20156
rect 2116 20100 2172 20156
rect 2172 20100 2176 20156
rect 2112 20096 2176 20100
rect 2192 20156 2256 20160
rect 2192 20100 2196 20156
rect 2196 20100 2252 20156
rect 2252 20100 2256 20156
rect 2192 20096 2256 20100
rect 6952 20156 7016 20160
rect 6952 20100 6956 20156
rect 6956 20100 7012 20156
rect 7012 20100 7016 20156
rect 6952 20096 7016 20100
rect 7032 20156 7096 20160
rect 7032 20100 7036 20156
rect 7036 20100 7092 20156
rect 7092 20100 7096 20156
rect 7032 20096 7096 20100
rect 7112 20156 7176 20160
rect 7112 20100 7116 20156
rect 7116 20100 7172 20156
rect 7172 20100 7176 20156
rect 7112 20096 7176 20100
rect 7192 20156 7256 20160
rect 7192 20100 7196 20156
rect 7196 20100 7252 20156
rect 7252 20100 7256 20156
rect 7192 20096 7256 20100
rect 11952 20156 12016 20160
rect 11952 20100 11956 20156
rect 11956 20100 12012 20156
rect 12012 20100 12016 20156
rect 11952 20096 12016 20100
rect 12032 20156 12096 20160
rect 12032 20100 12036 20156
rect 12036 20100 12092 20156
rect 12092 20100 12096 20156
rect 12032 20096 12096 20100
rect 12112 20156 12176 20160
rect 12112 20100 12116 20156
rect 12116 20100 12172 20156
rect 12172 20100 12176 20156
rect 12112 20096 12176 20100
rect 12192 20156 12256 20160
rect 12192 20100 12196 20156
rect 12196 20100 12252 20156
rect 12252 20100 12256 20156
rect 12192 20096 12256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 21952 20156 22016 20160
rect 21952 20100 21956 20156
rect 21956 20100 22012 20156
rect 22012 20100 22016 20156
rect 21952 20096 22016 20100
rect 22032 20156 22096 20160
rect 22032 20100 22036 20156
rect 22036 20100 22092 20156
rect 22092 20100 22096 20156
rect 22032 20096 22096 20100
rect 22112 20156 22176 20160
rect 22112 20100 22116 20156
rect 22116 20100 22172 20156
rect 22172 20100 22176 20156
rect 22112 20096 22176 20100
rect 22192 20156 22256 20160
rect 22192 20100 22196 20156
rect 22196 20100 22252 20156
rect 22252 20100 22256 20156
rect 22192 20096 22256 20100
rect 26952 20156 27016 20160
rect 26952 20100 26956 20156
rect 26956 20100 27012 20156
rect 27012 20100 27016 20156
rect 26952 20096 27016 20100
rect 27032 20156 27096 20160
rect 27032 20100 27036 20156
rect 27036 20100 27092 20156
rect 27092 20100 27096 20156
rect 27032 20096 27096 20100
rect 27112 20156 27176 20160
rect 27112 20100 27116 20156
rect 27116 20100 27172 20156
rect 27172 20100 27176 20156
rect 27112 20096 27176 20100
rect 27192 20156 27256 20160
rect 27192 20100 27196 20156
rect 27196 20100 27252 20156
rect 27252 20100 27256 20156
rect 27192 20096 27256 20100
rect 31952 20156 32016 20160
rect 31952 20100 31956 20156
rect 31956 20100 32012 20156
rect 32012 20100 32016 20156
rect 31952 20096 32016 20100
rect 32032 20156 32096 20160
rect 32032 20100 32036 20156
rect 32036 20100 32092 20156
rect 32092 20100 32096 20156
rect 32032 20096 32096 20100
rect 32112 20156 32176 20160
rect 32112 20100 32116 20156
rect 32116 20100 32172 20156
rect 32172 20100 32176 20156
rect 32112 20096 32176 20100
rect 32192 20156 32256 20160
rect 32192 20100 32196 20156
rect 32196 20100 32252 20156
rect 32252 20100 32256 20156
rect 32192 20096 32256 20100
rect 36952 20156 37016 20160
rect 36952 20100 36956 20156
rect 36956 20100 37012 20156
rect 37012 20100 37016 20156
rect 36952 20096 37016 20100
rect 37032 20156 37096 20160
rect 37032 20100 37036 20156
rect 37036 20100 37092 20156
rect 37092 20100 37096 20156
rect 37032 20096 37096 20100
rect 37112 20156 37176 20160
rect 37112 20100 37116 20156
rect 37116 20100 37172 20156
rect 37172 20100 37176 20156
rect 37112 20096 37176 20100
rect 37192 20156 37256 20160
rect 37192 20100 37196 20156
rect 37196 20100 37252 20156
rect 37252 20100 37256 20156
rect 37192 20096 37256 20100
rect 41952 20156 42016 20160
rect 41952 20100 41956 20156
rect 41956 20100 42012 20156
rect 42012 20100 42016 20156
rect 41952 20096 42016 20100
rect 42032 20156 42096 20160
rect 42032 20100 42036 20156
rect 42036 20100 42092 20156
rect 42092 20100 42096 20156
rect 42032 20096 42096 20100
rect 42112 20156 42176 20160
rect 42112 20100 42116 20156
rect 42116 20100 42172 20156
rect 42172 20100 42176 20156
rect 42112 20096 42176 20100
rect 42192 20156 42256 20160
rect 42192 20100 42196 20156
rect 42196 20100 42252 20156
rect 42252 20100 42256 20156
rect 42192 20096 42256 20100
rect 46952 20156 47016 20160
rect 46952 20100 46956 20156
rect 46956 20100 47012 20156
rect 47012 20100 47016 20156
rect 46952 20096 47016 20100
rect 47032 20156 47096 20160
rect 47032 20100 47036 20156
rect 47036 20100 47092 20156
rect 47092 20100 47096 20156
rect 47032 20096 47096 20100
rect 47112 20156 47176 20160
rect 47112 20100 47116 20156
rect 47116 20100 47172 20156
rect 47172 20100 47176 20156
rect 47112 20096 47176 20100
rect 47192 20156 47256 20160
rect 47192 20100 47196 20156
rect 47196 20100 47252 20156
rect 47252 20100 47256 20156
rect 47192 20096 47256 20100
rect 51952 20156 52016 20160
rect 51952 20100 51956 20156
rect 51956 20100 52012 20156
rect 52012 20100 52016 20156
rect 51952 20096 52016 20100
rect 52032 20156 52096 20160
rect 52032 20100 52036 20156
rect 52036 20100 52092 20156
rect 52092 20100 52096 20156
rect 52032 20096 52096 20100
rect 52112 20156 52176 20160
rect 52112 20100 52116 20156
rect 52116 20100 52172 20156
rect 52172 20100 52176 20156
rect 52112 20096 52176 20100
rect 52192 20156 52256 20160
rect 52192 20100 52196 20156
rect 52196 20100 52252 20156
rect 52252 20100 52256 20156
rect 52192 20096 52256 20100
rect 56952 20156 57016 20160
rect 56952 20100 56956 20156
rect 56956 20100 57012 20156
rect 57012 20100 57016 20156
rect 56952 20096 57016 20100
rect 57032 20156 57096 20160
rect 57032 20100 57036 20156
rect 57036 20100 57092 20156
rect 57092 20100 57096 20156
rect 57032 20096 57096 20100
rect 57112 20156 57176 20160
rect 57112 20100 57116 20156
rect 57116 20100 57172 20156
rect 57172 20100 57176 20156
rect 57112 20096 57176 20100
rect 57192 20156 57256 20160
rect 57192 20100 57196 20156
rect 57196 20100 57252 20156
rect 57252 20100 57256 20156
rect 57192 20096 57256 20100
rect 2612 19612 2676 19616
rect 2612 19556 2616 19612
rect 2616 19556 2672 19612
rect 2672 19556 2676 19612
rect 2612 19552 2676 19556
rect 2692 19612 2756 19616
rect 2692 19556 2696 19612
rect 2696 19556 2752 19612
rect 2752 19556 2756 19612
rect 2692 19552 2756 19556
rect 2772 19612 2836 19616
rect 2772 19556 2776 19612
rect 2776 19556 2832 19612
rect 2832 19556 2836 19612
rect 2772 19552 2836 19556
rect 2852 19612 2916 19616
rect 2852 19556 2856 19612
rect 2856 19556 2912 19612
rect 2912 19556 2916 19612
rect 2852 19552 2916 19556
rect 7612 19612 7676 19616
rect 7612 19556 7616 19612
rect 7616 19556 7672 19612
rect 7672 19556 7676 19612
rect 7612 19552 7676 19556
rect 7692 19612 7756 19616
rect 7692 19556 7696 19612
rect 7696 19556 7752 19612
rect 7752 19556 7756 19612
rect 7692 19552 7756 19556
rect 7772 19612 7836 19616
rect 7772 19556 7776 19612
rect 7776 19556 7832 19612
rect 7832 19556 7836 19612
rect 7772 19552 7836 19556
rect 7852 19612 7916 19616
rect 7852 19556 7856 19612
rect 7856 19556 7912 19612
rect 7912 19556 7916 19612
rect 7852 19552 7916 19556
rect 12612 19612 12676 19616
rect 12612 19556 12616 19612
rect 12616 19556 12672 19612
rect 12672 19556 12676 19612
rect 12612 19552 12676 19556
rect 12692 19612 12756 19616
rect 12692 19556 12696 19612
rect 12696 19556 12752 19612
rect 12752 19556 12756 19612
rect 12692 19552 12756 19556
rect 12772 19612 12836 19616
rect 12772 19556 12776 19612
rect 12776 19556 12832 19612
rect 12832 19556 12836 19612
rect 12772 19552 12836 19556
rect 12852 19612 12916 19616
rect 12852 19556 12856 19612
rect 12856 19556 12912 19612
rect 12912 19556 12916 19612
rect 12852 19552 12916 19556
rect 17612 19612 17676 19616
rect 17612 19556 17616 19612
rect 17616 19556 17672 19612
rect 17672 19556 17676 19612
rect 17612 19552 17676 19556
rect 17692 19612 17756 19616
rect 17692 19556 17696 19612
rect 17696 19556 17752 19612
rect 17752 19556 17756 19612
rect 17692 19552 17756 19556
rect 17772 19612 17836 19616
rect 17772 19556 17776 19612
rect 17776 19556 17832 19612
rect 17832 19556 17836 19612
rect 17772 19552 17836 19556
rect 17852 19612 17916 19616
rect 17852 19556 17856 19612
rect 17856 19556 17912 19612
rect 17912 19556 17916 19612
rect 17852 19552 17916 19556
rect 22612 19612 22676 19616
rect 22612 19556 22616 19612
rect 22616 19556 22672 19612
rect 22672 19556 22676 19612
rect 22612 19552 22676 19556
rect 22692 19612 22756 19616
rect 22692 19556 22696 19612
rect 22696 19556 22752 19612
rect 22752 19556 22756 19612
rect 22692 19552 22756 19556
rect 22772 19612 22836 19616
rect 22772 19556 22776 19612
rect 22776 19556 22832 19612
rect 22832 19556 22836 19612
rect 22772 19552 22836 19556
rect 22852 19612 22916 19616
rect 22852 19556 22856 19612
rect 22856 19556 22912 19612
rect 22912 19556 22916 19612
rect 22852 19552 22916 19556
rect 27612 19612 27676 19616
rect 27612 19556 27616 19612
rect 27616 19556 27672 19612
rect 27672 19556 27676 19612
rect 27612 19552 27676 19556
rect 27692 19612 27756 19616
rect 27692 19556 27696 19612
rect 27696 19556 27752 19612
rect 27752 19556 27756 19612
rect 27692 19552 27756 19556
rect 27772 19612 27836 19616
rect 27772 19556 27776 19612
rect 27776 19556 27832 19612
rect 27832 19556 27836 19612
rect 27772 19552 27836 19556
rect 27852 19612 27916 19616
rect 27852 19556 27856 19612
rect 27856 19556 27912 19612
rect 27912 19556 27916 19612
rect 27852 19552 27916 19556
rect 32612 19612 32676 19616
rect 32612 19556 32616 19612
rect 32616 19556 32672 19612
rect 32672 19556 32676 19612
rect 32612 19552 32676 19556
rect 32692 19612 32756 19616
rect 32692 19556 32696 19612
rect 32696 19556 32752 19612
rect 32752 19556 32756 19612
rect 32692 19552 32756 19556
rect 32772 19612 32836 19616
rect 32772 19556 32776 19612
rect 32776 19556 32832 19612
rect 32832 19556 32836 19612
rect 32772 19552 32836 19556
rect 32852 19612 32916 19616
rect 32852 19556 32856 19612
rect 32856 19556 32912 19612
rect 32912 19556 32916 19612
rect 32852 19552 32916 19556
rect 37612 19612 37676 19616
rect 37612 19556 37616 19612
rect 37616 19556 37672 19612
rect 37672 19556 37676 19612
rect 37612 19552 37676 19556
rect 37692 19612 37756 19616
rect 37692 19556 37696 19612
rect 37696 19556 37752 19612
rect 37752 19556 37756 19612
rect 37692 19552 37756 19556
rect 37772 19612 37836 19616
rect 37772 19556 37776 19612
rect 37776 19556 37832 19612
rect 37832 19556 37836 19612
rect 37772 19552 37836 19556
rect 37852 19612 37916 19616
rect 37852 19556 37856 19612
rect 37856 19556 37912 19612
rect 37912 19556 37916 19612
rect 37852 19552 37916 19556
rect 42612 19612 42676 19616
rect 42612 19556 42616 19612
rect 42616 19556 42672 19612
rect 42672 19556 42676 19612
rect 42612 19552 42676 19556
rect 42692 19612 42756 19616
rect 42692 19556 42696 19612
rect 42696 19556 42752 19612
rect 42752 19556 42756 19612
rect 42692 19552 42756 19556
rect 42772 19612 42836 19616
rect 42772 19556 42776 19612
rect 42776 19556 42832 19612
rect 42832 19556 42836 19612
rect 42772 19552 42836 19556
rect 42852 19612 42916 19616
rect 42852 19556 42856 19612
rect 42856 19556 42912 19612
rect 42912 19556 42916 19612
rect 42852 19552 42916 19556
rect 47612 19612 47676 19616
rect 47612 19556 47616 19612
rect 47616 19556 47672 19612
rect 47672 19556 47676 19612
rect 47612 19552 47676 19556
rect 47692 19612 47756 19616
rect 47692 19556 47696 19612
rect 47696 19556 47752 19612
rect 47752 19556 47756 19612
rect 47692 19552 47756 19556
rect 47772 19612 47836 19616
rect 47772 19556 47776 19612
rect 47776 19556 47832 19612
rect 47832 19556 47836 19612
rect 47772 19552 47836 19556
rect 47852 19612 47916 19616
rect 47852 19556 47856 19612
rect 47856 19556 47912 19612
rect 47912 19556 47916 19612
rect 47852 19552 47916 19556
rect 52612 19612 52676 19616
rect 52612 19556 52616 19612
rect 52616 19556 52672 19612
rect 52672 19556 52676 19612
rect 52612 19552 52676 19556
rect 52692 19612 52756 19616
rect 52692 19556 52696 19612
rect 52696 19556 52752 19612
rect 52752 19556 52756 19612
rect 52692 19552 52756 19556
rect 52772 19612 52836 19616
rect 52772 19556 52776 19612
rect 52776 19556 52832 19612
rect 52832 19556 52836 19612
rect 52772 19552 52836 19556
rect 52852 19612 52916 19616
rect 52852 19556 52856 19612
rect 52856 19556 52912 19612
rect 52912 19556 52916 19612
rect 52852 19552 52916 19556
rect 57612 19612 57676 19616
rect 57612 19556 57616 19612
rect 57616 19556 57672 19612
rect 57672 19556 57676 19612
rect 57612 19552 57676 19556
rect 57692 19612 57756 19616
rect 57692 19556 57696 19612
rect 57696 19556 57752 19612
rect 57752 19556 57756 19612
rect 57692 19552 57756 19556
rect 57772 19612 57836 19616
rect 57772 19556 57776 19612
rect 57776 19556 57832 19612
rect 57832 19556 57836 19612
rect 57772 19552 57836 19556
rect 57852 19612 57916 19616
rect 57852 19556 57856 19612
rect 57856 19556 57912 19612
rect 57912 19556 57916 19612
rect 57852 19552 57916 19556
rect 1952 19068 2016 19072
rect 1952 19012 1956 19068
rect 1956 19012 2012 19068
rect 2012 19012 2016 19068
rect 1952 19008 2016 19012
rect 2032 19068 2096 19072
rect 2032 19012 2036 19068
rect 2036 19012 2092 19068
rect 2092 19012 2096 19068
rect 2032 19008 2096 19012
rect 2112 19068 2176 19072
rect 2112 19012 2116 19068
rect 2116 19012 2172 19068
rect 2172 19012 2176 19068
rect 2112 19008 2176 19012
rect 2192 19068 2256 19072
rect 2192 19012 2196 19068
rect 2196 19012 2252 19068
rect 2252 19012 2256 19068
rect 2192 19008 2256 19012
rect 6952 19068 7016 19072
rect 6952 19012 6956 19068
rect 6956 19012 7012 19068
rect 7012 19012 7016 19068
rect 6952 19008 7016 19012
rect 7032 19068 7096 19072
rect 7032 19012 7036 19068
rect 7036 19012 7092 19068
rect 7092 19012 7096 19068
rect 7032 19008 7096 19012
rect 7112 19068 7176 19072
rect 7112 19012 7116 19068
rect 7116 19012 7172 19068
rect 7172 19012 7176 19068
rect 7112 19008 7176 19012
rect 7192 19068 7256 19072
rect 7192 19012 7196 19068
rect 7196 19012 7252 19068
rect 7252 19012 7256 19068
rect 7192 19008 7256 19012
rect 11952 19068 12016 19072
rect 11952 19012 11956 19068
rect 11956 19012 12012 19068
rect 12012 19012 12016 19068
rect 11952 19008 12016 19012
rect 12032 19068 12096 19072
rect 12032 19012 12036 19068
rect 12036 19012 12092 19068
rect 12092 19012 12096 19068
rect 12032 19008 12096 19012
rect 12112 19068 12176 19072
rect 12112 19012 12116 19068
rect 12116 19012 12172 19068
rect 12172 19012 12176 19068
rect 12112 19008 12176 19012
rect 12192 19068 12256 19072
rect 12192 19012 12196 19068
rect 12196 19012 12252 19068
rect 12252 19012 12256 19068
rect 12192 19008 12256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 21952 19068 22016 19072
rect 21952 19012 21956 19068
rect 21956 19012 22012 19068
rect 22012 19012 22016 19068
rect 21952 19008 22016 19012
rect 22032 19068 22096 19072
rect 22032 19012 22036 19068
rect 22036 19012 22092 19068
rect 22092 19012 22096 19068
rect 22032 19008 22096 19012
rect 22112 19068 22176 19072
rect 22112 19012 22116 19068
rect 22116 19012 22172 19068
rect 22172 19012 22176 19068
rect 22112 19008 22176 19012
rect 22192 19068 22256 19072
rect 22192 19012 22196 19068
rect 22196 19012 22252 19068
rect 22252 19012 22256 19068
rect 22192 19008 22256 19012
rect 26952 19068 27016 19072
rect 26952 19012 26956 19068
rect 26956 19012 27012 19068
rect 27012 19012 27016 19068
rect 26952 19008 27016 19012
rect 27032 19068 27096 19072
rect 27032 19012 27036 19068
rect 27036 19012 27092 19068
rect 27092 19012 27096 19068
rect 27032 19008 27096 19012
rect 27112 19068 27176 19072
rect 27112 19012 27116 19068
rect 27116 19012 27172 19068
rect 27172 19012 27176 19068
rect 27112 19008 27176 19012
rect 27192 19068 27256 19072
rect 27192 19012 27196 19068
rect 27196 19012 27252 19068
rect 27252 19012 27256 19068
rect 27192 19008 27256 19012
rect 31952 19068 32016 19072
rect 31952 19012 31956 19068
rect 31956 19012 32012 19068
rect 32012 19012 32016 19068
rect 31952 19008 32016 19012
rect 32032 19068 32096 19072
rect 32032 19012 32036 19068
rect 32036 19012 32092 19068
rect 32092 19012 32096 19068
rect 32032 19008 32096 19012
rect 32112 19068 32176 19072
rect 32112 19012 32116 19068
rect 32116 19012 32172 19068
rect 32172 19012 32176 19068
rect 32112 19008 32176 19012
rect 32192 19068 32256 19072
rect 32192 19012 32196 19068
rect 32196 19012 32252 19068
rect 32252 19012 32256 19068
rect 32192 19008 32256 19012
rect 36952 19068 37016 19072
rect 36952 19012 36956 19068
rect 36956 19012 37012 19068
rect 37012 19012 37016 19068
rect 36952 19008 37016 19012
rect 37032 19068 37096 19072
rect 37032 19012 37036 19068
rect 37036 19012 37092 19068
rect 37092 19012 37096 19068
rect 37032 19008 37096 19012
rect 37112 19068 37176 19072
rect 37112 19012 37116 19068
rect 37116 19012 37172 19068
rect 37172 19012 37176 19068
rect 37112 19008 37176 19012
rect 37192 19068 37256 19072
rect 37192 19012 37196 19068
rect 37196 19012 37252 19068
rect 37252 19012 37256 19068
rect 37192 19008 37256 19012
rect 41952 19068 42016 19072
rect 41952 19012 41956 19068
rect 41956 19012 42012 19068
rect 42012 19012 42016 19068
rect 41952 19008 42016 19012
rect 42032 19068 42096 19072
rect 42032 19012 42036 19068
rect 42036 19012 42092 19068
rect 42092 19012 42096 19068
rect 42032 19008 42096 19012
rect 42112 19068 42176 19072
rect 42112 19012 42116 19068
rect 42116 19012 42172 19068
rect 42172 19012 42176 19068
rect 42112 19008 42176 19012
rect 42192 19068 42256 19072
rect 42192 19012 42196 19068
rect 42196 19012 42252 19068
rect 42252 19012 42256 19068
rect 42192 19008 42256 19012
rect 46952 19068 47016 19072
rect 46952 19012 46956 19068
rect 46956 19012 47012 19068
rect 47012 19012 47016 19068
rect 46952 19008 47016 19012
rect 47032 19068 47096 19072
rect 47032 19012 47036 19068
rect 47036 19012 47092 19068
rect 47092 19012 47096 19068
rect 47032 19008 47096 19012
rect 47112 19068 47176 19072
rect 47112 19012 47116 19068
rect 47116 19012 47172 19068
rect 47172 19012 47176 19068
rect 47112 19008 47176 19012
rect 47192 19068 47256 19072
rect 47192 19012 47196 19068
rect 47196 19012 47252 19068
rect 47252 19012 47256 19068
rect 47192 19008 47256 19012
rect 51952 19068 52016 19072
rect 51952 19012 51956 19068
rect 51956 19012 52012 19068
rect 52012 19012 52016 19068
rect 51952 19008 52016 19012
rect 52032 19068 52096 19072
rect 52032 19012 52036 19068
rect 52036 19012 52092 19068
rect 52092 19012 52096 19068
rect 52032 19008 52096 19012
rect 52112 19068 52176 19072
rect 52112 19012 52116 19068
rect 52116 19012 52172 19068
rect 52172 19012 52176 19068
rect 52112 19008 52176 19012
rect 52192 19068 52256 19072
rect 52192 19012 52196 19068
rect 52196 19012 52252 19068
rect 52252 19012 52256 19068
rect 52192 19008 52256 19012
rect 56952 19068 57016 19072
rect 56952 19012 56956 19068
rect 56956 19012 57012 19068
rect 57012 19012 57016 19068
rect 56952 19008 57016 19012
rect 57032 19068 57096 19072
rect 57032 19012 57036 19068
rect 57036 19012 57092 19068
rect 57092 19012 57096 19068
rect 57032 19008 57096 19012
rect 57112 19068 57176 19072
rect 57112 19012 57116 19068
rect 57116 19012 57172 19068
rect 57172 19012 57176 19068
rect 57112 19008 57176 19012
rect 57192 19068 57256 19072
rect 57192 19012 57196 19068
rect 57196 19012 57252 19068
rect 57252 19012 57256 19068
rect 57192 19008 57256 19012
rect 2612 18524 2676 18528
rect 2612 18468 2616 18524
rect 2616 18468 2672 18524
rect 2672 18468 2676 18524
rect 2612 18464 2676 18468
rect 2692 18524 2756 18528
rect 2692 18468 2696 18524
rect 2696 18468 2752 18524
rect 2752 18468 2756 18524
rect 2692 18464 2756 18468
rect 2772 18524 2836 18528
rect 2772 18468 2776 18524
rect 2776 18468 2832 18524
rect 2832 18468 2836 18524
rect 2772 18464 2836 18468
rect 2852 18524 2916 18528
rect 2852 18468 2856 18524
rect 2856 18468 2912 18524
rect 2912 18468 2916 18524
rect 2852 18464 2916 18468
rect 7612 18524 7676 18528
rect 7612 18468 7616 18524
rect 7616 18468 7672 18524
rect 7672 18468 7676 18524
rect 7612 18464 7676 18468
rect 7692 18524 7756 18528
rect 7692 18468 7696 18524
rect 7696 18468 7752 18524
rect 7752 18468 7756 18524
rect 7692 18464 7756 18468
rect 7772 18524 7836 18528
rect 7772 18468 7776 18524
rect 7776 18468 7832 18524
rect 7832 18468 7836 18524
rect 7772 18464 7836 18468
rect 7852 18524 7916 18528
rect 7852 18468 7856 18524
rect 7856 18468 7912 18524
rect 7912 18468 7916 18524
rect 7852 18464 7916 18468
rect 12612 18524 12676 18528
rect 12612 18468 12616 18524
rect 12616 18468 12672 18524
rect 12672 18468 12676 18524
rect 12612 18464 12676 18468
rect 12692 18524 12756 18528
rect 12692 18468 12696 18524
rect 12696 18468 12752 18524
rect 12752 18468 12756 18524
rect 12692 18464 12756 18468
rect 12772 18524 12836 18528
rect 12772 18468 12776 18524
rect 12776 18468 12832 18524
rect 12832 18468 12836 18524
rect 12772 18464 12836 18468
rect 12852 18524 12916 18528
rect 12852 18468 12856 18524
rect 12856 18468 12912 18524
rect 12912 18468 12916 18524
rect 12852 18464 12916 18468
rect 17612 18524 17676 18528
rect 17612 18468 17616 18524
rect 17616 18468 17672 18524
rect 17672 18468 17676 18524
rect 17612 18464 17676 18468
rect 17692 18524 17756 18528
rect 17692 18468 17696 18524
rect 17696 18468 17752 18524
rect 17752 18468 17756 18524
rect 17692 18464 17756 18468
rect 17772 18524 17836 18528
rect 17772 18468 17776 18524
rect 17776 18468 17832 18524
rect 17832 18468 17836 18524
rect 17772 18464 17836 18468
rect 17852 18524 17916 18528
rect 17852 18468 17856 18524
rect 17856 18468 17912 18524
rect 17912 18468 17916 18524
rect 17852 18464 17916 18468
rect 22612 18524 22676 18528
rect 22612 18468 22616 18524
rect 22616 18468 22672 18524
rect 22672 18468 22676 18524
rect 22612 18464 22676 18468
rect 22692 18524 22756 18528
rect 22692 18468 22696 18524
rect 22696 18468 22752 18524
rect 22752 18468 22756 18524
rect 22692 18464 22756 18468
rect 22772 18524 22836 18528
rect 22772 18468 22776 18524
rect 22776 18468 22832 18524
rect 22832 18468 22836 18524
rect 22772 18464 22836 18468
rect 22852 18524 22916 18528
rect 22852 18468 22856 18524
rect 22856 18468 22912 18524
rect 22912 18468 22916 18524
rect 22852 18464 22916 18468
rect 27612 18524 27676 18528
rect 27612 18468 27616 18524
rect 27616 18468 27672 18524
rect 27672 18468 27676 18524
rect 27612 18464 27676 18468
rect 27692 18524 27756 18528
rect 27692 18468 27696 18524
rect 27696 18468 27752 18524
rect 27752 18468 27756 18524
rect 27692 18464 27756 18468
rect 27772 18524 27836 18528
rect 27772 18468 27776 18524
rect 27776 18468 27832 18524
rect 27832 18468 27836 18524
rect 27772 18464 27836 18468
rect 27852 18524 27916 18528
rect 27852 18468 27856 18524
rect 27856 18468 27912 18524
rect 27912 18468 27916 18524
rect 27852 18464 27916 18468
rect 32612 18524 32676 18528
rect 32612 18468 32616 18524
rect 32616 18468 32672 18524
rect 32672 18468 32676 18524
rect 32612 18464 32676 18468
rect 32692 18524 32756 18528
rect 32692 18468 32696 18524
rect 32696 18468 32752 18524
rect 32752 18468 32756 18524
rect 32692 18464 32756 18468
rect 32772 18524 32836 18528
rect 32772 18468 32776 18524
rect 32776 18468 32832 18524
rect 32832 18468 32836 18524
rect 32772 18464 32836 18468
rect 32852 18524 32916 18528
rect 32852 18468 32856 18524
rect 32856 18468 32912 18524
rect 32912 18468 32916 18524
rect 32852 18464 32916 18468
rect 37612 18524 37676 18528
rect 37612 18468 37616 18524
rect 37616 18468 37672 18524
rect 37672 18468 37676 18524
rect 37612 18464 37676 18468
rect 37692 18524 37756 18528
rect 37692 18468 37696 18524
rect 37696 18468 37752 18524
rect 37752 18468 37756 18524
rect 37692 18464 37756 18468
rect 37772 18524 37836 18528
rect 37772 18468 37776 18524
rect 37776 18468 37832 18524
rect 37832 18468 37836 18524
rect 37772 18464 37836 18468
rect 37852 18524 37916 18528
rect 37852 18468 37856 18524
rect 37856 18468 37912 18524
rect 37912 18468 37916 18524
rect 37852 18464 37916 18468
rect 42612 18524 42676 18528
rect 42612 18468 42616 18524
rect 42616 18468 42672 18524
rect 42672 18468 42676 18524
rect 42612 18464 42676 18468
rect 42692 18524 42756 18528
rect 42692 18468 42696 18524
rect 42696 18468 42752 18524
rect 42752 18468 42756 18524
rect 42692 18464 42756 18468
rect 42772 18524 42836 18528
rect 42772 18468 42776 18524
rect 42776 18468 42832 18524
rect 42832 18468 42836 18524
rect 42772 18464 42836 18468
rect 42852 18524 42916 18528
rect 42852 18468 42856 18524
rect 42856 18468 42912 18524
rect 42912 18468 42916 18524
rect 42852 18464 42916 18468
rect 47612 18524 47676 18528
rect 47612 18468 47616 18524
rect 47616 18468 47672 18524
rect 47672 18468 47676 18524
rect 47612 18464 47676 18468
rect 47692 18524 47756 18528
rect 47692 18468 47696 18524
rect 47696 18468 47752 18524
rect 47752 18468 47756 18524
rect 47692 18464 47756 18468
rect 47772 18524 47836 18528
rect 47772 18468 47776 18524
rect 47776 18468 47832 18524
rect 47832 18468 47836 18524
rect 47772 18464 47836 18468
rect 47852 18524 47916 18528
rect 47852 18468 47856 18524
rect 47856 18468 47912 18524
rect 47912 18468 47916 18524
rect 47852 18464 47916 18468
rect 52612 18524 52676 18528
rect 52612 18468 52616 18524
rect 52616 18468 52672 18524
rect 52672 18468 52676 18524
rect 52612 18464 52676 18468
rect 52692 18524 52756 18528
rect 52692 18468 52696 18524
rect 52696 18468 52752 18524
rect 52752 18468 52756 18524
rect 52692 18464 52756 18468
rect 52772 18524 52836 18528
rect 52772 18468 52776 18524
rect 52776 18468 52832 18524
rect 52832 18468 52836 18524
rect 52772 18464 52836 18468
rect 52852 18524 52916 18528
rect 52852 18468 52856 18524
rect 52856 18468 52912 18524
rect 52912 18468 52916 18524
rect 52852 18464 52916 18468
rect 57612 18524 57676 18528
rect 57612 18468 57616 18524
rect 57616 18468 57672 18524
rect 57672 18468 57676 18524
rect 57612 18464 57676 18468
rect 57692 18524 57756 18528
rect 57692 18468 57696 18524
rect 57696 18468 57752 18524
rect 57752 18468 57756 18524
rect 57692 18464 57756 18468
rect 57772 18524 57836 18528
rect 57772 18468 57776 18524
rect 57776 18468 57832 18524
rect 57832 18468 57836 18524
rect 57772 18464 57836 18468
rect 57852 18524 57916 18528
rect 57852 18468 57856 18524
rect 57856 18468 57912 18524
rect 57912 18468 57916 18524
rect 57852 18464 57916 18468
rect 1952 17980 2016 17984
rect 1952 17924 1956 17980
rect 1956 17924 2012 17980
rect 2012 17924 2016 17980
rect 1952 17920 2016 17924
rect 2032 17980 2096 17984
rect 2032 17924 2036 17980
rect 2036 17924 2092 17980
rect 2092 17924 2096 17980
rect 2032 17920 2096 17924
rect 2112 17980 2176 17984
rect 2112 17924 2116 17980
rect 2116 17924 2172 17980
rect 2172 17924 2176 17980
rect 2112 17920 2176 17924
rect 2192 17980 2256 17984
rect 2192 17924 2196 17980
rect 2196 17924 2252 17980
rect 2252 17924 2256 17980
rect 2192 17920 2256 17924
rect 6952 17980 7016 17984
rect 6952 17924 6956 17980
rect 6956 17924 7012 17980
rect 7012 17924 7016 17980
rect 6952 17920 7016 17924
rect 7032 17980 7096 17984
rect 7032 17924 7036 17980
rect 7036 17924 7092 17980
rect 7092 17924 7096 17980
rect 7032 17920 7096 17924
rect 7112 17980 7176 17984
rect 7112 17924 7116 17980
rect 7116 17924 7172 17980
rect 7172 17924 7176 17980
rect 7112 17920 7176 17924
rect 7192 17980 7256 17984
rect 7192 17924 7196 17980
rect 7196 17924 7252 17980
rect 7252 17924 7256 17980
rect 7192 17920 7256 17924
rect 11952 17980 12016 17984
rect 11952 17924 11956 17980
rect 11956 17924 12012 17980
rect 12012 17924 12016 17980
rect 11952 17920 12016 17924
rect 12032 17980 12096 17984
rect 12032 17924 12036 17980
rect 12036 17924 12092 17980
rect 12092 17924 12096 17980
rect 12032 17920 12096 17924
rect 12112 17980 12176 17984
rect 12112 17924 12116 17980
rect 12116 17924 12172 17980
rect 12172 17924 12176 17980
rect 12112 17920 12176 17924
rect 12192 17980 12256 17984
rect 12192 17924 12196 17980
rect 12196 17924 12252 17980
rect 12252 17924 12256 17980
rect 12192 17920 12256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 21952 17980 22016 17984
rect 21952 17924 21956 17980
rect 21956 17924 22012 17980
rect 22012 17924 22016 17980
rect 21952 17920 22016 17924
rect 22032 17980 22096 17984
rect 22032 17924 22036 17980
rect 22036 17924 22092 17980
rect 22092 17924 22096 17980
rect 22032 17920 22096 17924
rect 22112 17980 22176 17984
rect 22112 17924 22116 17980
rect 22116 17924 22172 17980
rect 22172 17924 22176 17980
rect 22112 17920 22176 17924
rect 22192 17980 22256 17984
rect 22192 17924 22196 17980
rect 22196 17924 22252 17980
rect 22252 17924 22256 17980
rect 22192 17920 22256 17924
rect 26952 17980 27016 17984
rect 26952 17924 26956 17980
rect 26956 17924 27012 17980
rect 27012 17924 27016 17980
rect 26952 17920 27016 17924
rect 27032 17980 27096 17984
rect 27032 17924 27036 17980
rect 27036 17924 27092 17980
rect 27092 17924 27096 17980
rect 27032 17920 27096 17924
rect 27112 17980 27176 17984
rect 27112 17924 27116 17980
rect 27116 17924 27172 17980
rect 27172 17924 27176 17980
rect 27112 17920 27176 17924
rect 27192 17980 27256 17984
rect 27192 17924 27196 17980
rect 27196 17924 27252 17980
rect 27252 17924 27256 17980
rect 27192 17920 27256 17924
rect 31952 17980 32016 17984
rect 31952 17924 31956 17980
rect 31956 17924 32012 17980
rect 32012 17924 32016 17980
rect 31952 17920 32016 17924
rect 32032 17980 32096 17984
rect 32032 17924 32036 17980
rect 32036 17924 32092 17980
rect 32092 17924 32096 17980
rect 32032 17920 32096 17924
rect 32112 17980 32176 17984
rect 32112 17924 32116 17980
rect 32116 17924 32172 17980
rect 32172 17924 32176 17980
rect 32112 17920 32176 17924
rect 32192 17980 32256 17984
rect 32192 17924 32196 17980
rect 32196 17924 32252 17980
rect 32252 17924 32256 17980
rect 32192 17920 32256 17924
rect 36952 17980 37016 17984
rect 36952 17924 36956 17980
rect 36956 17924 37012 17980
rect 37012 17924 37016 17980
rect 36952 17920 37016 17924
rect 37032 17980 37096 17984
rect 37032 17924 37036 17980
rect 37036 17924 37092 17980
rect 37092 17924 37096 17980
rect 37032 17920 37096 17924
rect 37112 17980 37176 17984
rect 37112 17924 37116 17980
rect 37116 17924 37172 17980
rect 37172 17924 37176 17980
rect 37112 17920 37176 17924
rect 37192 17980 37256 17984
rect 37192 17924 37196 17980
rect 37196 17924 37252 17980
rect 37252 17924 37256 17980
rect 37192 17920 37256 17924
rect 41952 17980 42016 17984
rect 41952 17924 41956 17980
rect 41956 17924 42012 17980
rect 42012 17924 42016 17980
rect 41952 17920 42016 17924
rect 42032 17980 42096 17984
rect 42032 17924 42036 17980
rect 42036 17924 42092 17980
rect 42092 17924 42096 17980
rect 42032 17920 42096 17924
rect 42112 17980 42176 17984
rect 42112 17924 42116 17980
rect 42116 17924 42172 17980
rect 42172 17924 42176 17980
rect 42112 17920 42176 17924
rect 42192 17980 42256 17984
rect 42192 17924 42196 17980
rect 42196 17924 42252 17980
rect 42252 17924 42256 17980
rect 42192 17920 42256 17924
rect 46952 17980 47016 17984
rect 46952 17924 46956 17980
rect 46956 17924 47012 17980
rect 47012 17924 47016 17980
rect 46952 17920 47016 17924
rect 47032 17980 47096 17984
rect 47032 17924 47036 17980
rect 47036 17924 47092 17980
rect 47092 17924 47096 17980
rect 47032 17920 47096 17924
rect 47112 17980 47176 17984
rect 47112 17924 47116 17980
rect 47116 17924 47172 17980
rect 47172 17924 47176 17980
rect 47112 17920 47176 17924
rect 47192 17980 47256 17984
rect 47192 17924 47196 17980
rect 47196 17924 47252 17980
rect 47252 17924 47256 17980
rect 47192 17920 47256 17924
rect 51952 17980 52016 17984
rect 51952 17924 51956 17980
rect 51956 17924 52012 17980
rect 52012 17924 52016 17980
rect 51952 17920 52016 17924
rect 52032 17980 52096 17984
rect 52032 17924 52036 17980
rect 52036 17924 52092 17980
rect 52092 17924 52096 17980
rect 52032 17920 52096 17924
rect 52112 17980 52176 17984
rect 52112 17924 52116 17980
rect 52116 17924 52172 17980
rect 52172 17924 52176 17980
rect 52112 17920 52176 17924
rect 52192 17980 52256 17984
rect 52192 17924 52196 17980
rect 52196 17924 52252 17980
rect 52252 17924 52256 17980
rect 52192 17920 52256 17924
rect 56952 17980 57016 17984
rect 56952 17924 56956 17980
rect 56956 17924 57012 17980
rect 57012 17924 57016 17980
rect 56952 17920 57016 17924
rect 57032 17980 57096 17984
rect 57032 17924 57036 17980
rect 57036 17924 57092 17980
rect 57092 17924 57096 17980
rect 57032 17920 57096 17924
rect 57112 17980 57176 17984
rect 57112 17924 57116 17980
rect 57116 17924 57172 17980
rect 57172 17924 57176 17980
rect 57112 17920 57176 17924
rect 57192 17980 57256 17984
rect 57192 17924 57196 17980
rect 57196 17924 57252 17980
rect 57252 17924 57256 17980
rect 57192 17920 57256 17924
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 22612 17436 22676 17440
rect 22612 17380 22616 17436
rect 22616 17380 22672 17436
rect 22672 17380 22676 17436
rect 22612 17376 22676 17380
rect 22692 17436 22756 17440
rect 22692 17380 22696 17436
rect 22696 17380 22752 17436
rect 22752 17380 22756 17436
rect 22692 17376 22756 17380
rect 22772 17436 22836 17440
rect 22772 17380 22776 17436
rect 22776 17380 22832 17436
rect 22832 17380 22836 17436
rect 22772 17376 22836 17380
rect 22852 17436 22916 17440
rect 22852 17380 22856 17436
rect 22856 17380 22912 17436
rect 22912 17380 22916 17436
rect 22852 17376 22916 17380
rect 27612 17436 27676 17440
rect 27612 17380 27616 17436
rect 27616 17380 27672 17436
rect 27672 17380 27676 17436
rect 27612 17376 27676 17380
rect 27692 17436 27756 17440
rect 27692 17380 27696 17436
rect 27696 17380 27752 17436
rect 27752 17380 27756 17436
rect 27692 17376 27756 17380
rect 27772 17436 27836 17440
rect 27772 17380 27776 17436
rect 27776 17380 27832 17436
rect 27832 17380 27836 17436
rect 27772 17376 27836 17380
rect 27852 17436 27916 17440
rect 27852 17380 27856 17436
rect 27856 17380 27912 17436
rect 27912 17380 27916 17436
rect 27852 17376 27916 17380
rect 32612 17436 32676 17440
rect 32612 17380 32616 17436
rect 32616 17380 32672 17436
rect 32672 17380 32676 17436
rect 32612 17376 32676 17380
rect 32692 17436 32756 17440
rect 32692 17380 32696 17436
rect 32696 17380 32752 17436
rect 32752 17380 32756 17436
rect 32692 17376 32756 17380
rect 32772 17436 32836 17440
rect 32772 17380 32776 17436
rect 32776 17380 32832 17436
rect 32832 17380 32836 17436
rect 32772 17376 32836 17380
rect 32852 17436 32916 17440
rect 32852 17380 32856 17436
rect 32856 17380 32912 17436
rect 32912 17380 32916 17436
rect 32852 17376 32916 17380
rect 37612 17436 37676 17440
rect 37612 17380 37616 17436
rect 37616 17380 37672 17436
rect 37672 17380 37676 17436
rect 37612 17376 37676 17380
rect 37692 17436 37756 17440
rect 37692 17380 37696 17436
rect 37696 17380 37752 17436
rect 37752 17380 37756 17436
rect 37692 17376 37756 17380
rect 37772 17436 37836 17440
rect 37772 17380 37776 17436
rect 37776 17380 37832 17436
rect 37832 17380 37836 17436
rect 37772 17376 37836 17380
rect 37852 17436 37916 17440
rect 37852 17380 37856 17436
rect 37856 17380 37912 17436
rect 37912 17380 37916 17436
rect 37852 17376 37916 17380
rect 42612 17436 42676 17440
rect 42612 17380 42616 17436
rect 42616 17380 42672 17436
rect 42672 17380 42676 17436
rect 42612 17376 42676 17380
rect 42692 17436 42756 17440
rect 42692 17380 42696 17436
rect 42696 17380 42752 17436
rect 42752 17380 42756 17436
rect 42692 17376 42756 17380
rect 42772 17436 42836 17440
rect 42772 17380 42776 17436
rect 42776 17380 42832 17436
rect 42832 17380 42836 17436
rect 42772 17376 42836 17380
rect 42852 17436 42916 17440
rect 42852 17380 42856 17436
rect 42856 17380 42912 17436
rect 42912 17380 42916 17436
rect 42852 17376 42916 17380
rect 47612 17436 47676 17440
rect 47612 17380 47616 17436
rect 47616 17380 47672 17436
rect 47672 17380 47676 17436
rect 47612 17376 47676 17380
rect 47692 17436 47756 17440
rect 47692 17380 47696 17436
rect 47696 17380 47752 17436
rect 47752 17380 47756 17436
rect 47692 17376 47756 17380
rect 47772 17436 47836 17440
rect 47772 17380 47776 17436
rect 47776 17380 47832 17436
rect 47832 17380 47836 17436
rect 47772 17376 47836 17380
rect 47852 17436 47916 17440
rect 47852 17380 47856 17436
rect 47856 17380 47912 17436
rect 47912 17380 47916 17436
rect 47852 17376 47916 17380
rect 52612 17436 52676 17440
rect 52612 17380 52616 17436
rect 52616 17380 52672 17436
rect 52672 17380 52676 17436
rect 52612 17376 52676 17380
rect 52692 17436 52756 17440
rect 52692 17380 52696 17436
rect 52696 17380 52752 17436
rect 52752 17380 52756 17436
rect 52692 17376 52756 17380
rect 52772 17436 52836 17440
rect 52772 17380 52776 17436
rect 52776 17380 52832 17436
rect 52832 17380 52836 17436
rect 52772 17376 52836 17380
rect 52852 17436 52916 17440
rect 52852 17380 52856 17436
rect 52856 17380 52912 17436
rect 52912 17380 52916 17436
rect 52852 17376 52916 17380
rect 57612 17436 57676 17440
rect 57612 17380 57616 17436
rect 57616 17380 57672 17436
rect 57672 17380 57676 17436
rect 57612 17376 57676 17380
rect 57692 17436 57756 17440
rect 57692 17380 57696 17436
rect 57696 17380 57752 17436
rect 57752 17380 57756 17436
rect 57692 17376 57756 17380
rect 57772 17436 57836 17440
rect 57772 17380 57776 17436
rect 57776 17380 57832 17436
rect 57832 17380 57836 17436
rect 57772 17376 57836 17380
rect 57852 17436 57916 17440
rect 57852 17380 57856 17436
rect 57856 17380 57912 17436
rect 57912 17380 57916 17436
rect 57852 17376 57916 17380
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 21952 16892 22016 16896
rect 21952 16836 21956 16892
rect 21956 16836 22012 16892
rect 22012 16836 22016 16892
rect 21952 16832 22016 16836
rect 22032 16892 22096 16896
rect 22032 16836 22036 16892
rect 22036 16836 22092 16892
rect 22092 16836 22096 16892
rect 22032 16832 22096 16836
rect 22112 16892 22176 16896
rect 22112 16836 22116 16892
rect 22116 16836 22172 16892
rect 22172 16836 22176 16892
rect 22112 16832 22176 16836
rect 22192 16892 22256 16896
rect 22192 16836 22196 16892
rect 22196 16836 22252 16892
rect 22252 16836 22256 16892
rect 22192 16832 22256 16836
rect 26952 16892 27016 16896
rect 26952 16836 26956 16892
rect 26956 16836 27012 16892
rect 27012 16836 27016 16892
rect 26952 16832 27016 16836
rect 27032 16892 27096 16896
rect 27032 16836 27036 16892
rect 27036 16836 27092 16892
rect 27092 16836 27096 16892
rect 27032 16832 27096 16836
rect 27112 16892 27176 16896
rect 27112 16836 27116 16892
rect 27116 16836 27172 16892
rect 27172 16836 27176 16892
rect 27112 16832 27176 16836
rect 27192 16892 27256 16896
rect 27192 16836 27196 16892
rect 27196 16836 27252 16892
rect 27252 16836 27256 16892
rect 27192 16832 27256 16836
rect 31952 16892 32016 16896
rect 31952 16836 31956 16892
rect 31956 16836 32012 16892
rect 32012 16836 32016 16892
rect 31952 16832 32016 16836
rect 32032 16892 32096 16896
rect 32032 16836 32036 16892
rect 32036 16836 32092 16892
rect 32092 16836 32096 16892
rect 32032 16832 32096 16836
rect 32112 16892 32176 16896
rect 32112 16836 32116 16892
rect 32116 16836 32172 16892
rect 32172 16836 32176 16892
rect 32112 16832 32176 16836
rect 32192 16892 32256 16896
rect 32192 16836 32196 16892
rect 32196 16836 32252 16892
rect 32252 16836 32256 16892
rect 32192 16832 32256 16836
rect 36952 16892 37016 16896
rect 36952 16836 36956 16892
rect 36956 16836 37012 16892
rect 37012 16836 37016 16892
rect 36952 16832 37016 16836
rect 37032 16892 37096 16896
rect 37032 16836 37036 16892
rect 37036 16836 37092 16892
rect 37092 16836 37096 16892
rect 37032 16832 37096 16836
rect 37112 16892 37176 16896
rect 37112 16836 37116 16892
rect 37116 16836 37172 16892
rect 37172 16836 37176 16892
rect 37112 16832 37176 16836
rect 37192 16892 37256 16896
rect 37192 16836 37196 16892
rect 37196 16836 37252 16892
rect 37252 16836 37256 16892
rect 37192 16832 37256 16836
rect 41952 16892 42016 16896
rect 41952 16836 41956 16892
rect 41956 16836 42012 16892
rect 42012 16836 42016 16892
rect 41952 16832 42016 16836
rect 42032 16892 42096 16896
rect 42032 16836 42036 16892
rect 42036 16836 42092 16892
rect 42092 16836 42096 16892
rect 42032 16832 42096 16836
rect 42112 16892 42176 16896
rect 42112 16836 42116 16892
rect 42116 16836 42172 16892
rect 42172 16836 42176 16892
rect 42112 16832 42176 16836
rect 42192 16892 42256 16896
rect 42192 16836 42196 16892
rect 42196 16836 42252 16892
rect 42252 16836 42256 16892
rect 42192 16832 42256 16836
rect 46952 16892 47016 16896
rect 46952 16836 46956 16892
rect 46956 16836 47012 16892
rect 47012 16836 47016 16892
rect 46952 16832 47016 16836
rect 47032 16892 47096 16896
rect 47032 16836 47036 16892
rect 47036 16836 47092 16892
rect 47092 16836 47096 16892
rect 47032 16832 47096 16836
rect 47112 16892 47176 16896
rect 47112 16836 47116 16892
rect 47116 16836 47172 16892
rect 47172 16836 47176 16892
rect 47112 16832 47176 16836
rect 47192 16892 47256 16896
rect 47192 16836 47196 16892
rect 47196 16836 47252 16892
rect 47252 16836 47256 16892
rect 47192 16832 47256 16836
rect 51952 16892 52016 16896
rect 51952 16836 51956 16892
rect 51956 16836 52012 16892
rect 52012 16836 52016 16892
rect 51952 16832 52016 16836
rect 52032 16892 52096 16896
rect 52032 16836 52036 16892
rect 52036 16836 52092 16892
rect 52092 16836 52096 16892
rect 52032 16832 52096 16836
rect 52112 16892 52176 16896
rect 52112 16836 52116 16892
rect 52116 16836 52172 16892
rect 52172 16836 52176 16892
rect 52112 16832 52176 16836
rect 52192 16892 52256 16896
rect 52192 16836 52196 16892
rect 52196 16836 52252 16892
rect 52252 16836 52256 16892
rect 52192 16832 52256 16836
rect 56952 16892 57016 16896
rect 56952 16836 56956 16892
rect 56956 16836 57012 16892
rect 57012 16836 57016 16892
rect 56952 16832 57016 16836
rect 57032 16892 57096 16896
rect 57032 16836 57036 16892
rect 57036 16836 57092 16892
rect 57092 16836 57096 16892
rect 57032 16832 57096 16836
rect 57112 16892 57176 16896
rect 57112 16836 57116 16892
rect 57116 16836 57172 16892
rect 57172 16836 57176 16892
rect 57112 16832 57176 16836
rect 57192 16892 57256 16896
rect 57192 16836 57196 16892
rect 57196 16836 57252 16892
rect 57252 16836 57256 16892
rect 57192 16832 57256 16836
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 22612 16348 22676 16352
rect 22612 16292 22616 16348
rect 22616 16292 22672 16348
rect 22672 16292 22676 16348
rect 22612 16288 22676 16292
rect 22692 16348 22756 16352
rect 22692 16292 22696 16348
rect 22696 16292 22752 16348
rect 22752 16292 22756 16348
rect 22692 16288 22756 16292
rect 22772 16348 22836 16352
rect 22772 16292 22776 16348
rect 22776 16292 22832 16348
rect 22832 16292 22836 16348
rect 22772 16288 22836 16292
rect 22852 16348 22916 16352
rect 22852 16292 22856 16348
rect 22856 16292 22912 16348
rect 22912 16292 22916 16348
rect 22852 16288 22916 16292
rect 27612 16348 27676 16352
rect 27612 16292 27616 16348
rect 27616 16292 27672 16348
rect 27672 16292 27676 16348
rect 27612 16288 27676 16292
rect 27692 16348 27756 16352
rect 27692 16292 27696 16348
rect 27696 16292 27752 16348
rect 27752 16292 27756 16348
rect 27692 16288 27756 16292
rect 27772 16348 27836 16352
rect 27772 16292 27776 16348
rect 27776 16292 27832 16348
rect 27832 16292 27836 16348
rect 27772 16288 27836 16292
rect 27852 16348 27916 16352
rect 27852 16292 27856 16348
rect 27856 16292 27912 16348
rect 27912 16292 27916 16348
rect 27852 16288 27916 16292
rect 32612 16348 32676 16352
rect 32612 16292 32616 16348
rect 32616 16292 32672 16348
rect 32672 16292 32676 16348
rect 32612 16288 32676 16292
rect 32692 16348 32756 16352
rect 32692 16292 32696 16348
rect 32696 16292 32752 16348
rect 32752 16292 32756 16348
rect 32692 16288 32756 16292
rect 32772 16348 32836 16352
rect 32772 16292 32776 16348
rect 32776 16292 32832 16348
rect 32832 16292 32836 16348
rect 32772 16288 32836 16292
rect 32852 16348 32916 16352
rect 32852 16292 32856 16348
rect 32856 16292 32912 16348
rect 32912 16292 32916 16348
rect 32852 16288 32916 16292
rect 37612 16348 37676 16352
rect 37612 16292 37616 16348
rect 37616 16292 37672 16348
rect 37672 16292 37676 16348
rect 37612 16288 37676 16292
rect 37692 16348 37756 16352
rect 37692 16292 37696 16348
rect 37696 16292 37752 16348
rect 37752 16292 37756 16348
rect 37692 16288 37756 16292
rect 37772 16348 37836 16352
rect 37772 16292 37776 16348
rect 37776 16292 37832 16348
rect 37832 16292 37836 16348
rect 37772 16288 37836 16292
rect 37852 16348 37916 16352
rect 37852 16292 37856 16348
rect 37856 16292 37912 16348
rect 37912 16292 37916 16348
rect 37852 16288 37916 16292
rect 42612 16348 42676 16352
rect 42612 16292 42616 16348
rect 42616 16292 42672 16348
rect 42672 16292 42676 16348
rect 42612 16288 42676 16292
rect 42692 16348 42756 16352
rect 42692 16292 42696 16348
rect 42696 16292 42752 16348
rect 42752 16292 42756 16348
rect 42692 16288 42756 16292
rect 42772 16348 42836 16352
rect 42772 16292 42776 16348
rect 42776 16292 42832 16348
rect 42832 16292 42836 16348
rect 42772 16288 42836 16292
rect 42852 16348 42916 16352
rect 42852 16292 42856 16348
rect 42856 16292 42912 16348
rect 42912 16292 42916 16348
rect 42852 16288 42916 16292
rect 47612 16348 47676 16352
rect 47612 16292 47616 16348
rect 47616 16292 47672 16348
rect 47672 16292 47676 16348
rect 47612 16288 47676 16292
rect 47692 16348 47756 16352
rect 47692 16292 47696 16348
rect 47696 16292 47752 16348
rect 47752 16292 47756 16348
rect 47692 16288 47756 16292
rect 47772 16348 47836 16352
rect 47772 16292 47776 16348
rect 47776 16292 47832 16348
rect 47832 16292 47836 16348
rect 47772 16288 47836 16292
rect 47852 16348 47916 16352
rect 47852 16292 47856 16348
rect 47856 16292 47912 16348
rect 47912 16292 47916 16348
rect 47852 16288 47916 16292
rect 52612 16348 52676 16352
rect 52612 16292 52616 16348
rect 52616 16292 52672 16348
rect 52672 16292 52676 16348
rect 52612 16288 52676 16292
rect 52692 16348 52756 16352
rect 52692 16292 52696 16348
rect 52696 16292 52752 16348
rect 52752 16292 52756 16348
rect 52692 16288 52756 16292
rect 52772 16348 52836 16352
rect 52772 16292 52776 16348
rect 52776 16292 52832 16348
rect 52832 16292 52836 16348
rect 52772 16288 52836 16292
rect 52852 16348 52916 16352
rect 52852 16292 52856 16348
rect 52856 16292 52912 16348
rect 52912 16292 52916 16348
rect 52852 16288 52916 16292
rect 57612 16348 57676 16352
rect 57612 16292 57616 16348
rect 57616 16292 57672 16348
rect 57672 16292 57676 16348
rect 57612 16288 57676 16292
rect 57692 16348 57756 16352
rect 57692 16292 57696 16348
rect 57696 16292 57752 16348
rect 57752 16292 57756 16348
rect 57692 16288 57756 16292
rect 57772 16348 57836 16352
rect 57772 16292 57776 16348
rect 57776 16292 57832 16348
rect 57832 16292 57836 16348
rect 57772 16288 57836 16292
rect 57852 16348 57916 16352
rect 57852 16292 57856 16348
rect 57856 16292 57912 16348
rect 57912 16292 57916 16348
rect 57852 16288 57916 16292
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 21952 15804 22016 15808
rect 21952 15748 21956 15804
rect 21956 15748 22012 15804
rect 22012 15748 22016 15804
rect 21952 15744 22016 15748
rect 22032 15804 22096 15808
rect 22032 15748 22036 15804
rect 22036 15748 22092 15804
rect 22092 15748 22096 15804
rect 22032 15744 22096 15748
rect 22112 15804 22176 15808
rect 22112 15748 22116 15804
rect 22116 15748 22172 15804
rect 22172 15748 22176 15804
rect 22112 15744 22176 15748
rect 22192 15804 22256 15808
rect 22192 15748 22196 15804
rect 22196 15748 22252 15804
rect 22252 15748 22256 15804
rect 22192 15744 22256 15748
rect 26952 15804 27016 15808
rect 26952 15748 26956 15804
rect 26956 15748 27012 15804
rect 27012 15748 27016 15804
rect 26952 15744 27016 15748
rect 27032 15804 27096 15808
rect 27032 15748 27036 15804
rect 27036 15748 27092 15804
rect 27092 15748 27096 15804
rect 27032 15744 27096 15748
rect 27112 15804 27176 15808
rect 27112 15748 27116 15804
rect 27116 15748 27172 15804
rect 27172 15748 27176 15804
rect 27112 15744 27176 15748
rect 27192 15804 27256 15808
rect 27192 15748 27196 15804
rect 27196 15748 27252 15804
rect 27252 15748 27256 15804
rect 27192 15744 27256 15748
rect 31952 15804 32016 15808
rect 31952 15748 31956 15804
rect 31956 15748 32012 15804
rect 32012 15748 32016 15804
rect 31952 15744 32016 15748
rect 32032 15804 32096 15808
rect 32032 15748 32036 15804
rect 32036 15748 32092 15804
rect 32092 15748 32096 15804
rect 32032 15744 32096 15748
rect 32112 15804 32176 15808
rect 32112 15748 32116 15804
rect 32116 15748 32172 15804
rect 32172 15748 32176 15804
rect 32112 15744 32176 15748
rect 32192 15804 32256 15808
rect 32192 15748 32196 15804
rect 32196 15748 32252 15804
rect 32252 15748 32256 15804
rect 32192 15744 32256 15748
rect 36952 15804 37016 15808
rect 36952 15748 36956 15804
rect 36956 15748 37012 15804
rect 37012 15748 37016 15804
rect 36952 15744 37016 15748
rect 37032 15804 37096 15808
rect 37032 15748 37036 15804
rect 37036 15748 37092 15804
rect 37092 15748 37096 15804
rect 37032 15744 37096 15748
rect 37112 15804 37176 15808
rect 37112 15748 37116 15804
rect 37116 15748 37172 15804
rect 37172 15748 37176 15804
rect 37112 15744 37176 15748
rect 37192 15804 37256 15808
rect 37192 15748 37196 15804
rect 37196 15748 37252 15804
rect 37252 15748 37256 15804
rect 37192 15744 37256 15748
rect 41952 15804 42016 15808
rect 41952 15748 41956 15804
rect 41956 15748 42012 15804
rect 42012 15748 42016 15804
rect 41952 15744 42016 15748
rect 42032 15804 42096 15808
rect 42032 15748 42036 15804
rect 42036 15748 42092 15804
rect 42092 15748 42096 15804
rect 42032 15744 42096 15748
rect 42112 15804 42176 15808
rect 42112 15748 42116 15804
rect 42116 15748 42172 15804
rect 42172 15748 42176 15804
rect 42112 15744 42176 15748
rect 42192 15804 42256 15808
rect 42192 15748 42196 15804
rect 42196 15748 42252 15804
rect 42252 15748 42256 15804
rect 42192 15744 42256 15748
rect 46952 15804 47016 15808
rect 46952 15748 46956 15804
rect 46956 15748 47012 15804
rect 47012 15748 47016 15804
rect 46952 15744 47016 15748
rect 47032 15804 47096 15808
rect 47032 15748 47036 15804
rect 47036 15748 47092 15804
rect 47092 15748 47096 15804
rect 47032 15744 47096 15748
rect 47112 15804 47176 15808
rect 47112 15748 47116 15804
rect 47116 15748 47172 15804
rect 47172 15748 47176 15804
rect 47112 15744 47176 15748
rect 47192 15804 47256 15808
rect 47192 15748 47196 15804
rect 47196 15748 47252 15804
rect 47252 15748 47256 15804
rect 47192 15744 47256 15748
rect 51952 15804 52016 15808
rect 51952 15748 51956 15804
rect 51956 15748 52012 15804
rect 52012 15748 52016 15804
rect 51952 15744 52016 15748
rect 52032 15804 52096 15808
rect 52032 15748 52036 15804
rect 52036 15748 52092 15804
rect 52092 15748 52096 15804
rect 52032 15744 52096 15748
rect 52112 15804 52176 15808
rect 52112 15748 52116 15804
rect 52116 15748 52172 15804
rect 52172 15748 52176 15804
rect 52112 15744 52176 15748
rect 52192 15804 52256 15808
rect 52192 15748 52196 15804
rect 52196 15748 52252 15804
rect 52252 15748 52256 15804
rect 52192 15744 52256 15748
rect 56952 15804 57016 15808
rect 56952 15748 56956 15804
rect 56956 15748 57012 15804
rect 57012 15748 57016 15804
rect 56952 15744 57016 15748
rect 57032 15804 57096 15808
rect 57032 15748 57036 15804
rect 57036 15748 57092 15804
rect 57092 15748 57096 15804
rect 57032 15744 57096 15748
rect 57112 15804 57176 15808
rect 57112 15748 57116 15804
rect 57116 15748 57172 15804
rect 57172 15748 57176 15804
rect 57112 15744 57176 15748
rect 57192 15804 57256 15808
rect 57192 15748 57196 15804
rect 57196 15748 57252 15804
rect 57252 15748 57256 15804
rect 57192 15744 57256 15748
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 22612 15260 22676 15264
rect 22612 15204 22616 15260
rect 22616 15204 22672 15260
rect 22672 15204 22676 15260
rect 22612 15200 22676 15204
rect 22692 15260 22756 15264
rect 22692 15204 22696 15260
rect 22696 15204 22752 15260
rect 22752 15204 22756 15260
rect 22692 15200 22756 15204
rect 22772 15260 22836 15264
rect 22772 15204 22776 15260
rect 22776 15204 22832 15260
rect 22832 15204 22836 15260
rect 22772 15200 22836 15204
rect 22852 15260 22916 15264
rect 22852 15204 22856 15260
rect 22856 15204 22912 15260
rect 22912 15204 22916 15260
rect 22852 15200 22916 15204
rect 27612 15260 27676 15264
rect 27612 15204 27616 15260
rect 27616 15204 27672 15260
rect 27672 15204 27676 15260
rect 27612 15200 27676 15204
rect 27692 15260 27756 15264
rect 27692 15204 27696 15260
rect 27696 15204 27752 15260
rect 27752 15204 27756 15260
rect 27692 15200 27756 15204
rect 27772 15260 27836 15264
rect 27772 15204 27776 15260
rect 27776 15204 27832 15260
rect 27832 15204 27836 15260
rect 27772 15200 27836 15204
rect 27852 15260 27916 15264
rect 27852 15204 27856 15260
rect 27856 15204 27912 15260
rect 27912 15204 27916 15260
rect 27852 15200 27916 15204
rect 32612 15260 32676 15264
rect 32612 15204 32616 15260
rect 32616 15204 32672 15260
rect 32672 15204 32676 15260
rect 32612 15200 32676 15204
rect 32692 15260 32756 15264
rect 32692 15204 32696 15260
rect 32696 15204 32752 15260
rect 32752 15204 32756 15260
rect 32692 15200 32756 15204
rect 32772 15260 32836 15264
rect 32772 15204 32776 15260
rect 32776 15204 32832 15260
rect 32832 15204 32836 15260
rect 32772 15200 32836 15204
rect 32852 15260 32916 15264
rect 32852 15204 32856 15260
rect 32856 15204 32912 15260
rect 32912 15204 32916 15260
rect 32852 15200 32916 15204
rect 37612 15260 37676 15264
rect 37612 15204 37616 15260
rect 37616 15204 37672 15260
rect 37672 15204 37676 15260
rect 37612 15200 37676 15204
rect 37692 15260 37756 15264
rect 37692 15204 37696 15260
rect 37696 15204 37752 15260
rect 37752 15204 37756 15260
rect 37692 15200 37756 15204
rect 37772 15260 37836 15264
rect 37772 15204 37776 15260
rect 37776 15204 37832 15260
rect 37832 15204 37836 15260
rect 37772 15200 37836 15204
rect 37852 15260 37916 15264
rect 37852 15204 37856 15260
rect 37856 15204 37912 15260
rect 37912 15204 37916 15260
rect 37852 15200 37916 15204
rect 42612 15260 42676 15264
rect 42612 15204 42616 15260
rect 42616 15204 42672 15260
rect 42672 15204 42676 15260
rect 42612 15200 42676 15204
rect 42692 15260 42756 15264
rect 42692 15204 42696 15260
rect 42696 15204 42752 15260
rect 42752 15204 42756 15260
rect 42692 15200 42756 15204
rect 42772 15260 42836 15264
rect 42772 15204 42776 15260
rect 42776 15204 42832 15260
rect 42832 15204 42836 15260
rect 42772 15200 42836 15204
rect 42852 15260 42916 15264
rect 42852 15204 42856 15260
rect 42856 15204 42912 15260
rect 42912 15204 42916 15260
rect 42852 15200 42916 15204
rect 47612 15260 47676 15264
rect 47612 15204 47616 15260
rect 47616 15204 47672 15260
rect 47672 15204 47676 15260
rect 47612 15200 47676 15204
rect 47692 15260 47756 15264
rect 47692 15204 47696 15260
rect 47696 15204 47752 15260
rect 47752 15204 47756 15260
rect 47692 15200 47756 15204
rect 47772 15260 47836 15264
rect 47772 15204 47776 15260
rect 47776 15204 47832 15260
rect 47832 15204 47836 15260
rect 47772 15200 47836 15204
rect 47852 15260 47916 15264
rect 47852 15204 47856 15260
rect 47856 15204 47912 15260
rect 47912 15204 47916 15260
rect 47852 15200 47916 15204
rect 52612 15260 52676 15264
rect 52612 15204 52616 15260
rect 52616 15204 52672 15260
rect 52672 15204 52676 15260
rect 52612 15200 52676 15204
rect 52692 15260 52756 15264
rect 52692 15204 52696 15260
rect 52696 15204 52752 15260
rect 52752 15204 52756 15260
rect 52692 15200 52756 15204
rect 52772 15260 52836 15264
rect 52772 15204 52776 15260
rect 52776 15204 52832 15260
rect 52832 15204 52836 15260
rect 52772 15200 52836 15204
rect 52852 15260 52916 15264
rect 52852 15204 52856 15260
rect 52856 15204 52912 15260
rect 52912 15204 52916 15260
rect 52852 15200 52916 15204
rect 57612 15260 57676 15264
rect 57612 15204 57616 15260
rect 57616 15204 57672 15260
rect 57672 15204 57676 15260
rect 57612 15200 57676 15204
rect 57692 15260 57756 15264
rect 57692 15204 57696 15260
rect 57696 15204 57752 15260
rect 57752 15204 57756 15260
rect 57692 15200 57756 15204
rect 57772 15260 57836 15264
rect 57772 15204 57776 15260
rect 57776 15204 57832 15260
rect 57832 15204 57836 15260
rect 57772 15200 57836 15204
rect 57852 15260 57916 15264
rect 57852 15204 57856 15260
rect 57856 15204 57912 15260
rect 57912 15204 57916 15260
rect 57852 15200 57916 15204
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 21952 14716 22016 14720
rect 21952 14660 21956 14716
rect 21956 14660 22012 14716
rect 22012 14660 22016 14716
rect 21952 14656 22016 14660
rect 22032 14716 22096 14720
rect 22032 14660 22036 14716
rect 22036 14660 22092 14716
rect 22092 14660 22096 14716
rect 22032 14656 22096 14660
rect 22112 14716 22176 14720
rect 22112 14660 22116 14716
rect 22116 14660 22172 14716
rect 22172 14660 22176 14716
rect 22112 14656 22176 14660
rect 22192 14716 22256 14720
rect 22192 14660 22196 14716
rect 22196 14660 22252 14716
rect 22252 14660 22256 14716
rect 22192 14656 22256 14660
rect 26952 14716 27016 14720
rect 26952 14660 26956 14716
rect 26956 14660 27012 14716
rect 27012 14660 27016 14716
rect 26952 14656 27016 14660
rect 27032 14716 27096 14720
rect 27032 14660 27036 14716
rect 27036 14660 27092 14716
rect 27092 14660 27096 14716
rect 27032 14656 27096 14660
rect 27112 14716 27176 14720
rect 27112 14660 27116 14716
rect 27116 14660 27172 14716
rect 27172 14660 27176 14716
rect 27112 14656 27176 14660
rect 27192 14716 27256 14720
rect 27192 14660 27196 14716
rect 27196 14660 27252 14716
rect 27252 14660 27256 14716
rect 27192 14656 27256 14660
rect 31952 14716 32016 14720
rect 31952 14660 31956 14716
rect 31956 14660 32012 14716
rect 32012 14660 32016 14716
rect 31952 14656 32016 14660
rect 32032 14716 32096 14720
rect 32032 14660 32036 14716
rect 32036 14660 32092 14716
rect 32092 14660 32096 14716
rect 32032 14656 32096 14660
rect 32112 14716 32176 14720
rect 32112 14660 32116 14716
rect 32116 14660 32172 14716
rect 32172 14660 32176 14716
rect 32112 14656 32176 14660
rect 32192 14716 32256 14720
rect 32192 14660 32196 14716
rect 32196 14660 32252 14716
rect 32252 14660 32256 14716
rect 32192 14656 32256 14660
rect 36952 14716 37016 14720
rect 36952 14660 36956 14716
rect 36956 14660 37012 14716
rect 37012 14660 37016 14716
rect 36952 14656 37016 14660
rect 37032 14716 37096 14720
rect 37032 14660 37036 14716
rect 37036 14660 37092 14716
rect 37092 14660 37096 14716
rect 37032 14656 37096 14660
rect 37112 14716 37176 14720
rect 37112 14660 37116 14716
rect 37116 14660 37172 14716
rect 37172 14660 37176 14716
rect 37112 14656 37176 14660
rect 37192 14716 37256 14720
rect 37192 14660 37196 14716
rect 37196 14660 37252 14716
rect 37252 14660 37256 14716
rect 37192 14656 37256 14660
rect 41952 14716 42016 14720
rect 41952 14660 41956 14716
rect 41956 14660 42012 14716
rect 42012 14660 42016 14716
rect 41952 14656 42016 14660
rect 42032 14716 42096 14720
rect 42032 14660 42036 14716
rect 42036 14660 42092 14716
rect 42092 14660 42096 14716
rect 42032 14656 42096 14660
rect 42112 14716 42176 14720
rect 42112 14660 42116 14716
rect 42116 14660 42172 14716
rect 42172 14660 42176 14716
rect 42112 14656 42176 14660
rect 42192 14716 42256 14720
rect 42192 14660 42196 14716
rect 42196 14660 42252 14716
rect 42252 14660 42256 14716
rect 42192 14656 42256 14660
rect 46952 14716 47016 14720
rect 46952 14660 46956 14716
rect 46956 14660 47012 14716
rect 47012 14660 47016 14716
rect 46952 14656 47016 14660
rect 47032 14716 47096 14720
rect 47032 14660 47036 14716
rect 47036 14660 47092 14716
rect 47092 14660 47096 14716
rect 47032 14656 47096 14660
rect 47112 14716 47176 14720
rect 47112 14660 47116 14716
rect 47116 14660 47172 14716
rect 47172 14660 47176 14716
rect 47112 14656 47176 14660
rect 47192 14716 47256 14720
rect 47192 14660 47196 14716
rect 47196 14660 47252 14716
rect 47252 14660 47256 14716
rect 47192 14656 47256 14660
rect 51952 14716 52016 14720
rect 51952 14660 51956 14716
rect 51956 14660 52012 14716
rect 52012 14660 52016 14716
rect 51952 14656 52016 14660
rect 52032 14716 52096 14720
rect 52032 14660 52036 14716
rect 52036 14660 52092 14716
rect 52092 14660 52096 14716
rect 52032 14656 52096 14660
rect 52112 14716 52176 14720
rect 52112 14660 52116 14716
rect 52116 14660 52172 14716
rect 52172 14660 52176 14716
rect 52112 14656 52176 14660
rect 52192 14716 52256 14720
rect 52192 14660 52196 14716
rect 52196 14660 52252 14716
rect 52252 14660 52256 14716
rect 52192 14656 52256 14660
rect 56952 14716 57016 14720
rect 56952 14660 56956 14716
rect 56956 14660 57012 14716
rect 57012 14660 57016 14716
rect 56952 14656 57016 14660
rect 57032 14716 57096 14720
rect 57032 14660 57036 14716
rect 57036 14660 57092 14716
rect 57092 14660 57096 14716
rect 57032 14656 57096 14660
rect 57112 14716 57176 14720
rect 57112 14660 57116 14716
rect 57116 14660 57172 14716
rect 57172 14660 57176 14716
rect 57112 14656 57176 14660
rect 57192 14716 57256 14720
rect 57192 14660 57196 14716
rect 57196 14660 57252 14716
rect 57252 14660 57256 14716
rect 57192 14656 57256 14660
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 22612 14172 22676 14176
rect 22612 14116 22616 14172
rect 22616 14116 22672 14172
rect 22672 14116 22676 14172
rect 22612 14112 22676 14116
rect 22692 14172 22756 14176
rect 22692 14116 22696 14172
rect 22696 14116 22752 14172
rect 22752 14116 22756 14172
rect 22692 14112 22756 14116
rect 22772 14172 22836 14176
rect 22772 14116 22776 14172
rect 22776 14116 22832 14172
rect 22832 14116 22836 14172
rect 22772 14112 22836 14116
rect 22852 14172 22916 14176
rect 22852 14116 22856 14172
rect 22856 14116 22912 14172
rect 22912 14116 22916 14172
rect 22852 14112 22916 14116
rect 27612 14172 27676 14176
rect 27612 14116 27616 14172
rect 27616 14116 27672 14172
rect 27672 14116 27676 14172
rect 27612 14112 27676 14116
rect 27692 14172 27756 14176
rect 27692 14116 27696 14172
rect 27696 14116 27752 14172
rect 27752 14116 27756 14172
rect 27692 14112 27756 14116
rect 27772 14172 27836 14176
rect 27772 14116 27776 14172
rect 27776 14116 27832 14172
rect 27832 14116 27836 14172
rect 27772 14112 27836 14116
rect 27852 14172 27916 14176
rect 27852 14116 27856 14172
rect 27856 14116 27912 14172
rect 27912 14116 27916 14172
rect 27852 14112 27916 14116
rect 32612 14172 32676 14176
rect 32612 14116 32616 14172
rect 32616 14116 32672 14172
rect 32672 14116 32676 14172
rect 32612 14112 32676 14116
rect 32692 14172 32756 14176
rect 32692 14116 32696 14172
rect 32696 14116 32752 14172
rect 32752 14116 32756 14172
rect 32692 14112 32756 14116
rect 32772 14172 32836 14176
rect 32772 14116 32776 14172
rect 32776 14116 32832 14172
rect 32832 14116 32836 14172
rect 32772 14112 32836 14116
rect 32852 14172 32916 14176
rect 32852 14116 32856 14172
rect 32856 14116 32912 14172
rect 32912 14116 32916 14172
rect 32852 14112 32916 14116
rect 37612 14172 37676 14176
rect 37612 14116 37616 14172
rect 37616 14116 37672 14172
rect 37672 14116 37676 14172
rect 37612 14112 37676 14116
rect 37692 14172 37756 14176
rect 37692 14116 37696 14172
rect 37696 14116 37752 14172
rect 37752 14116 37756 14172
rect 37692 14112 37756 14116
rect 37772 14172 37836 14176
rect 37772 14116 37776 14172
rect 37776 14116 37832 14172
rect 37832 14116 37836 14172
rect 37772 14112 37836 14116
rect 37852 14172 37916 14176
rect 37852 14116 37856 14172
rect 37856 14116 37912 14172
rect 37912 14116 37916 14172
rect 37852 14112 37916 14116
rect 42612 14172 42676 14176
rect 42612 14116 42616 14172
rect 42616 14116 42672 14172
rect 42672 14116 42676 14172
rect 42612 14112 42676 14116
rect 42692 14172 42756 14176
rect 42692 14116 42696 14172
rect 42696 14116 42752 14172
rect 42752 14116 42756 14172
rect 42692 14112 42756 14116
rect 42772 14172 42836 14176
rect 42772 14116 42776 14172
rect 42776 14116 42832 14172
rect 42832 14116 42836 14172
rect 42772 14112 42836 14116
rect 42852 14172 42916 14176
rect 42852 14116 42856 14172
rect 42856 14116 42912 14172
rect 42912 14116 42916 14172
rect 42852 14112 42916 14116
rect 47612 14172 47676 14176
rect 47612 14116 47616 14172
rect 47616 14116 47672 14172
rect 47672 14116 47676 14172
rect 47612 14112 47676 14116
rect 47692 14172 47756 14176
rect 47692 14116 47696 14172
rect 47696 14116 47752 14172
rect 47752 14116 47756 14172
rect 47692 14112 47756 14116
rect 47772 14172 47836 14176
rect 47772 14116 47776 14172
rect 47776 14116 47832 14172
rect 47832 14116 47836 14172
rect 47772 14112 47836 14116
rect 47852 14172 47916 14176
rect 47852 14116 47856 14172
rect 47856 14116 47912 14172
rect 47912 14116 47916 14172
rect 47852 14112 47916 14116
rect 52612 14172 52676 14176
rect 52612 14116 52616 14172
rect 52616 14116 52672 14172
rect 52672 14116 52676 14172
rect 52612 14112 52676 14116
rect 52692 14172 52756 14176
rect 52692 14116 52696 14172
rect 52696 14116 52752 14172
rect 52752 14116 52756 14172
rect 52692 14112 52756 14116
rect 52772 14172 52836 14176
rect 52772 14116 52776 14172
rect 52776 14116 52832 14172
rect 52832 14116 52836 14172
rect 52772 14112 52836 14116
rect 52852 14172 52916 14176
rect 52852 14116 52856 14172
rect 52856 14116 52912 14172
rect 52912 14116 52916 14172
rect 52852 14112 52916 14116
rect 57612 14172 57676 14176
rect 57612 14116 57616 14172
rect 57616 14116 57672 14172
rect 57672 14116 57676 14172
rect 57612 14112 57676 14116
rect 57692 14172 57756 14176
rect 57692 14116 57696 14172
rect 57696 14116 57752 14172
rect 57752 14116 57756 14172
rect 57692 14112 57756 14116
rect 57772 14172 57836 14176
rect 57772 14116 57776 14172
rect 57776 14116 57832 14172
rect 57832 14116 57836 14172
rect 57772 14112 57836 14116
rect 57852 14172 57916 14176
rect 57852 14116 57856 14172
rect 57856 14116 57912 14172
rect 57912 14116 57916 14172
rect 57852 14112 57916 14116
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 21952 13628 22016 13632
rect 21952 13572 21956 13628
rect 21956 13572 22012 13628
rect 22012 13572 22016 13628
rect 21952 13568 22016 13572
rect 22032 13628 22096 13632
rect 22032 13572 22036 13628
rect 22036 13572 22092 13628
rect 22092 13572 22096 13628
rect 22032 13568 22096 13572
rect 22112 13628 22176 13632
rect 22112 13572 22116 13628
rect 22116 13572 22172 13628
rect 22172 13572 22176 13628
rect 22112 13568 22176 13572
rect 22192 13628 22256 13632
rect 22192 13572 22196 13628
rect 22196 13572 22252 13628
rect 22252 13572 22256 13628
rect 22192 13568 22256 13572
rect 26952 13628 27016 13632
rect 26952 13572 26956 13628
rect 26956 13572 27012 13628
rect 27012 13572 27016 13628
rect 26952 13568 27016 13572
rect 27032 13628 27096 13632
rect 27032 13572 27036 13628
rect 27036 13572 27092 13628
rect 27092 13572 27096 13628
rect 27032 13568 27096 13572
rect 27112 13628 27176 13632
rect 27112 13572 27116 13628
rect 27116 13572 27172 13628
rect 27172 13572 27176 13628
rect 27112 13568 27176 13572
rect 27192 13628 27256 13632
rect 27192 13572 27196 13628
rect 27196 13572 27252 13628
rect 27252 13572 27256 13628
rect 27192 13568 27256 13572
rect 31952 13628 32016 13632
rect 31952 13572 31956 13628
rect 31956 13572 32012 13628
rect 32012 13572 32016 13628
rect 31952 13568 32016 13572
rect 32032 13628 32096 13632
rect 32032 13572 32036 13628
rect 32036 13572 32092 13628
rect 32092 13572 32096 13628
rect 32032 13568 32096 13572
rect 32112 13628 32176 13632
rect 32112 13572 32116 13628
rect 32116 13572 32172 13628
rect 32172 13572 32176 13628
rect 32112 13568 32176 13572
rect 32192 13628 32256 13632
rect 32192 13572 32196 13628
rect 32196 13572 32252 13628
rect 32252 13572 32256 13628
rect 32192 13568 32256 13572
rect 36952 13628 37016 13632
rect 36952 13572 36956 13628
rect 36956 13572 37012 13628
rect 37012 13572 37016 13628
rect 36952 13568 37016 13572
rect 37032 13628 37096 13632
rect 37032 13572 37036 13628
rect 37036 13572 37092 13628
rect 37092 13572 37096 13628
rect 37032 13568 37096 13572
rect 37112 13628 37176 13632
rect 37112 13572 37116 13628
rect 37116 13572 37172 13628
rect 37172 13572 37176 13628
rect 37112 13568 37176 13572
rect 37192 13628 37256 13632
rect 37192 13572 37196 13628
rect 37196 13572 37252 13628
rect 37252 13572 37256 13628
rect 37192 13568 37256 13572
rect 41952 13628 42016 13632
rect 41952 13572 41956 13628
rect 41956 13572 42012 13628
rect 42012 13572 42016 13628
rect 41952 13568 42016 13572
rect 42032 13628 42096 13632
rect 42032 13572 42036 13628
rect 42036 13572 42092 13628
rect 42092 13572 42096 13628
rect 42032 13568 42096 13572
rect 42112 13628 42176 13632
rect 42112 13572 42116 13628
rect 42116 13572 42172 13628
rect 42172 13572 42176 13628
rect 42112 13568 42176 13572
rect 42192 13628 42256 13632
rect 42192 13572 42196 13628
rect 42196 13572 42252 13628
rect 42252 13572 42256 13628
rect 42192 13568 42256 13572
rect 46952 13628 47016 13632
rect 46952 13572 46956 13628
rect 46956 13572 47012 13628
rect 47012 13572 47016 13628
rect 46952 13568 47016 13572
rect 47032 13628 47096 13632
rect 47032 13572 47036 13628
rect 47036 13572 47092 13628
rect 47092 13572 47096 13628
rect 47032 13568 47096 13572
rect 47112 13628 47176 13632
rect 47112 13572 47116 13628
rect 47116 13572 47172 13628
rect 47172 13572 47176 13628
rect 47112 13568 47176 13572
rect 47192 13628 47256 13632
rect 47192 13572 47196 13628
rect 47196 13572 47252 13628
rect 47252 13572 47256 13628
rect 47192 13568 47256 13572
rect 51952 13628 52016 13632
rect 51952 13572 51956 13628
rect 51956 13572 52012 13628
rect 52012 13572 52016 13628
rect 51952 13568 52016 13572
rect 52032 13628 52096 13632
rect 52032 13572 52036 13628
rect 52036 13572 52092 13628
rect 52092 13572 52096 13628
rect 52032 13568 52096 13572
rect 52112 13628 52176 13632
rect 52112 13572 52116 13628
rect 52116 13572 52172 13628
rect 52172 13572 52176 13628
rect 52112 13568 52176 13572
rect 52192 13628 52256 13632
rect 52192 13572 52196 13628
rect 52196 13572 52252 13628
rect 52252 13572 52256 13628
rect 52192 13568 52256 13572
rect 56952 13628 57016 13632
rect 56952 13572 56956 13628
rect 56956 13572 57012 13628
rect 57012 13572 57016 13628
rect 56952 13568 57016 13572
rect 57032 13628 57096 13632
rect 57032 13572 57036 13628
rect 57036 13572 57092 13628
rect 57092 13572 57096 13628
rect 57032 13568 57096 13572
rect 57112 13628 57176 13632
rect 57112 13572 57116 13628
rect 57116 13572 57172 13628
rect 57172 13572 57176 13628
rect 57112 13568 57176 13572
rect 57192 13628 57256 13632
rect 57192 13572 57196 13628
rect 57196 13572 57252 13628
rect 57252 13572 57256 13628
rect 57192 13568 57256 13572
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 22612 13084 22676 13088
rect 22612 13028 22616 13084
rect 22616 13028 22672 13084
rect 22672 13028 22676 13084
rect 22612 13024 22676 13028
rect 22692 13084 22756 13088
rect 22692 13028 22696 13084
rect 22696 13028 22752 13084
rect 22752 13028 22756 13084
rect 22692 13024 22756 13028
rect 22772 13084 22836 13088
rect 22772 13028 22776 13084
rect 22776 13028 22832 13084
rect 22832 13028 22836 13084
rect 22772 13024 22836 13028
rect 22852 13084 22916 13088
rect 22852 13028 22856 13084
rect 22856 13028 22912 13084
rect 22912 13028 22916 13084
rect 22852 13024 22916 13028
rect 27612 13084 27676 13088
rect 27612 13028 27616 13084
rect 27616 13028 27672 13084
rect 27672 13028 27676 13084
rect 27612 13024 27676 13028
rect 27692 13084 27756 13088
rect 27692 13028 27696 13084
rect 27696 13028 27752 13084
rect 27752 13028 27756 13084
rect 27692 13024 27756 13028
rect 27772 13084 27836 13088
rect 27772 13028 27776 13084
rect 27776 13028 27832 13084
rect 27832 13028 27836 13084
rect 27772 13024 27836 13028
rect 27852 13084 27916 13088
rect 27852 13028 27856 13084
rect 27856 13028 27912 13084
rect 27912 13028 27916 13084
rect 27852 13024 27916 13028
rect 32612 13084 32676 13088
rect 32612 13028 32616 13084
rect 32616 13028 32672 13084
rect 32672 13028 32676 13084
rect 32612 13024 32676 13028
rect 32692 13084 32756 13088
rect 32692 13028 32696 13084
rect 32696 13028 32752 13084
rect 32752 13028 32756 13084
rect 32692 13024 32756 13028
rect 32772 13084 32836 13088
rect 32772 13028 32776 13084
rect 32776 13028 32832 13084
rect 32832 13028 32836 13084
rect 32772 13024 32836 13028
rect 32852 13084 32916 13088
rect 32852 13028 32856 13084
rect 32856 13028 32912 13084
rect 32912 13028 32916 13084
rect 32852 13024 32916 13028
rect 37612 13084 37676 13088
rect 37612 13028 37616 13084
rect 37616 13028 37672 13084
rect 37672 13028 37676 13084
rect 37612 13024 37676 13028
rect 37692 13084 37756 13088
rect 37692 13028 37696 13084
rect 37696 13028 37752 13084
rect 37752 13028 37756 13084
rect 37692 13024 37756 13028
rect 37772 13084 37836 13088
rect 37772 13028 37776 13084
rect 37776 13028 37832 13084
rect 37832 13028 37836 13084
rect 37772 13024 37836 13028
rect 37852 13084 37916 13088
rect 37852 13028 37856 13084
rect 37856 13028 37912 13084
rect 37912 13028 37916 13084
rect 37852 13024 37916 13028
rect 42612 13084 42676 13088
rect 42612 13028 42616 13084
rect 42616 13028 42672 13084
rect 42672 13028 42676 13084
rect 42612 13024 42676 13028
rect 42692 13084 42756 13088
rect 42692 13028 42696 13084
rect 42696 13028 42752 13084
rect 42752 13028 42756 13084
rect 42692 13024 42756 13028
rect 42772 13084 42836 13088
rect 42772 13028 42776 13084
rect 42776 13028 42832 13084
rect 42832 13028 42836 13084
rect 42772 13024 42836 13028
rect 42852 13084 42916 13088
rect 42852 13028 42856 13084
rect 42856 13028 42912 13084
rect 42912 13028 42916 13084
rect 42852 13024 42916 13028
rect 47612 13084 47676 13088
rect 47612 13028 47616 13084
rect 47616 13028 47672 13084
rect 47672 13028 47676 13084
rect 47612 13024 47676 13028
rect 47692 13084 47756 13088
rect 47692 13028 47696 13084
rect 47696 13028 47752 13084
rect 47752 13028 47756 13084
rect 47692 13024 47756 13028
rect 47772 13084 47836 13088
rect 47772 13028 47776 13084
rect 47776 13028 47832 13084
rect 47832 13028 47836 13084
rect 47772 13024 47836 13028
rect 47852 13084 47916 13088
rect 47852 13028 47856 13084
rect 47856 13028 47912 13084
rect 47912 13028 47916 13084
rect 47852 13024 47916 13028
rect 52612 13084 52676 13088
rect 52612 13028 52616 13084
rect 52616 13028 52672 13084
rect 52672 13028 52676 13084
rect 52612 13024 52676 13028
rect 52692 13084 52756 13088
rect 52692 13028 52696 13084
rect 52696 13028 52752 13084
rect 52752 13028 52756 13084
rect 52692 13024 52756 13028
rect 52772 13084 52836 13088
rect 52772 13028 52776 13084
rect 52776 13028 52832 13084
rect 52832 13028 52836 13084
rect 52772 13024 52836 13028
rect 52852 13084 52916 13088
rect 52852 13028 52856 13084
rect 52856 13028 52912 13084
rect 52912 13028 52916 13084
rect 52852 13024 52916 13028
rect 57612 13084 57676 13088
rect 57612 13028 57616 13084
rect 57616 13028 57672 13084
rect 57672 13028 57676 13084
rect 57612 13024 57676 13028
rect 57692 13084 57756 13088
rect 57692 13028 57696 13084
rect 57696 13028 57752 13084
rect 57752 13028 57756 13084
rect 57692 13024 57756 13028
rect 57772 13084 57836 13088
rect 57772 13028 57776 13084
rect 57776 13028 57832 13084
rect 57832 13028 57836 13084
rect 57772 13024 57836 13028
rect 57852 13084 57916 13088
rect 57852 13028 57856 13084
rect 57856 13028 57912 13084
rect 57912 13028 57916 13084
rect 57852 13024 57916 13028
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 21952 12540 22016 12544
rect 21952 12484 21956 12540
rect 21956 12484 22012 12540
rect 22012 12484 22016 12540
rect 21952 12480 22016 12484
rect 22032 12540 22096 12544
rect 22032 12484 22036 12540
rect 22036 12484 22092 12540
rect 22092 12484 22096 12540
rect 22032 12480 22096 12484
rect 22112 12540 22176 12544
rect 22112 12484 22116 12540
rect 22116 12484 22172 12540
rect 22172 12484 22176 12540
rect 22112 12480 22176 12484
rect 22192 12540 22256 12544
rect 22192 12484 22196 12540
rect 22196 12484 22252 12540
rect 22252 12484 22256 12540
rect 22192 12480 22256 12484
rect 26952 12540 27016 12544
rect 26952 12484 26956 12540
rect 26956 12484 27012 12540
rect 27012 12484 27016 12540
rect 26952 12480 27016 12484
rect 27032 12540 27096 12544
rect 27032 12484 27036 12540
rect 27036 12484 27092 12540
rect 27092 12484 27096 12540
rect 27032 12480 27096 12484
rect 27112 12540 27176 12544
rect 27112 12484 27116 12540
rect 27116 12484 27172 12540
rect 27172 12484 27176 12540
rect 27112 12480 27176 12484
rect 27192 12540 27256 12544
rect 27192 12484 27196 12540
rect 27196 12484 27252 12540
rect 27252 12484 27256 12540
rect 27192 12480 27256 12484
rect 31952 12540 32016 12544
rect 31952 12484 31956 12540
rect 31956 12484 32012 12540
rect 32012 12484 32016 12540
rect 31952 12480 32016 12484
rect 32032 12540 32096 12544
rect 32032 12484 32036 12540
rect 32036 12484 32092 12540
rect 32092 12484 32096 12540
rect 32032 12480 32096 12484
rect 32112 12540 32176 12544
rect 32112 12484 32116 12540
rect 32116 12484 32172 12540
rect 32172 12484 32176 12540
rect 32112 12480 32176 12484
rect 32192 12540 32256 12544
rect 32192 12484 32196 12540
rect 32196 12484 32252 12540
rect 32252 12484 32256 12540
rect 32192 12480 32256 12484
rect 36952 12540 37016 12544
rect 36952 12484 36956 12540
rect 36956 12484 37012 12540
rect 37012 12484 37016 12540
rect 36952 12480 37016 12484
rect 37032 12540 37096 12544
rect 37032 12484 37036 12540
rect 37036 12484 37092 12540
rect 37092 12484 37096 12540
rect 37032 12480 37096 12484
rect 37112 12540 37176 12544
rect 37112 12484 37116 12540
rect 37116 12484 37172 12540
rect 37172 12484 37176 12540
rect 37112 12480 37176 12484
rect 37192 12540 37256 12544
rect 37192 12484 37196 12540
rect 37196 12484 37252 12540
rect 37252 12484 37256 12540
rect 37192 12480 37256 12484
rect 41952 12540 42016 12544
rect 41952 12484 41956 12540
rect 41956 12484 42012 12540
rect 42012 12484 42016 12540
rect 41952 12480 42016 12484
rect 42032 12540 42096 12544
rect 42032 12484 42036 12540
rect 42036 12484 42092 12540
rect 42092 12484 42096 12540
rect 42032 12480 42096 12484
rect 42112 12540 42176 12544
rect 42112 12484 42116 12540
rect 42116 12484 42172 12540
rect 42172 12484 42176 12540
rect 42112 12480 42176 12484
rect 42192 12540 42256 12544
rect 42192 12484 42196 12540
rect 42196 12484 42252 12540
rect 42252 12484 42256 12540
rect 42192 12480 42256 12484
rect 46952 12540 47016 12544
rect 46952 12484 46956 12540
rect 46956 12484 47012 12540
rect 47012 12484 47016 12540
rect 46952 12480 47016 12484
rect 47032 12540 47096 12544
rect 47032 12484 47036 12540
rect 47036 12484 47092 12540
rect 47092 12484 47096 12540
rect 47032 12480 47096 12484
rect 47112 12540 47176 12544
rect 47112 12484 47116 12540
rect 47116 12484 47172 12540
rect 47172 12484 47176 12540
rect 47112 12480 47176 12484
rect 47192 12540 47256 12544
rect 47192 12484 47196 12540
rect 47196 12484 47252 12540
rect 47252 12484 47256 12540
rect 47192 12480 47256 12484
rect 51952 12540 52016 12544
rect 51952 12484 51956 12540
rect 51956 12484 52012 12540
rect 52012 12484 52016 12540
rect 51952 12480 52016 12484
rect 52032 12540 52096 12544
rect 52032 12484 52036 12540
rect 52036 12484 52092 12540
rect 52092 12484 52096 12540
rect 52032 12480 52096 12484
rect 52112 12540 52176 12544
rect 52112 12484 52116 12540
rect 52116 12484 52172 12540
rect 52172 12484 52176 12540
rect 52112 12480 52176 12484
rect 52192 12540 52256 12544
rect 52192 12484 52196 12540
rect 52196 12484 52252 12540
rect 52252 12484 52256 12540
rect 52192 12480 52256 12484
rect 56952 12540 57016 12544
rect 56952 12484 56956 12540
rect 56956 12484 57012 12540
rect 57012 12484 57016 12540
rect 56952 12480 57016 12484
rect 57032 12540 57096 12544
rect 57032 12484 57036 12540
rect 57036 12484 57092 12540
rect 57092 12484 57096 12540
rect 57032 12480 57096 12484
rect 57112 12540 57176 12544
rect 57112 12484 57116 12540
rect 57116 12484 57172 12540
rect 57172 12484 57176 12540
rect 57112 12480 57176 12484
rect 57192 12540 57256 12544
rect 57192 12484 57196 12540
rect 57196 12484 57252 12540
rect 57252 12484 57256 12540
rect 57192 12480 57256 12484
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 22612 11996 22676 12000
rect 22612 11940 22616 11996
rect 22616 11940 22672 11996
rect 22672 11940 22676 11996
rect 22612 11936 22676 11940
rect 22692 11996 22756 12000
rect 22692 11940 22696 11996
rect 22696 11940 22752 11996
rect 22752 11940 22756 11996
rect 22692 11936 22756 11940
rect 22772 11996 22836 12000
rect 22772 11940 22776 11996
rect 22776 11940 22832 11996
rect 22832 11940 22836 11996
rect 22772 11936 22836 11940
rect 22852 11996 22916 12000
rect 22852 11940 22856 11996
rect 22856 11940 22912 11996
rect 22912 11940 22916 11996
rect 22852 11936 22916 11940
rect 27612 11996 27676 12000
rect 27612 11940 27616 11996
rect 27616 11940 27672 11996
rect 27672 11940 27676 11996
rect 27612 11936 27676 11940
rect 27692 11996 27756 12000
rect 27692 11940 27696 11996
rect 27696 11940 27752 11996
rect 27752 11940 27756 11996
rect 27692 11936 27756 11940
rect 27772 11996 27836 12000
rect 27772 11940 27776 11996
rect 27776 11940 27832 11996
rect 27832 11940 27836 11996
rect 27772 11936 27836 11940
rect 27852 11996 27916 12000
rect 27852 11940 27856 11996
rect 27856 11940 27912 11996
rect 27912 11940 27916 11996
rect 27852 11936 27916 11940
rect 32612 11996 32676 12000
rect 32612 11940 32616 11996
rect 32616 11940 32672 11996
rect 32672 11940 32676 11996
rect 32612 11936 32676 11940
rect 32692 11996 32756 12000
rect 32692 11940 32696 11996
rect 32696 11940 32752 11996
rect 32752 11940 32756 11996
rect 32692 11936 32756 11940
rect 32772 11996 32836 12000
rect 32772 11940 32776 11996
rect 32776 11940 32832 11996
rect 32832 11940 32836 11996
rect 32772 11936 32836 11940
rect 32852 11996 32916 12000
rect 32852 11940 32856 11996
rect 32856 11940 32912 11996
rect 32912 11940 32916 11996
rect 32852 11936 32916 11940
rect 37612 11996 37676 12000
rect 37612 11940 37616 11996
rect 37616 11940 37672 11996
rect 37672 11940 37676 11996
rect 37612 11936 37676 11940
rect 37692 11996 37756 12000
rect 37692 11940 37696 11996
rect 37696 11940 37752 11996
rect 37752 11940 37756 11996
rect 37692 11936 37756 11940
rect 37772 11996 37836 12000
rect 37772 11940 37776 11996
rect 37776 11940 37832 11996
rect 37832 11940 37836 11996
rect 37772 11936 37836 11940
rect 37852 11996 37916 12000
rect 37852 11940 37856 11996
rect 37856 11940 37912 11996
rect 37912 11940 37916 11996
rect 37852 11936 37916 11940
rect 42612 11996 42676 12000
rect 42612 11940 42616 11996
rect 42616 11940 42672 11996
rect 42672 11940 42676 11996
rect 42612 11936 42676 11940
rect 42692 11996 42756 12000
rect 42692 11940 42696 11996
rect 42696 11940 42752 11996
rect 42752 11940 42756 11996
rect 42692 11936 42756 11940
rect 42772 11996 42836 12000
rect 42772 11940 42776 11996
rect 42776 11940 42832 11996
rect 42832 11940 42836 11996
rect 42772 11936 42836 11940
rect 42852 11996 42916 12000
rect 42852 11940 42856 11996
rect 42856 11940 42912 11996
rect 42912 11940 42916 11996
rect 42852 11936 42916 11940
rect 47612 11996 47676 12000
rect 47612 11940 47616 11996
rect 47616 11940 47672 11996
rect 47672 11940 47676 11996
rect 47612 11936 47676 11940
rect 47692 11996 47756 12000
rect 47692 11940 47696 11996
rect 47696 11940 47752 11996
rect 47752 11940 47756 11996
rect 47692 11936 47756 11940
rect 47772 11996 47836 12000
rect 47772 11940 47776 11996
rect 47776 11940 47832 11996
rect 47832 11940 47836 11996
rect 47772 11936 47836 11940
rect 47852 11996 47916 12000
rect 47852 11940 47856 11996
rect 47856 11940 47912 11996
rect 47912 11940 47916 11996
rect 47852 11936 47916 11940
rect 52612 11996 52676 12000
rect 52612 11940 52616 11996
rect 52616 11940 52672 11996
rect 52672 11940 52676 11996
rect 52612 11936 52676 11940
rect 52692 11996 52756 12000
rect 52692 11940 52696 11996
rect 52696 11940 52752 11996
rect 52752 11940 52756 11996
rect 52692 11936 52756 11940
rect 52772 11996 52836 12000
rect 52772 11940 52776 11996
rect 52776 11940 52832 11996
rect 52832 11940 52836 11996
rect 52772 11936 52836 11940
rect 52852 11996 52916 12000
rect 52852 11940 52856 11996
rect 52856 11940 52912 11996
rect 52912 11940 52916 11996
rect 52852 11936 52916 11940
rect 57612 11996 57676 12000
rect 57612 11940 57616 11996
rect 57616 11940 57672 11996
rect 57672 11940 57676 11996
rect 57612 11936 57676 11940
rect 57692 11996 57756 12000
rect 57692 11940 57696 11996
rect 57696 11940 57752 11996
rect 57752 11940 57756 11996
rect 57692 11936 57756 11940
rect 57772 11996 57836 12000
rect 57772 11940 57776 11996
rect 57776 11940 57832 11996
rect 57832 11940 57836 11996
rect 57772 11936 57836 11940
rect 57852 11996 57916 12000
rect 57852 11940 57856 11996
rect 57856 11940 57912 11996
rect 57912 11940 57916 11996
rect 57852 11936 57916 11940
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 21952 11452 22016 11456
rect 21952 11396 21956 11452
rect 21956 11396 22012 11452
rect 22012 11396 22016 11452
rect 21952 11392 22016 11396
rect 22032 11452 22096 11456
rect 22032 11396 22036 11452
rect 22036 11396 22092 11452
rect 22092 11396 22096 11452
rect 22032 11392 22096 11396
rect 22112 11452 22176 11456
rect 22112 11396 22116 11452
rect 22116 11396 22172 11452
rect 22172 11396 22176 11452
rect 22112 11392 22176 11396
rect 22192 11452 22256 11456
rect 22192 11396 22196 11452
rect 22196 11396 22252 11452
rect 22252 11396 22256 11452
rect 22192 11392 22256 11396
rect 26952 11452 27016 11456
rect 26952 11396 26956 11452
rect 26956 11396 27012 11452
rect 27012 11396 27016 11452
rect 26952 11392 27016 11396
rect 27032 11452 27096 11456
rect 27032 11396 27036 11452
rect 27036 11396 27092 11452
rect 27092 11396 27096 11452
rect 27032 11392 27096 11396
rect 27112 11452 27176 11456
rect 27112 11396 27116 11452
rect 27116 11396 27172 11452
rect 27172 11396 27176 11452
rect 27112 11392 27176 11396
rect 27192 11452 27256 11456
rect 27192 11396 27196 11452
rect 27196 11396 27252 11452
rect 27252 11396 27256 11452
rect 27192 11392 27256 11396
rect 31952 11452 32016 11456
rect 31952 11396 31956 11452
rect 31956 11396 32012 11452
rect 32012 11396 32016 11452
rect 31952 11392 32016 11396
rect 32032 11452 32096 11456
rect 32032 11396 32036 11452
rect 32036 11396 32092 11452
rect 32092 11396 32096 11452
rect 32032 11392 32096 11396
rect 32112 11452 32176 11456
rect 32112 11396 32116 11452
rect 32116 11396 32172 11452
rect 32172 11396 32176 11452
rect 32112 11392 32176 11396
rect 32192 11452 32256 11456
rect 32192 11396 32196 11452
rect 32196 11396 32252 11452
rect 32252 11396 32256 11452
rect 32192 11392 32256 11396
rect 36952 11452 37016 11456
rect 36952 11396 36956 11452
rect 36956 11396 37012 11452
rect 37012 11396 37016 11452
rect 36952 11392 37016 11396
rect 37032 11452 37096 11456
rect 37032 11396 37036 11452
rect 37036 11396 37092 11452
rect 37092 11396 37096 11452
rect 37032 11392 37096 11396
rect 37112 11452 37176 11456
rect 37112 11396 37116 11452
rect 37116 11396 37172 11452
rect 37172 11396 37176 11452
rect 37112 11392 37176 11396
rect 37192 11452 37256 11456
rect 37192 11396 37196 11452
rect 37196 11396 37252 11452
rect 37252 11396 37256 11452
rect 37192 11392 37256 11396
rect 41952 11452 42016 11456
rect 41952 11396 41956 11452
rect 41956 11396 42012 11452
rect 42012 11396 42016 11452
rect 41952 11392 42016 11396
rect 42032 11452 42096 11456
rect 42032 11396 42036 11452
rect 42036 11396 42092 11452
rect 42092 11396 42096 11452
rect 42032 11392 42096 11396
rect 42112 11452 42176 11456
rect 42112 11396 42116 11452
rect 42116 11396 42172 11452
rect 42172 11396 42176 11452
rect 42112 11392 42176 11396
rect 42192 11452 42256 11456
rect 42192 11396 42196 11452
rect 42196 11396 42252 11452
rect 42252 11396 42256 11452
rect 42192 11392 42256 11396
rect 46952 11452 47016 11456
rect 46952 11396 46956 11452
rect 46956 11396 47012 11452
rect 47012 11396 47016 11452
rect 46952 11392 47016 11396
rect 47032 11452 47096 11456
rect 47032 11396 47036 11452
rect 47036 11396 47092 11452
rect 47092 11396 47096 11452
rect 47032 11392 47096 11396
rect 47112 11452 47176 11456
rect 47112 11396 47116 11452
rect 47116 11396 47172 11452
rect 47172 11396 47176 11452
rect 47112 11392 47176 11396
rect 47192 11452 47256 11456
rect 47192 11396 47196 11452
rect 47196 11396 47252 11452
rect 47252 11396 47256 11452
rect 47192 11392 47256 11396
rect 51952 11452 52016 11456
rect 51952 11396 51956 11452
rect 51956 11396 52012 11452
rect 52012 11396 52016 11452
rect 51952 11392 52016 11396
rect 52032 11452 52096 11456
rect 52032 11396 52036 11452
rect 52036 11396 52092 11452
rect 52092 11396 52096 11452
rect 52032 11392 52096 11396
rect 52112 11452 52176 11456
rect 52112 11396 52116 11452
rect 52116 11396 52172 11452
rect 52172 11396 52176 11452
rect 52112 11392 52176 11396
rect 52192 11452 52256 11456
rect 52192 11396 52196 11452
rect 52196 11396 52252 11452
rect 52252 11396 52256 11452
rect 52192 11392 52256 11396
rect 56952 11452 57016 11456
rect 56952 11396 56956 11452
rect 56956 11396 57012 11452
rect 57012 11396 57016 11452
rect 56952 11392 57016 11396
rect 57032 11452 57096 11456
rect 57032 11396 57036 11452
rect 57036 11396 57092 11452
rect 57092 11396 57096 11452
rect 57032 11392 57096 11396
rect 57112 11452 57176 11456
rect 57112 11396 57116 11452
rect 57116 11396 57172 11452
rect 57172 11396 57176 11452
rect 57112 11392 57176 11396
rect 57192 11452 57256 11456
rect 57192 11396 57196 11452
rect 57196 11396 57252 11452
rect 57252 11396 57256 11452
rect 57192 11392 57256 11396
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 22612 10908 22676 10912
rect 22612 10852 22616 10908
rect 22616 10852 22672 10908
rect 22672 10852 22676 10908
rect 22612 10848 22676 10852
rect 22692 10908 22756 10912
rect 22692 10852 22696 10908
rect 22696 10852 22752 10908
rect 22752 10852 22756 10908
rect 22692 10848 22756 10852
rect 22772 10908 22836 10912
rect 22772 10852 22776 10908
rect 22776 10852 22832 10908
rect 22832 10852 22836 10908
rect 22772 10848 22836 10852
rect 22852 10908 22916 10912
rect 22852 10852 22856 10908
rect 22856 10852 22912 10908
rect 22912 10852 22916 10908
rect 22852 10848 22916 10852
rect 27612 10908 27676 10912
rect 27612 10852 27616 10908
rect 27616 10852 27672 10908
rect 27672 10852 27676 10908
rect 27612 10848 27676 10852
rect 27692 10908 27756 10912
rect 27692 10852 27696 10908
rect 27696 10852 27752 10908
rect 27752 10852 27756 10908
rect 27692 10848 27756 10852
rect 27772 10908 27836 10912
rect 27772 10852 27776 10908
rect 27776 10852 27832 10908
rect 27832 10852 27836 10908
rect 27772 10848 27836 10852
rect 27852 10908 27916 10912
rect 27852 10852 27856 10908
rect 27856 10852 27912 10908
rect 27912 10852 27916 10908
rect 27852 10848 27916 10852
rect 32612 10908 32676 10912
rect 32612 10852 32616 10908
rect 32616 10852 32672 10908
rect 32672 10852 32676 10908
rect 32612 10848 32676 10852
rect 32692 10908 32756 10912
rect 32692 10852 32696 10908
rect 32696 10852 32752 10908
rect 32752 10852 32756 10908
rect 32692 10848 32756 10852
rect 32772 10908 32836 10912
rect 32772 10852 32776 10908
rect 32776 10852 32832 10908
rect 32832 10852 32836 10908
rect 32772 10848 32836 10852
rect 32852 10908 32916 10912
rect 32852 10852 32856 10908
rect 32856 10852 32912 10908
rect 32912 10852 32916 10908
rect 32852 10848 32916 10852
rect 37612 10908 37676 10912
rect 37612 10852 37616 10908
rect 37616 10852 37672 10908
rect 37672 10852 37676 10908
rect 37612 10848 37676 10852
rect 37692 10908 37756 10912
rect 37692 10852 37696 10908
rect 37696 10852 37752 10908
rect 37752 10852 37756 10908
rect 37692 10848 37756 10852
rect 37772 10908 37836 10912
rect 37772 10852 37776 10908
rect 37776 10852 37832 10908
rect 37832 10852 37836 10908
rect 37772 10848 37836 10852
rect 37852 10908 37916 10912
rect 37852 10852 37856 10908
rect 37856 10852 37912 10908
rect 37912 10852 37916 10908
rect 37852 10848 37916 10852
rect 42612 10908 42676 10912
rect 42612 10852 42616 10908
rect 42616 10852 42672 10908
rect 42672 10852 42676 10908
rect 42612 10848 42676 10852
rect 42692 10908 42756 10912
rect 42692 10852 42696 10908
rect 42696 10852 42752 10908
rect 42752 10852 42756 10908
rect 42692 10848 42756 10852
rect 42772 10908 42836 10912
rect 42772 10852 42776 10908
rect 42776 10852 42832 10908
rect 42832 10852 42836 10908
rect 42772 10848 42836 10852
rect 42852 10908 42916 10912
rect 42852 10852 42856 10908
rect 42856 10852 42912 10908
rect 42912 10852 42916 10908
rect 42852 10848 42916 10852
rect 47612 10908 47676 10912
rect 47612 10852 47616 10908
rect 47616 10852 47672 10908
rect 47672 10852 47676 10908
rect 47612 10848 47676 10852
rect 47692 10908 47756 10912
rect 47692 10852 47696 10908
rect 47696 10852 47752 10908
rect 47752 10852 47756 10908
rect 47692 10848 47756 10852
rect 47772 10908 47836 10912
rect 47772 10852 47776 10908
rect 47776 10852 47832 10908
rect 47832 10852 47836 10908
rect 47772 10848 47836 10852
rect 47852 10908 47916 10912
rect 47852 10852 47856 10908
rect 47856 10852 47912 10908
rect 47912 10852 47916 10908
rect 47852 10848 47916 10852
rect 52612 10908 52676 10912
rect 52612 10852 52616 10908
rect 52616 10852 52672 10908
rect 52672 10852 52676 10908
rect 52612 10848 52676 10852
rect 52692 10908 52756 10912
rect 52692 10852 52696 10908
rect 52696 10852 52752 10908
rect 52752 10852 52756 10908
rect 52692 10848 52756 10852
rect 52772 10908 52836 10912
rect 52772 10852 52776 10908
rect 52776 10852 52832 10908
rect 52832 10852 52836 10908
rect 52772 10848 52836 10852
rect 52852 10908 52916 10912
rect 52852 10852 52856 10908
rect 52856 10852 52912 10908
rect 52912 10852 52916 10908
rect 52852 10848 52916 10852
rect 57612 10908 57676 10912
rect 57612 10852 57616 10908
rect 57616 10852 57672 10908
rect 57672 10852 57676 10908
rect 57612 10848 57676 10852
rect 57692 10908 57756 10912
rect 57692 10852 57696 10908
rect 57696 10852 57752 10908
rect 57752 10852 57756 10908
rect 57692 10848 57756 10852
rect 57772 10908 57836 10912
rect 57772 10852 57776 10908
rect 57776 10852 57832 10908
rect 57832 10852 57836 10908
rect 57772 10848 57836 10852
rect 57852 10908 57916 10912
rect 57852 10852 57856 10908
rect 57856 10852 57912 10908
rect 57912 10852 57916 10908
rect 57852 10848 57916 10852
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 21952 10364 22016 10368
rect 21952 10308 21956 10364
rect 21956 10308 22012 10364
rect 22012 10308 22016 10364
rect 21952 10304 22016 10308
rect 22032 10364 22096 10368
rect 22032 10308 22036 10364
rect 22036 10308 22092 10364
rect 22092 10308 22096 10364
rect 22032 10304 22096 10308
rect 22112 10364 22176 10368
rect 22112 10308 22116 10364
rect 22116 10308 22172 10364
rect 22172 10308 22176 10364
rect 22112 10304 22176 10308
rect 22192 10364 22256 10368
rect 22192 10308 22196 10364
rect 22196 10308 22252 10364
rect 22252 10308 22256 10364
rect 22192 10304 22256 10308
rect 26952 10364 27016 10368
rect 26952 10308 26956 10364
rect 26956 10308 27012 10364
rect 27012 10308 27016 10364
rect 26952 10304 27016 10308
rect 27032 10364 27096 10368
rect 27032 10308 27036 10364
rect 27036 10308 27092 10364
rect 27092 10308 27096 10364
rect 27032 10304 27096 10308
rect 27112 10364 27176 10368
rect 27112 10308 27116 10364
rect 27116 10308 27172 10364
rect 27172 10308 27176 10364
rect 27112 10304 27176 10308
rect 27192 10364 27256 10368
rect 27192 10308 27196 10364
rect 27196 10308 27252 10364
rect 27252 10308 27256 10364
rect 27192 10304 27256 10308
rect 31952 10364 32016 10368
rect 31952 10308 31956 10364
rect 31956 10308 32012 10364
rect 32012 10308 32016 10364
rect 31952 10304 32016 10308
rect 32032 10364 32096 10368
rect 32032 10308 32036 10364
rect 32036 10308 32092 10364
rect 32092 10308 32096 10364
rect 32032 10304 32096 10308
rect 32112 10364 32176 10368
rect 32112 10308 32116 10364
rect 32116 10308 32172 10364
rect 32172 10308 32176 10364
rect 32112 10304 32176 10308
rect 32192 10364 32256 10368
rect 32192 10308 32196 10364
rect 32196 10308 32252 10364
rect 32252 10308 32256 10364
rect 32192 10304 32256 10308
rect 36952 10364 37016 10368
rect 36952 10308 36956 10364
rect 36956 10308 37012 10364
rect 37012 10308 37016 10364
rect 36952 10304 37016 10308
rect 37032 10364 37096 10368
rect 37032 10308 37036 10364
rect 37036 10308 37092 10364
rect 37092 10308 37096 10364
rect 37032 10304 37096 10308
rect 37112 10364 37176 10368
rect 37112 10308 37116 10364
rect 37116 10308 37172 10364
rect 37172 10308 37176 10364
rect 37112 10304 37176 10308
rect 37192 10364 37256 10368
rect 37192 10308 37196 10364
rect 37196 10308 37252 10364
rect 37252 10308 37256 10364
rect 37192 10304 37256 10308
rect 41952 10364 42016 10368
rect 41952 10308 41956 10364
rect 41956 10308 42012 10364
rect 42012 10308 42016 10364
rect 41952 10304 42016 10308
rect 42032 10364 42096 10368
rect 42032 10308 42036 10364
rect 42036 10308 42092 10364
rect 42092 10308 42096 10364
rect 42032 10304 42096 10308
rect 42112 10364 42176 10368
rect 42112 10308 42116 10364
rect 42116 10308 42172 10364
rect 42172 10308 42176 10364
rect 42112 10304 42176 10308
rect 42192 10364 42256 10368
rect 42192 10308 42196 10364
rect 42196 10308 42252 10364
rect 42252 10308 42256 10364
rect 42192 10304 42256 10308
rect 46952 10364 47016 10368
rect 46952 10308 46956 10364
rect 46956 10308 47012 10364
rect 47012 10308 47016 10364
rect 46952 10304 47016 10308
rect 47032 10364 47096 10368
rect 47032 10308 47036 10364
rect 47036 10308 47092 10364
rect 47092 10308 47096 10364
rect 47032 10304 47096 10308
rect 47112 10364 47176 10368
rect 47112 10308 47116 10364
rect 47116 10308 47172 10364
rect 47172 10308 47176 10364
rect 47112 10304 47176 10308
rect 47192 10364 47256 10368
rect 47192 10308 47196 10364
rect 47196 10308 47252 10364
rect 47252 10308 47256 10364
rect 47192 10304 47256 10308
rect 51952 10364 52016 10368
rect 51952 10308 51956 10364
rect 51956 10308 52012 10364
rect 52012 10308 52016 10364
rect 51952 10304 52016 10308
rect 52032 10364 52096 10368
rect 52032 10308 52036 10364
rect 52036 10308 52092 10364
rect 52092 10308 52096 10364
rect 52032 10304 52096 10308
rect 52112 10364 52176 10368
rect 52112 10308 52116 10364
rect 52116 10308 52172 10364
rect 52172 10308 52176 10364
rect 52112 10304 52176 10308
rect 52192 10364 52256 10368
rect 52192 10308 52196 10364
rect 52196 10308 52252 10364
rect 52252 10308 52256 10364
rect 52192 10304 52256 10308
rect 56952 10364 57016 10368
rect 56952 10308 56956 10364
rect 56956 10308 57012 10364
rect 57012 10308 57016 10364
rect 56952 10304 57016 10308
rect 57032 10364 57096 10368
rect 57032 10308 57036 10364
rect 57036 10308 57092 10364
rect 57092 10308 57096 10364
rect 57032 10304 57096 10308
rect 57112 10364 57176 10368
rect 57112 10308 57116 10364
rect 57116 10308 57172 10364
rect 57172 10308 57176 10364
rect 57112 10304 57176 10308
rect 57192 10364 57256 10368
rect 57192 10308 57196 10364
rect 57196 10308 57252 10364
rect 57252 10308 57256 10364
rect 57192 10304 57256 10308
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 22612 9820 22676 9824
rect 22612 9764 22616 9820
rect 22616 9764 22672 9820
rect 22672 9764 22676 9820
rect 22612 9760 22676 9764
rect 22692 9820 22756 9824
rect 22692 9764 22696 9820
rect 22696 9764 22752 9820
rect 22752 9764 22756 9820
rect 22692 9760 22756 9764
rect 22772 9820 22836 9824
rect 22772 9764 22776 9820
rect 22776 9764 22832 9820
rect 22832 9764 22836 9820
rect 22772 9760 22836 9764
rect 22852 9820 22916 9824
rect 22852 9764 22856 9820
rect 22856 9764 22912 9820
rect 22912 9764 22916 9820
rect 22852 9760 22916 9764
rect 27612 9820 27676 9824
rect 27612 9764 27616 9820
rect 27616 9764 27672 9820
rect 27672 9764 27676 9820
rect 27612 9760 27676 9764
rect 27692 9820 27756 9824
rect 27692 9764 27696 9820
rect 27696 9764 27752 9820
rect 27752 9764 27756 9820
rect 27692 9760 27756 9764
rect 27772 9820 27836 9824
rect 27772 9764 27776 9820
rect 27776 9764 27832 9820
rect 27832 9764 27836 9820
rect 27772 9760 27836 9764
rect 27852 9820 27916 9824
rect 27852 9764 27856 9820
rect 27856 9764 27912 9820
rect 27912 9764 27916 9820
rect 27852 9760 27916 9764
rect 32612 9820 32676 9824
rect 32612 9764 32616 9820
rect 32616 9764 32672 9820
rect 32672 9764 32676 9820
rect 32612 9760 32676 9764
rect 32692 9820 32756 9824
rect 32692 9764 32696 9820
rect 32696 9764 32752 9820
rect 32752 9764 32756 9820
rect 32692 9760 32756 9764
rect 32772 9820 32836 9824
rect 32772 9764 32776 9820
rect 32776 9764 32832 9820
rect 32832 9764 32836 9820
rect 32772 9760 32836 9764
rect 32852 9820 32916 9824
rect 32852 9764 32856 9820
rect 32856 9764 32912 9820
rect 32912 9764 32916 9820
rect 32852 9760 32916 9764
rect 37612 9820 37676 9824
rect 37612 9764 37616 9820
rect 37616 9764 37672 9820
rect 37672 9764 37676 9820
rect 37612 9760 37676 9764
rect 37692 9820 37756 9824
rect 37692 9764 37696 9820
rect 37696 9764 37752 9820
rect 37752 9764 37756 9820
rect 37692 9760 37756 9764
rect 37772 9820 37836 9824
rect 37772 9764 37776 9820
rect 37776 9764 37832 9820
rect 37832 9764 37836 9820
rect 37772 9760 37836 9764
rect 37852 9820 37916 9824
rect 37852 9764 37856 9820
rect 37856 9764 37912 9820
rect 37912 9764 37916 9820
rect 37852 9760 37916 9764
rect 42612 9820 42676 9824
rect 42612 9764 42616 9820
rect 42616 9764 42672 9820
rect 42672 9764 42676 9820
rect 42612 9760 42676 9764
rect 42692 9820 42756 9824
rect 42692 9764 42696 9820
rect 42696 9764 42752 9820
rect 42752 9764 42756 9820
rect 42692 9760 42756 9764
rect 42772 9820 42836 9824
rect 42772 9764 42776 9820
rect 42776 9764 42832 9820
rect 42832 9764 42836 9820
rect 42772 9760 42836 9764
rect 42852 9820 42916 9824
rect 42852 9764 42856 9820
rect 42856 9764 42912 9820
rect 42912 9764 42916 9820
rect 42852 9760 42916 9764
rect 47612 9820 47676 9824
rect 47612 9764 47616 9820
rect 47616 9764 47672 9820
rect 47672 9764 47676 9820
rect 47612 9760 47676 9764
rect 47692 9820 47756 9824
rect 47692 9764 47696 9820
rect 47696 9764 47752 9820
rect 47752 9764 47756 9820
rect 47692 9760 47756 9764
rect 47772 9820 47836 9824
rect 47772 9764 47776 9820
rect 47776 9764 47832 9820
rect 47832 9764 47836 9820
rect 47772 9760 47836 9764
rect 47852 9820 47916 9824
rect 47852 9764 47856 9820
rect 47856 9764 47912 9820
rect 47912 9764 47916 9820
rect 47852 9760 47916 9764
rect 52612 9820 52676 9824
rect 52612 9764 52616 9820
rect 52616 9764 52672 9820
rect 52672 9764 52676 9820
rect 52612 9760 52676 9764
rect 52692 9820 52756 9824
rect 52692 9764 52696 9820
rect 52696 9764 52752 9820
rect 52752 9764 52756 9820
rect 52692 9760 52756 9764
rect 52772 9820 52836 9824
rect 52772 9764 52776 9820
rect 52776 9764 52832 9820
rect 52832 9764 52836 9820
rect 52772 9760 52836 9764
rect 52852 9820 52916 9824
rect 52852 9764 52856 9820
rect 52856 9764 52912 9820
rect 52912 9764 52916 9820
rect 52852 9760 52916 9764
rect 57612 9820 57676 9824
rect 57612 9764 57616 9820
rect 57616 9764 57672 9820
rect 57672 9764 57676 9820
rect 57612 9760 57676 9764
rect 57692 9820 57756 9824
rect 57692 9764 57696 9820
rect 57696 9764 57752 9820
rect 57752 9764 57756 9820
rect 57692 9760 57756 9764
rect 57772 9820 57836 9824
rect 57772 9764 57776 9820
rect 57776 9764 57832 9820
rect 57832 9764 57836 9820
rect 57772 9760 57836 9764
rect 57852 9820 57916 9824
rect 57852 9764 57856 9820
rect 57856 9764 57912 9820
rect 57912 9764 57916 9820
rect 57852 9760 57916 9764
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 21952 9276 22016 9280
rect 21952 9220 21956 9276
rect 21956 9220 22012 9276
rect 22012 9220 22016 9276
rect 21952 9216 22016 9220
rect 22032 9276 22096 9280
rect 22032 9220 22036 9276
rect 22036 9220 22092 9276
rect 22092 9220 22096 9276
rect 22032 9216 22096 9220
rect 22112 9276 22176 9280
rect 22112 9220 22116 9276
rect 22116 9220 22172 9276
rect 22172 9220 22176 9276
rect 22112 9216 22176 9220
rect 22192 9276 22256 9280
rect 22192 9220 22196 9276
rect 22196 9220 22252 9276
rect 22252 9220 22256 9276
rect 22192 9216 22256 9220
rect 26952 9276 27016 9280
rect 26952 9220 26956 9276
rect 26956 9220 27012 9276
rect 27012 9220 27016 9276
rect 26952 9216 27016 9220
rect 27032 9276 27096 9280
rect 27032 9220 27036 9276
rect 27036 9220 27092 9276
rect 27092 9220 27096 9276
rect 27032 9216 27096 9220
rect 27112 9276 27176 9280
rect 27112 9220 27116 9276
rect 27116 9220 27172 9276
rect 27172 9220 27176 9276
rect 27112 9216 27176 9220
rect 27192 9276 27256 9280
rect 27192 9220 27196 9276
rect 27196 9220 27252 9276
rect 27252 9220 27256 9276
rect 27192 9216 27256 9220
rect 31952 9276 32016 9280
rect 31952 9220 31956 9276
rect 31956 9220 32012 9276
rect 32012 9220 32016 9276
rect 31952 9216 32016 9220
rect 32032 9276 32096 9280
rect 32032 9220 32036 9276
rect 32036 9220 32092 9276
rect 32092 9220 32096 9276
rect 32032 9216 32096 9220
rect 32112 9276 32176 9280
rect 32112 9220 32116 9276
rect 32116 9220 32172 9276
rect 32172 9220 32176 9276
rect 32112 9216 32176 9220
rect 32192 9276 32256 9280
rect 32192 9220 32196 9276
rect 32196 9220 32252 9276
rect 32252 9220 32256 9276
rect 32192 9216 32256 9220
rect 36952 9276 37016 9280
rect 36952 9220 36956 9276
rect 36956 9220 37012 9276
rect 37012 9220 37016 9276
rect 36952 9216 37016 9220
rect 37032 9276 37096 9280
rect 37032 9220 37036 9276
rect 37036 9220 37092 9276
rect 37092 9220 37096 9276
rect 37032 9216 37096 9220
rect 37112 9276 37176 9280
rect 37112 9220 37116 9276
rect 37116 9220 37172 9276
rect 37172 9220 37176 9276
rect 37112 9216 37176 9220
rect 37192 9276 37256 9280
rect 37192 9220 37196 9276
rect 37196 9220 37252 9276
rect 37252 9220 37256 9276
rect 37192 9216 37256 9220
rect 41952 9276 42016 9280
rect 41952 9220 41956 9276
rect 41956 9220 42012 9276
rect 42012 9220 42016 9276
rect 41952 9216 42016 9220
rect 42032 9276 42096 9280
rect 42032 9220 42036 9276
rect 42036 9220 42092 9276
rect 42092 9220 42096 9276
rect 42032 9216 42096 9220
rect 42112 9276 42176 9280
rect 42112 9220 42116 9276
rect 42116 9220 42172 9276
rect 42172 9220 42176 9276
rect 42112 9216 42176 9220
rect 42192 9276 42256 9280
rect 42192 9220 42196 9276
rect 42196 9220 42252 9276
rect 42252 9220 42256 9276
rect 42192 9216 42256 9220
rect 46952 9276 47016 9280
rect 46952 9220 46956 9276
rect 46956 9220 47012 9276
rect 47012 9220 47016 9276
rect 46952 9216 47016 9220
rect 47032 9276 47096 9280
rect 47032 9220 47036 9276
rect 47036 9220 47092 9276
rect 47092 9220 47096 9276
rect 47032 9216 47096 9220
rect 47112 9276 47176 9280
rect 47112 9220 47116 9276
rect 47116 9220 47172 9276
rect 47172 9220 47176 9276
rect 47112 9216 47176 9220
rect 47192 9276 47256 9280
rect 47192 9220 47196 9276
rect 47196 9220 47252 9276
rect 47252 9220 47256 9276
rect 47192 9216 47256 9220
rect 51952 9276 52016 9280
rect 51952 9220 51956 9276
rect 51956 9220 52012 9276
rect 52012 9220 52016 9276
rect 51952 9216 52016 9220
rect 52032 9276 52096 9280
rect 52032 9220 52036 9276
rect 52036 9220 52092 9276
rect 52092 9220 52096 9276
rect 52032 9216 52096 9220
rect 52112 9276 52176 9280
rect 52112 9220 52116 9276
rect 52116 9220 52172 9276
rect 52172 9220 52176 9276
rect 52112 9216 52176 9220
rect 52192 9276 52256 9280
rect 52192 9220 52196 9276
rect 52196 9220 52252 9276
rect 52252 9220 52256 9276
rect 52192 9216 52256 9220
rect 56952 9276 57016 9280
rect 56952 9220 56956 9276
rect 56956 9220 57012 9276
rect 57012 9220 57016 9276
rect 56952 9216 57016 9220
rect 57032 9276 57096 9280
rect 57032 9220 57036 9276
rect 57036 9220 57092 9276
rect 57092 9220 57096 9276
rect 57032 9216 57096 9220
rect 57112 9276 57176 9280
rect 57112 9220 57116 9276
rect 57116 9220 57172 9276
rect 57172 9220 57176 9276
rect 57112 9216 57176 9220
rect 57192 9276 57256 9280
rect 57192 9220 57196 9276
rect 57196 9220 57252 9276
rect 57252 9220 57256 9276
rect 57192 9216 57256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 22612 8732 22676 8736
rect 22612 8676 22616 8732
rect 22616 8676 22672 8732
rect 22672 8676 22676 8732
rect 22612 8672 22676 8676
rect 22692 8732 22756 8736
rect 22692 8676 22696 8732
rect 22696 8676 22752 8732
rect 22752 8676 22756 8732
rect 22692 8672 22756 8676
rect 22772 8732 22836 8736
rect 22772 8676 22776 8732
rect 22776 8676 22832 8732
rect 22832 8676 22836 8732
rect 22772 8672 22836 8676
rect 22852 8732 22916 8736
rect 22852 8676 22856 8732
rect 22856 8676 22912 8732
rect 22912 8676 22916 8732
rect 22852 8672 22916 8676
rect 27612 8732 27676 8736
rect 27612 8676 27616 8732
rect 27616 8676 27672 8732
rect 27672 8676 27676 8732
rect 27612 8672 27676 8676
rect 27692 8732 27756 8736
rect 27692 8676 27696 8732
rect 27696 8676 27752 8732
rect 27752 8676 27756 8732
rect 27692 8672 27756 8676
rect 27772 8732 27836 8736
rect 27772 8676 27776 8732
rect 27776 8676 27832 8732
rect 27832 8676 27836 8732
rect 27772 8672 27836 8676
rect 27852 8732 27916 8736
rect 27852 8676 27856 8732
rect 27856 8676 27912 8732
rect 27912 8676 27916 8732
rect 27852 8672 27916 8676
rect 32612 8732 32676 8736
rect 32612 8676 32616 8732
rect 32616 8676 32672 8732
rect 32672 8676 32676 8732
rect 32612 8672 32676 8676
rect 32692 8732 32756 8736
rect 32692 8676 32696 8732
rect 32696 8676 32752 8732
rect 32752 8676 32756 8732
rect 32692 8672 32756 8676
rect 32772 8732 32836 8736
rect 32772 8676 32776 8732
rect 32776 8676 32832 8732
rect 32832 8676 32836 8732
rect 32772 8672 32836 8676
rect 32852 8732 32916 8736
rect 32852 8676 32856 8732
rect 32856 8676 32912 8732
rect 32912 8676 32916 8732
rect 32852 8672 32916 8676
rect 37612 8732 37676 8736
rect 37612 8676 37616 8732
rect 37616 8676 37672 8732
rect 37672 8676 37676 8732
rect 37612 8672 37676 8676
rect 37692 8732 37756 8736
rect 37692 8676 37696 8732
rect 37696 8676 37752 8732
rect 37752 8676 37756 8732
rect 37692 8672 37756 8676
rect 37772 8732 37836 8736
rect 37772 8676 37776 8732
rect 37776 8676 37832 8732
rect 37832 8676 37836 8732
rect 37772 8672 37836 8676
rect 37852 8732 37916 8736
rect 37852 8676 37856 8732
rect 37856 8676 37912 8732
rect 37912 8676 37916 8732
rect 37852 8672 37916 8676
rect 42612 8732 42676 8736
rect 42612 8676 42616 8732
rect 42616 8676 42672 8732
rect 42672 8676 42676 8732
rect 42612 8672 42676 8676
rect 42692 8732 42756 8736
rect 42692 8676 42696 8732
rect 42696 8676 42752 8732
rect 42752 8676 42756 8732
rect 42692 8672 42756 8676
rect 42772 8732 42836 8736
rect 42772 8676 42776 8732
rect 42776 8676 42832 8732
rect 42832 8676 42836 8732
rect 42772 8672 42836 8676
rect 42852 8732 42916 8736
rect 42852 8676 42856 8732
rect 42856 8676 42912 8732
rect 42912 8676 42916 8732
rect 42852 8672 42916 8676
rect 47612 8732 47676 8736
rect 47612 8676 47616 8732
rect 47616 8676 47672 8732
rect 47672 8676 47676 8732
rect 47612 8672 47676 8676
rect 47692 8732 47756 8736
rect 47692 8676 47696 8732
rect 47696 8676 47752 8732
rect 47752 8676 47756 8732
rect 47692 8672 47756 8676
rect 47772 8732 47836 8736
rect 47772 8676 47776 8732
rect 47776 8676 47832 8732
rect 47832 8676 47836 8732
rect 47772 8672 47836 8676
rect 47852 8732 47916 8736
rect 47852 8676 47856 8732
rect 47856 8676 47912 8732
rect 47912 8676 47916 8732
rect 47852 8672 47916 8676
rect 52612 8732 52676 8736
rect 52612 8676 52616 8732
rect 52616 8676 52672 8732
rect 52672 8676 52676 8732
rect 52612 8672 52676 8676
rect 52692 8732 52756 8736
rect 52692 8676 52696 8732
rect 52696 8676 52752 8732
rect 52752 8676 52756 8732
rect 52692 8672 52756 8676
rect 52772 8732 52836 8736
rect 52772 8676 52776 8732
rect 52776 8676 52832 8732
rect 52832 8676 52836 8732
rect 52772 8672 52836 8676
rect 52852 8732 52916 8736
rect 52852 8676 52856 8732
rect 52856 8676 52912 8732
rect 52912 8676 52916 8732
rect 52852 8672 52916 8676
rect 57612 8732 57676 8736
rect 57612 8676 57616 8732
rect 57616 8676 57672 8732
rect 57672 8676 57676 8732
rect 57612 8672 57676 8676
rect 57692 8732 57756 8736
rect 57692 8676 57696 8732
rect 57696 8676 57752 8732
rect 57752 8676 57756 8732
rect 57692 8672 57756 8676
rect 57772 8732 57836 8736
rect 57772 8676 57776 8732
rect 57776 8676 57832 8732
rect 57832 8676 57836 8732
rect 57772 8672 57836 8676
rect 57852 8732 57916 8736
rect 57852 8676 57856 8732
rect 57856 8676 57912 8732
rect 57912 8676 57916 8732
rect 57852 8672 57916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 21952 8188 22016 8192
rect 21952 8132 21956 8188
rect 21956 8132 22012 8188
rect 22012 8132 22016 8188
rect 21952 8128 22016 8132
rect 22032 8188 22096 8192
rect 22032 8132 22036 8188
rect 22036 8132 22092 8188
rect 22092 8132 22096 8188
rect 22032 8128 22096 8132
rect 22112 8188 22176 8192
rect 22112 8132 22116 8188
rect 22116 8132 22172 8188
rect 22172 8132 22176 8188
rect 22112 8128 22176 8132
rect 22192 8188 22256 8192
rect 22192 8132 22196 8188
rect 22196 8132 22252 8188
rect 22252 8132 22256 8188
rect 22192 8128 22256 8132
rect 26952 8188 27016 8192
rect 26952 8132 26956 8188
rect 26956 8132 27012 8188
rect 27012 8132 27016 8188
rect 26952 8128 27016 8132
rect 27032 8188 27096 8192
rect 27032 8132 27036 8188
rect 27036 8132 27092 8188
rect 27092 8132 27096 8188
rect 27032 8128 27096 8132
rect 27112 8188 27176 8192
rect 27112 8132 27116 8188
rect 27116 8132 27172 8188
rect 27172 8132 27176 8188
rect 27112 8128 27176 8132
rect 27192 8188 27256 8192
rect 27192 8132 27196 8188
rect 27196 8132 27252 8188
rect 27252 8132 27256 8188
rect 27192 8128 27256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 36952 8188 37016 8192
rect 36952 8132 36956 8188
rect 36956 8132 37012 8188
rect 37012 8132 37016 8188
rect 36952 8128 37016 8132
rect 37032 8188 37096 8192
rect 37032 8132 37036 8188
rect 37036 8132 37092 8188
rect 37092 8132 37096 8188
rect 37032 8128 37096 8132
rect 37112 8188 37176 8192
rect 37112 8132 37116 8188
rect 37116 8132 37172 8188
rect 37172 8132 37176 8188
rect 37112 8128 37176 8132
rect 37192 8188 37256 8192
rect 37192 8132 37196 8188
rect 37196 8132 37252 8188
rect 37252 8132 37256 8188
rect 37192 8128 37256 8132
rect 41952 8188 42016 8192
rect 41952 8132 41956 8188
rect 41956 8132 42012 8188
rect 42012 8132 42016 8188
rect 41952 8128 42016 8132
rect 42032 8188 42096 8192
rect 42032 8132 42036 8188
rect 42036 8132 42092 8188
rect 42092 8132 42096 8188
rect 42032 8128 42096 8132
rect 42112 8188 42176 8192
rect 42112 8132 42116 8188
rect 42116 8132 42172 8188
rect 42172 8132 42176 8188
rect 42112 8128 42176 8132
rect 42192 8188 42256 8192
rect 42192 8132 42196 8188
rect 42196 8132 42252 8188
rect 42252 8132 42256 8188
rect 42192 8128 42256 8132
rect 46952 8188 47016 8192
rect 46952 8132 46956 8188
rect 46956 8132 47012 8188
rect 47012 8132 47016 8188
rect 46952 8128 47016 8132
rect 47032 8188 47096 8192
rect 47032 8132 47036 8188
rect 47036 8132 47092 8188
rect 47092 8132 47096 8188
rect 47032 8128 47096 8132
rect 47112 8188 47176 8192
rect 47112 8132 47116 8188
rect 47116 8132 47172 8188
rect 47172 8132 47176 8188
rect 47112 8128 47176 8132
rect 47192 8188 47256 8192
rect 47192 8132 47196 8188
rect 47196 8132 47252 8188
rect 47252 8132 47256 8188
rect 47192 8128 47256 8132
rect 51952 8188 52016 8192
rect 51952 8132 51956 8188
rect 51956 8132 52012 8188
rect 52012 8132 52016 8188
rect 51952 8128 52016 8132
rect 52032 8188 52096 8192
rect 52032 8132 52036 8188
rect 52036 8132 52092 8188
rect 52092 8132 52096 8188
rect 52032 8128 52096 8132
rect 52112 8188 52176 8192
rect 52112 8132 52116 8188
rect 52116 8132 52172 8188
rect 52172 8132 52176 8188
rect 52112 8128 52176 8132
rect 52192 8188 52256 8192
rect 52192 8132 52196 8188
rect 52196 8132 52252 8188
rect 52252 8132 52256 8188
rect 52192 8128 52256 8132
rect 56952 8188 57016 8192
rect 56952 8132 56956 8188
rect 56956 8132 57012 8188
rect 57012 8132 57016 8188
rect 56952 8128 57016 8132
rect 57032 8188 57096 8192
rect 57032 8132 57036 8188
rect 57036 8132 57092 8188
rect 57092 8132 57096 8188
rect 57032 8128 57096 8132
rect 57112 8188 57176 8192
rect 57112 8132 57116 8188
rect 57116 8132 57172 8188
rect 57172 8132 57176 8188
rect 57112 8128 57176 8132
rect 57192 8188 57256 8192
rect 57192 8132 57196 8188
rect 57196 8132 57252 8188
rect 57252 8132 57256 8188
rect 57192 8128 57256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 22612 7644 22676 7648
rect 22612 7588 22616 7644
rect 22616 7588 22672 7644
rect 22672 7588 22676 7644
rect 22612 7584 22676 7588
rect 22692 7644 22756 7648
rect 22692 7588 22696 7644
rect 22696 7588 22752 7644
rect 22752 7588 22756 7644
rect 22692 7584 22756 7588
rect 22772 7644 22836 7648
rect 22772 7588 22776 7644
rect 22776 7588 22832 7644
rect 22832 7588 22836 7644
rect 22772 7584 22836 7588
rect 22852 7644 22916 7648
rect 22852 7588 22856 7644
rect 22856 7588 22912 7644
rect 22912 7588 22916 7644
rect 22852 7584 22916 7588
rect 27612 7644 27676 7648
rect 27612 7588 27616 7644
rect 27616 7588 27672 7644
rect 27672 7588 27676 7644
rect 27612 7584 27676 7588
rect 27692 7644 27756 7648
rect 27692 7588 27696 7644
rect 27696 7588 27752 7644
rect 27752 7588 27756 7644
rect 27692 7584 27756 7588
rect 27772 7644 27836 7648
rect 27772 7588 27776 7644
rect 27776 7588 27832 7644
rect 27832 7588 27836 7644
rect 27772 7584 27836 7588
rect 27852 7644 27916 7648
rect 27852 7588 27856 7644
rect 27856 7588 27912 7644
rect 27912 7588 27916 7644
rect 27852 7584 27916 7588
rect 32612 7644 32676 7648
rect 32612 7588 32616 7644
rect 32616 7588 32672 7644
rect 32672 7588 32676 7644
rect 32612 7584 32676 7588
rect 32692 7644 32756 7648
rect 32692 7588 32696 7644
rect 32696 7588 32752 7644
rect 32752 7588 32756 7644
rect 32692 7584 32756 7588
rect 32772 7644 32836 7648
rect 32772 7588 32776 7644
rect 32776 7588 32832 7644
rect 32832 7588 32836 7644
rect 32772 7584 32836 7588
rect 32852 7644 32916 7648
rect 32852 7588 32856 7644
rect 32856 7588 32912 7644
rect 32912 7588 32916 7644
rect 32852 7584 32916 7588
rect 37612 7644 37676 7648
rect 37612 7588 37616 7644
rect 37616 7588 37672 7644
rect 37672 7588 37676 7644
rect 37612 7584 37676 7588
rect 37692 7644 37756 7648
rect 37692 7588 37696 7644
rect 37696 7588 37752 7644
rect 37752 7588 37756 7644
rect 37692 7584 37756 7588
rect 37772 7644 37836 7648
rect 37772 7588 37776 7644
rect 37776 7588 37832 7644
rect 37832 7588 37836 7644
rect 37772 7584 37836 7588
rect 37852 7644 37916 7648
rect 37852 7588 37856 7644
rect 37856 7588 37912 7644
rect 37912 7588 37916 7644
rect 37852 7584 37916 7588
rect 42612 7644 42676 7648
rect 42612 7588 42616 7644
rect 42616 7588 42672 7644
rect 42672 7588 42676 7644
rect 42612 7584 42676 7588
rect 42692 7644 42756 7648
rect 42692 7588 42696 7644
rect 42696 7588 42752 7644
rect 42752 7588 42756 7644
rect 42692 7584 42756 7588
rect 42772 7644 42836 7648
rect 42772 7588 42776 7644
rect 42776 7588 42832 7644
rect 42832 7588 42836 7644
rect 42772 7584 42836 7588
rect 42852 7644 42916 7648
rect 42852 7588 42856 7644
rect 42856 7588 42912 7644
rect 42912 7588 42916 7644
rect 42852 7584 42916 7588
rect 47612 7644 47676 7648
rect 47612 7588 47616 7644
rect 47616 7588 47672 7644
rect 47672 7588 47676 7644
rect 47612 7584 47676 7588
rect 47692 7644 47756 7648
rect 47692 7588 47696 7644
rect 47696 7588 47752 7644
rect 47752 7588 47756 7644
rect 47692 7584 47756 7588
rect 47772 7644 47836 7648
rect 47772 7588 47776 7644
rect 47776 7588 47832 7644
rect 47832 7588 47836 7644
rect 47772 7584 47836 7588
rect 47852 7644 47916 7648
rect 47852 7588 47856 7644
rect 47856 7588 47912 7644
rect 47912 7588 47916 7644
rect 47852 7584 47916 7588
rect 52612 7644 52676 7648
rect 52612 7588 52616 7644
rect 52616 7588 52672 7644
rect 52672 7588 52676 7644
rect 52612 7584 52676 7588
rect 52692 7644 52756 7648
rect 52692 7588 52696 7644
rect 52696 7588 52752 7644
rect 52752 7588 52756 7644
rect 52692 7584 52756 7588
rect 52772 7644 52836 7648
rect 52772 7588 52776 7644
rect 52776 7588 52832 7644
rect 52832 7588 52836 7644
rect 52772 7584 52836 7588
rect 52852 7644 52916 7648
rect 52852 7588 52856 7644
rect 52856 7588 52912 7644
rect 52912 7588 52916 7644
rect 52852 7584 52916 7588
rect 57612 7644 57676 7648
rect 57612 7588 57616 7644
rect 57616 7588 57672 7644
rect 57672 7588 57676 7644
rect 57612 7584 57676 7588
rect 57692 7644 57756 7648
rect 57692 7588 57696 7644
rect 57696 7588 57752 7644
rect 57752 7588 57756 7644
rect 57692 7584 57756 7588
rect 57772 7644 57836 7648
rect 57772 7588 57776 7644
rect 57776 7588 57832 7644
rect 57832 7588 57836 7644
rect 57772 7584 57836 7588
rect 57852 7644 57916 7648
rect 57852 7588 57856 7644
rect 57856 7588 57912 7644
rect 57912 7588 57916 7644
rect 57852 7584 57916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 21952 7100 22016 7104
rect 21952 7044 21956 7100
rect 21956 7044 22012 7100
rect 22012 7044 22016 7100
rect 21952 7040 22016 7044
rect 22032 7100 22096 7104
rect 22032 7044 22036 7100
rect 22036 7044 22092 7100
rect 22092 7044 22096 7100
rect 22032 7040 22096 7044
rect 22112 7100 22176 7104
rect 22112 7044 22116 7100
rect 22116 7044 22172 7100
rect 22172 7044 22176 7100
rect 22112 7040 22176 7044
rect 22192 7100 22256 7104
rect 22192 7044 22196 7100
rect 22196 7044 22252 7100
rect 22252 7044 22256 7100
rect 22192 7040 22256 7044
rect 26952 7100 27016 7104
rect 26952 7044 26956 7100
rect 26956 7044 27012 7100
rect 27012 7044 27016 7100
rect 26952 7040 27016 7044
rect 27032 7100 27096 7104
rect 27032 7044 27036 7100
rect 27036 7044 27092 7100
rect 27092 7044 27096 7100
rect 27032 7040 27096 7044
rect 27112 7100 27176 7104
rect 27112 7044 27116 7100
rect 27116 7044 27172 7100
rect 27172 7044 27176 7100
rect 27112 7040 27176 7044
rect 27192 7100 27256 7104
rect 27192 7044 27196 7100
rect 27196 7044 27252 7100
rect 27252 7044 27256 7100
rect 27192 7040 27256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 36952 7100 37016 7104
rect 36952 7044 36956 7100
rect 36956 7044 37012 7100
rect 37012 7044 37016 7100
rect 36952 7040 37016 7044
rect 37032 7100 37096 7104
rect 37032 7044 37036 7100
rect 37036 7044 37092 7100
rect 37092 7044 37096 7100
rect 37032 7040 37096 7044
rect 37112 7100 37176 7104
rect 37112 7044 37116 7100
rect 37116 7044 37172 7100
rect 37172 7044 37176 7100
rect 37112 7040 37176 7044
rect 37192 7100 37256 7104
rect 37192 7044 37196 7100
rect 37196 7044 37252 7100
rect 37252 7044 37256 7100
rect 37192 7040 37256 7044
rect 41952 7100 42016 7104
rect 41952 7044 41956 7100
rect 41956 7044 42012 7100
rect 42012 7044 42016 7100
rect 41952 7040 42016 7044
rect 42032 7100 42096 7104
rect 42032 7044 42036 7100
rect 42036 7044 42092 7100
rect 42092 7044 42096 7100
rect 42032 7040 42096 7044
rect 42112 7100 42176 7104
rect 42112 7044 42116 7100
rect 42116 7044 42172 7100
rect 42172 7044 42176 7100
rect 42112 7040 42176 7044
rect 42192 7100 42256 7104
rect 42192 7044 42196 7100
rect 42196 7044 42252 7100
rect 42252 7044 42256 7100
rect 42192 7040 42256 7044
rect 46952 7100 47016 7104
rect 46952 7044 46956 7100
rect 46956 7044 47012 7100
rect 47012 7044 47016 7100
rect 46952 7040 47016 7044
rect 47032 7100 47096 7104
rect 47032 7044 47036 7100
rect 47036 7044 47092 7100
rect 47092 7044 47096 7100
rect 47032 7040 47096 7044
rect 47112 7100 47176 7104
rect 47112 7044 47116 7100
rect 47116 7044 47172 7100
rect 47172 7044 47176 7100
rect 47112 7040 47176 7044
rect 47192 7100 47256 7104
rect 47192 7044 47196 7100
rect 47196 7044 47252 7100
rect 47252 7044 47256 7100
rect 47192 7040 47256 7044
rect 51952 7100 52016 7104
rect 51952 7044 51956 7100
rect 51956 7044 52012 7100
rect 52012 7044 52016 7100
rect 51952 7040 52016 7044
rect 52032 7100 52096 7104
rect 52032 7044 52036 7100
rect 52036 7044 52092 7100
rect 52092 7044 52096 7100
rect 52032 7040 52096 7044
rect 52112 7100 52176 7104
rect 52112 7044 52116 7100
rect 52116 7044 52172 7100
rect 52172 7044 52176 7100
rect 52112 7040 52176 7044
rect 52192 7100 52256 7104
rect 52192 7044 52196 7100
rect 52196 7044 52252 7100
rect 52252 7044 52256 7100
rect 52192 7040 52256 7044
rect 56952 7100 57016 7104
rect 56952 7044 56956 7100
rect 56956 7044 57012 7100
rect 57012 7044 57016 7100
rect 56952 7040 57016 7044
rect 57032 7100 57096 7104
rect 57032 7044 57036 7100
rect 57036 7044 57092 7100
rect 57092 7044 57096 7100
rect 57032 7040 57096 7044
rect 57112 7100 57176 7104
rect 57112 7044 57116 7100
rect 57116 7044 57172 7100
rect 57172 7044 57176 7100
rect 57112 7040 57176 7044
rect 57192 7100 57256 7104
rect 57192 7044 57196 7100
rect 57196 7044 57252 7100
rect 57252 7044 57256 7100
rect 57192 7040 57256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 22612 6556 22676 6560
rect 22612 6500 22616 6556
rect 22616 6500 22672 6556
rect 22672 6500 22676 6556
rect 22612 6496 22676 6500
rect 22692 6556 22756 6560
rect 22692 6500 22696 6556
rect 22696 6500 22752 6556
rect 22752 6500 22756 6556
rect 22692 6496 22756 6500
rect 22772 6556 22836 6560
rect 22772 6500 22776 6556
rect 22776 6500 22832 6556
rect 22832 6500 22836 6556
rect 22772 6496 22836 6500
rect 22852 6556 22916 6560
rect 22852 6500 22856 6556
rect 22856 6500 22912 6556
rect 22912 6500 22916 6556
rect 22852 6496 22916 6500
rect 27612 6556 27676 6560
rect 27612 6500 27616 6556
rect 27616 6500 27672 6556
rect 27672 6500 27676 6556
rect 27612 6496 27676 6500
rect 27692 6556 27756 6560
rect 27692 6500 27696 6556
rect 27696 6500 27752 6556
rect 27752 6500 27756 6556
rect 27692 6496 27756 6500
rect 27772 6556 27836 6560
rect 27772 6500 27776 6556
rect 27776 6500 27832 6556
rect 27832 6500 27836 6556
rect 27772 6496 27836 6500
rect 27852 6556 27916 6560
rect 27852 6500 27856 6556
rect 27856 6500 27912 6556
rect 27912 6500 27916 6556
rect 27852 6496 27916 6500
rect 32612 6556 32676 6560
rect 32612 6500 32616 6556
rect 32616 6500 32672 6556
rect 32672 6500 32676 6556
rect 32612 6496 32676 6500
rect 32692 6556 32756 6560
rect 32692 6500 32696 6556
rect 32696 6500 32752 6556
rect 32752 6500 32756 6556
rect 32692 6496 32756 6500
rect 32772 6556 32836 6560
rect 32772 6500 32776 6556
rect 32776 6500 32832 6556
rect 32832 6500 32836 6556
rect 32772 6496 32836 6500
rect 32852 6556 32916 6560
rect 32852 6500 32856 6556
rect 32856 6500 32912 6556
rect 32912 6500 32916 6556
rect 32852 6496 32916 6500
rect 37612 6556 37676 6560
rect 37612 6500 37616 6556
rect 37616 6500 37672 6556
rect 37672 6500 37676 6556
rect 37612 6496 37676 6500
rect 37692 6556 37756 6560
rect 37692 6500 37696 6556
rect 37696 6500 37752 6556
rect 37752 6500 37756 6556
rect 37692 6496 37756 6500
rect 37772 6556 37836 6560
rect 37772 6500 37776 6556
rect 37776 6500 37832 6556
rect 37832 6500 37836 6556
rect 37772 6496 37836 6500
rect 37852 6556 37916 6560
rect 37852 6500 37856 6556
rect 37856 6500 37912 6556
rect 37912 6500 37916 6556
rect 37852 6496 37916 6500
rect 42612 6556 42676 6560
rect 42612 6500 42616 6556
rect 42616 6500 42672 6556
rect 42672 6500 42676 6556
rect 42612 6496 42676 6500
rect 42692 6556 42756 6560
rect 42692 6500 42696 6556
rect 42696 6500 42752 6556
rect 42752 6500 42756 6556
rect 42692 6496 42756 6500
rect 42772 6556 42836 6560
rect 42772 6500 42776 6556
rect 42776 6500 42832 6556
rect 42832 6500 42836 6556
rect 42772 6496 42836 6500
rect 42852 6556 42916 6560
rect 42852 6500 42856 6556
rect 42856 6500 42912 6556
rect 42912 6500 42916 6556
rect 42852 6496 42916 6500
rect 47612 6556 47676 6560
rect 47612 6500 47616 6556
rect 47616 6500 47672 6556
rect 47672 6500 47676 6556
rect 47612 6496 47676 6500
rect 47692 6556 47756 6560
rect 47692 6500 47696 6556
rect 47696 6500 47752 6556
rect 47752 6500 47756 6556
rect 47692 6496 47756 6500
rect 47772 6556 47836 6560
rect 47772 6500 47776 6556
rect 47776 6500 47832 6556
rect 47832 6500 47836 6556
rect 47772 6496 47836 6500
rect 47852 6556 47916 6560
rect 47852 6500 47856 6556
rect 47856 6500 47912 6556
rect 47912 6500 47916 6556
rect 47852 6496 47916 6500
rect 52612 6556 52676 6560
rect 52612 6500 52616 6556
rect 52616 6500 52672 6556
rect 52672 6500 52676 6556
rect 52612 6496 52676 6500
rect 52692 6556 52756 6560
rect 52692 6500 52696 6556
rect 52696 6500 52752 6556
rect 52752 6500 52756 6556
rect 52692 6496 52756 6500
rect 52772 6556 52836 6560
rect 52772 6500 52776 6556
rect 52776 6500 52832 6556
rect 52832 6500 52836 6556
rect 52772 6496 52836 6500
rect 52852 6556 52916 6560
rect 52852 6500 52856 6556
rect 52856 6500 52912 6556
rect 52912 6500 52916 6556
rect 52852 6496 52916 6500
rect 57612 6556 57676 6560
rect 57612 6500 57616 6556
rect 57616 6500 57672 6556
rect 57672 6500 57676 6556
rect 57612 6496 57676 6500
rect 57692 6556 57756 6560
rect 57692 6500 57696 6556
rect 57696 6500 57752 6556
rect 57752 6500 57756 6556
rect 57692 6496 57756 6500
rect 57772 6556 57836 6560
rect 57772 6500 57776 6556
rect 57776 6500 57832 6556
rect 57832 6500 57836 6556
rect 57772 6496 57836 6500
rect 57852 6556 57916 6560
rect 57852 6500 57856 6556
rect 57856 6500 57912 6556
rect 57912 6500 57916 6556
rect 57852 6496 57916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 21952 6012 22016 6016
rect 21952 5956 21956 6012
rect 21956 5956 22012 6012
rect 22012 5956 22016 6012
rect 21952 5952 22016 5956
rect 22032 6012 22096 6016
rect 22032 5956 22036 6012
rect 22036 5956 22092 6012
rect 22092 5956 22096 6012
rect 22032 5952 22096 5956
rect 22112 6012 22176 6016
rect 22112 5956 22116 6012
rect 22116 5956 22172 6012
rect 22172 5956 22176 6012
rect 22112 5952 22176 5956
rect 22192 6012 22256 6016
rect 22192 5956 22196 6012
rect 22196 5956 22252 6012
rect 22252 5956 22256 6012
rect 22192 5952 22256 5956
rect 26952 6012 27016 6016
rect 26952 5956 26956 6012
rect 26956 5956 27012 6012
rect 27012 5956 27016 6012
rect 26952 5952 27016 5956
rect 27032 6012 27096 6016
rect 27032 5956 27036 6012
rect 27036 5956 27092 6012
rect 27092 5956 27096 6012
rect 27032 5952 27096 5956
rect 27112 6012 27176 6016
rect 27112 5956 27116 6012
rect 27116 5956 27172 6012
rect 27172 5956 27176 6012
rect 27112 5952 27176 5956
rect 27192 6012 27256 6016
rect 27192 5956 27196 6012
rect 27196 5956 27252 6012
rect 27252 5956 27256 6012
rect 27192 5952 27256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 36952 6012 37016 6016
rect 36952 5956 36956 6012
rect 36956 5956 37012 6012
rect 37012 5956 37016 6012
rect 36952 5952 37016 5956
rect 37032 6012 37096 6016
rect 37032 5956 37036 6012
rect 37036 5956 37092 6012
rect 37092 5956 37096 6012
rect 37032 5952 37096 5956
rect 37112 6012 37176 6016
rect 37112 5956 37116 6012
rect 37116 5956 37172 6012
rect 37172 5956 37176 6012
rect 37112 5952 37176 5956
rect 37192 6012 37256 6016
rect 37192 5956 37196 6012
rect 37196 5956 37252 6012
rect 37252 5956 37256 6012
rect 37192 5952 37256 5956
rect 41952 6012 42016 6016
rect 41952 5956 41956 6012
rect 41956 5956 42012 6012
rect 42012 5956 42016 6012
rect 41952 5952 42016 5956
rect 42032 6012 42096 6016
rect 42032 5956 42036 6012
rect 42036 5956 42092 6012
rect 42092 5956 42096 6012
rect 42032 5952 42096 5956
rect 42112 6012 42176 6016
rect 42112 5956 42116 6012
rect 42116 5956 42172 6012
rect 42172 5956 42176 6012
rect 42112 5952 42176 5956
rect 42192 6012 42256 6016
rect 42192 5956 42196 6012
rect 42196 5956 42252 6012
rect 42252 5956 42256 6012
rect 42192 5952 42256 5956
rect 46952 6012 47016 6016
rect 46952 5956 46956 6012
rect 46956 5956 47012 6012
rect 47012 5956 47016 6012
rect 46952 5952 47016 5956
rect 47032 6012 47096 6016
rect 47032 5956 47036 6012
rect 47036 5956 47092 6012
rect 47092 5956 47096 6012
rect 47032 5952 47096 5956
rect 47112 6012 47176 6016
rect 47112 5956 47116 6012
rect 47116 5956 47172 6012
rect 47172 5956 47176 6012
rect 47112 5952 47176 5956
rect 47192 6012 47256 6016
rect 47192 5956 47196 6012
rect 47196 5956 47252 6012
rect 47252 5956 47256 6012
rect 47192 5952 47256 5956
rect 51952 6012 52016 6016
rect 51952 5956 51956 6012
rect 51956 5956 52012 6012
rect 52012 5956 52016 6012
rect 51952 5952 52016 5956
rect 52032 6012 52096 6016
rect 52032 5956 52036 6012
rect 52036 5956 52092 6012
rect 52092 5956 52096 6012
rect 52032 5952 52096 5956
rect 52112 6012 52176 6016
rect 52112 5956 52116 6012
rect 52116 5956 52172 6012
rect 52172 5956 52176 6012
rect 52112 5952 52176 5956
rect 52192 6012 52256 6016
rect 52192 5956 52196 6012
rect 52196 5956 52252 6012
rect 52252 5956 52256 6012
rect 52192 5952 52256 5956
rect 56952 6012 57016 6016
rect 56952 5956 56956 6012
rect 56956 5956 57012 6012
rect 57012 5956 57016 6012
rect 56952 5952 57016 5956
rect 57032 6012 57096 6016
rect 57032 5956 57036 6012
rect 57036 5956 57092 6012
rect 57092 5956 57096 6012
rect 57032 5952 57096 5956
rect 57112 6012 57176 6016
rect 57112 5956 57116 6012
rect 57116 5956 57172 6012
rect 57172 5956 57176 6012
rect 57112 5952 57176 5956
rect 57192 6012 57256 6016
rect 57192 5956 57196 6012
rect 57196 5956 57252 6012
rect 57252 5956 57256 6012
rect 57192 5952 57256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 22612 5468 22676 5472
rect 22612 5412 22616 5468
rect 22616 5412 22672 5468
rect 22672 5412 22676 5468
rect 22612 5408 22676 5412
rect 22692 5468 22756 5472
rect 22692 5412 22696 5468
rect 22696 5412 22752 5468
rect 22752 5412 22756 5468
rect 22692 5408 22756 5412
rect 22772 5468 22836 5472
rect 22772 5412 22776 5468
rect 22776 5412 22832 5468
rect 22832 5412 22836 5468
rect 22772 5408 22836 5412
rect 22852 5468 22916 5472
rect 22852 5412 22856 5468
rect 22856 5412 22912 5468
rect 22912 5412 22916 5468
rect 22852 5408 22916 5412
rect 27612 5468 27676 5472
rect 27612 5412 27616 5468
rect 27616 5412 27672 5468
rect 27672 5412 27676 5468
rect 27612 5408 27676 5412
rect 27692 5468 27756 5472
rect 27692 5412 27696 5468
rect 27696 5412 27752 5468
rect 27752 5412 27756 5468
rect 27692 5408 27756 5412
rect 27772 5468 27836 5472
rect 27772 5412 27776 5468
rect 27776 5412 27832 5468
rect 27832 5412 27836 5468
rect 27772 5408 27836 5412
rect 27852 5468 27916 5472
rect 27852 5412 27856 5468
rect 27856 5412 27912 5468
rect 27912 5412 27916 5468
rect 27852 5408 27916 5412
rect 32612 5468 32676 5472
rect 32612 5412 32616 5468
rect 32616 5412 32672 5468
rect 32672 5412 32676 5468
rect 32612 5408 32676 5412
rect 32692 5468 32756 5472
rect 32692 5412 32696 5468
rect 32696 5412 32752 5468
rect 32752 5412 32756 5468
rect 32692 5408 32756 5412
rect 32772 5468 32836 5472
rect 32772 5412 32776 5468
rect 32776 5412 32832 5468
rect 32832 5412 32836 5468
rect 32772 5408 32836 5412
rect 32852 5468 32916 5472
rect 32852 5412 32856 5468
rect 32856 5412 32912 5468
rect 32912 5412 32916 5468
rect 32852 5408 32916 5412
rect 37612 5468 37676 5472
rect 37612 5412 37616 5468
rect 37616 5412 37672 5468
rect 37672 5412 37676 5468
rect 37612 5408 37676 5412
rect 37692 5468 37756 5472
rect 37692 5412 37696 5468
rect 37696 5412 37752 5468
rect 37752 5412 37756 5468
rect 37692 5408 37756 5412
rect 37772 5468 37836 5472
rect 37772 5412 37776 5468
rect 37776 5412 37832 5468
rect 37832 5412 37836 5468
rect 37772 5408 37836 5412
rect 37852 5468 37916 5472
rect 37852 5412 37856 5468
rect 37856 5412 37912 5468
rect 37912 5412 37916 5468
rect 37852 5408 37916 5412
rect 42612 5468 42676 5472
rect 42612 5412 42616 5468
rect 42616 5412 42672 5468
rect 42672 5412 42676 5468
rect 42612 5408 42676 5412
rect 42692 5468 42756 5472
rect 42692 5412 42696 5468
rect 42696 5412 42752 5468
rect 42752 5412 42756 5468
rect 42692 5408 42756 5412
rect 42772 5468 42836 5472
rect 42772 5412 42776 5468
rect 42776 5412 42832 5468
rect 42832 5412 42836 5468
rect 42772 5408 42836 5412
rect 42852 5468 42916 5472
rect 42852 5412 42856 5468
rect 42856 5412 42912 5468
rect 42912 5412 42916 5468
rect 42852 5408 42916 5412
rect 47612 5468 47676 5472
rect 47612 5412 47616 5468
rect 47616 5412 47672 5468
rect 47672 5412 47676 5468
rect 47612 5408 47676 5412
rect 47692 5468 47756 5472
rect 47692 5412 47696 5468
rect 47696 5412 47752 5468
rect 47752 5412 47756 5468
rect 47692 5408 47756 5412
rect 47772 5468 47836 5472
rect 47772 5412 47776 5468
rect 47776 5412 47832 5468
rect 47832 5412 47836 5468
rect 47772 5408 47836 5412
rect 47852 5468 47916 5472
rect 47852 5412 47856 5468
rect 47856 5412 47912 5468
rect 47912 5412 47916 5468
rect 47852 5408 47916 5412
rect 52612 5468 52676 5472
rect 52612 5412 52616 5468
rect 52616 5412 52672 5468
rect 52672 5412 52676 5468
rect 52612 5408 52676 5412
rect 52692 5468 52756 5472
rect 52692 5412 52696 5468
rect 52696 5412 52752 5468
rect 52752 5412 52756 5468
rect 52692 5408 52756 5412
rect 52772 5468 52836 5472
rect 52772 5412 52776 5468
rect 52776 5412 52832 5468
rect 52832 5412 52836 5468
rect 52772 5408 52836 5412
rect 52852 5468 52916 5472
rect 52852 5412 52856 5468
rect 52856 5412 52912 5468
rect 52912 5412 52916 5468
rect 52852 5408 52916 5412
rect 57612 5468 57676 5472
rect 57612 5412 57616 5468
rect 57616 5412 57672 5468
rect 57672 5412 57676 5468
rect 57612 5408 57676 5412
rect 57692 5468 57756 5472
rect 57692 5412 57696 5468
rect 57696 5412 57752 5468
rect 57752 5412 57756 5468
rect 57692 5408 57756 5412
rect 57772 5468 57836 5472
rect 57772 5412 57776 5468
rect 57776 5412 57832 5468
rect 57832 5412 57836 5468
rect 57772 5408 57836 5412
rect 57852 5468 57916 5472
rect 57852 5412 57856 5468
rect 57856 5412 57912 5468
rect 57912 5412 57916 5468
rect 57852 5408 57916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 21952 4924 22016 4928
rect 21952 4868 21956 4924
rect 21956 4868 22012 4924
rect 22012 4868 22016 4924
rect 21952 4864 22016 4868
rect 22032 4924 22096 4928
rect 22032 4868 22036 4924
rect 22036 4868 22092 4924
rect 22092 4868 22096 4924
rect 22032 4864 22096 4868
rect 22112 4924 22176 4928
rect 22112 4868 22116 4924
rect 22116 4868 22172 4924
rect 22172 4868 22176 4924
rect 22112 4864 22176 4868
rect 22192 4924 22256 4928
rect 22192 4868 22196 4924
rect 22196 4868 22252 4924
rect 22252 4868 22256 4924
rect 22192 4864 22256 4868
rect 26952 4924 27016 4928
rect 26952 4868 26956 4924
rect 26956 4868 27012 4924
rect 27012 4868 27016 4924
rect 26952 4864 27016 4868
rect 27032 4924 27096 4928
rect 27032 4868 27036 4924
rect 27036 4868 27092 4924
rect 27092 4868 27096 4924
rect 27032 4864 27096 4868
rect 27112 4924 27176 4928
rect 27112 4868 27116 4924
rect 27116 4868 27172 4924
rect 27172 4868 27176 4924
rect 27112 4864 27176 4868
rect 27192 4924 27256 4928
rect 27192 4868 27196 4924
rect 27196 4868 27252 4924
rect 27252 4868 27256 4924
rect 27192 4864 27256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 36952 4924 37016 4928
rect 36952 4868 36956 4924
rect 36956 4868 37012 4924
rect 37012 4868 37016 4924
rect 36952 4864 37016 4868
rect 37032 4924 37096 4928
rect 37032 4868 37036 4924
rect 37036 4868 37092 4924
rect 37092 4868 37096 4924
rect 37032 4864 37096 4868
rect 37112 4924 37176 4928
rect 37112 4868 37116 4924
rect 37116 4868 37172 4924
rect 37172 4868 37176 4924
rect 37112 4864 37176 4868
rect 37192 4924 37256 4928
rect 37192 4868 37196 4924
rect 37196 4868 37252 4924
rect 37252 4868 37256 4924
rect 37192 4864 37256 4868
rect 41952 4924 42016 4928
rect 41952 4868 41956 4924
rect 41956 4868 42012 4924
rect 42012 4868 42016 4924
rect 41952 4864 42016 4868
rect 42032 4924 42096 4928
rect 42032 4868 42036 4924
rect 42036 4868 42092 4924
rect 42092 4868 42096 4924
rect 42032 4864 42096 4868
rect 42112 4924 42176 4928
rect 42112 4868 42116 4924
rect 42116 4868 42172 4924
rect 42172 4868 42176 4924
rect 42112 4864 42176 4868
rect 42192 4924 42256 4928
rect 42192 4868 42196 4924
rect 42196 4868 42252 4924
rect 42252 4868 42256 4924
rect 42192 4864 42256 4868
rect 46952 4924 47016 4928
rect 46952 4868 46956 4924
rect 46956 4868 47012 4924
rect 47012 4868 47016 4924
rect 46952 4864 47016 4868
rect 47032 4924 47096 4928
rect 47032 4868 47036 4924
rect 47036 4868 47092 4924
rect 47092 4868 47096 4924
rect 47032 4864 47096 4868
rect 47112 4924 47176 4928
rect 47112 4868 47116 4924
rect 47116 4868 47172 4924
rect 47172 4868 47176 4924
rect 47112 4864 47176 4868
rect 47192 4924 47256 4928
rect 47192 4868 47196 4924
rect 47196 4868 47252 4924
rect 47252 4868 47256 4924
rect 47192 4864 47256 4868
rect 51952 4924 52016 4928
rect 51952 4868 51956 4924
rect 51956 4868 52012 4924
rect 52012 4868 52016 4924
rect 51952 4864 52016 4868
rect 52032 4924 52096 4928
rect 52032 4868 52036 4924
rect 52036 4868 52092 4924
rect 52092 4868 52096 4924
rect 52032 4864 52096 4868
rect 52112 4924 52176 4928
rect 52112 4868 52116 4924
rect 52116 4868 52172 4924
rect 52172 4868 52176 4924
rect 52112 4864 52176 4868
rect 52192 4924 52256 4928
rect 52192 4868 52196 4924
rect 52196 4868 52252 4924
rect 52252 4868 52256 4924
rect 52192 4864 52256 4868
rect 56952 4924 57016 4928
rect 56952 4868 56956 4924
rect 56956 4868 57012 4924
rect 57012 4868 57016 4924
rect 56952 4864 57016 4868
rect 57032 4924 57096 4928
rect 57032 4868 57036 4924
rect 57036 4868 57092 4924
rect 57092 4868 57096 4924
rect 57032 4864 57096 4868
rect 57112 4924 57176 4928
rect 57112 4868 57116 4924
rect 57116 4868 57172 4924
rect 57172 4868 57176 4924
rect 57112 4864 57176 4868
rect 57192 4924 57256 4928
rect 57192 4868 57196 4924
rect 57196 4868 57252 4924
rect 57252 4868 57256 4924
rect 57192 4864 57256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 22612 4380 22676 4384
rect 22612 4324 22616 4380
rect 22616 4324 22672 4380
rect 22672 4324 22676 4380
rect 22612 4320 22676 4324
rect 22692 4380 22756 4384
rect 22692 4324 22696 4380
rect 22696 4324 22752 4380
rect 22752 4324 22756 4380
rect 22692 4320 22756 4324
rect 22772 4380 22836 4384
rect 22772 4324 22776 4380
rect 22776 4324 22832 4380
rect 22832 4324 22836 4380
rect 22772 4320 22836 4324
rect 22852 4380 22916 4384
rect 22852 4324 22856 4380
rect 22856 4324 22912 4380
rect 22912 4324 22916 4380
rect 22852 4320 22916 4324
rect 27612 4380 27676 4384
rect 27612 4324 27616 4380
rect 27616 4324 27672 4380
rect 27672 4324 27676 4380
rect 27612 4320 27676 4324
rect 27692 4380 27756 4384
rect 27692 4324 27696 4380
rect 27696 4324 27752 4380
rect 27752 4324 27756 4380
rect 27692 4320 27756 4324
rect 27772 4380 27836 4384
rect 27772 4324 27776 4380
rect 27776 4324 27832 4380
rect 27832 4324 27836 4380
rect 27772 4320 27836 4324
rect 27852 4380 27916 4384
rect 27852 4324 27856 4380
rect 27856 4324 27912 4380
rect 27912 4324 27916 4380
rect 27852 4320 27916 4324
rect 32612 4380 32676 4384
rect 32612 4324 32616 4380
rect 32616 4324 32672 4380
rect 32672 4324 32676 4380
rect 32612 4320 32676 4324
rect 32692 4380 32756 4384
rect 32692 4324 32696 4380
rect 32696 4324 32752 4380
rect 32752 4324 32756 4380
rect 32692 4320 32756 4324
rect 32772 4380 32836 4384
rect 32772 4324 32776 4380
rect 32776 4324 32832 4380
rect 32832 4324 32836 4380
rect 32772 4320 32836 4324
rect 32852 4380 32916 4384
rect 32852 4324 32856 4380
rect 32856 4324 32912 4380
rect 32912 4324 32916 4380
rect 32852 4320 32916 4324
rect 37612 4380 37676 4384
rect 37612 4324 37616 4380
rect 37616 4324 37672 4380
rect 37672 4324 37676 4380
rect 37612 4320 37676 4324
rect 37692 4380 37756 4384
rect 37692 4324 37696 4380
rect 37696 4324 37752 4380
rect 37752 4324 37756 4380
rect 37692 4320 37756 4324
rect 37772 4380 37836 4384
rect 37772 4324 37776 4380
rect 37776 4324 37832 4380
rect 37832 4324 37836 4380
rect 37772 4320 37836 4324
rect 37852 4380 37916 4384
rect 37852 4324 37856 4380
rect 37856 4324 37912 4380
rect 37912 4324 37916 4380
rect 37852 4320 37916 4324
rect 42612 4380 42676 4384
rect 42612 4324 42616 4380
rect 42616 4324 42672 4380
rect 42672 4324 42676 4380
rect 42612 4320 42676 4324
rect 42692 4380 42756 4384
rect 42692 4324 42696 4380
rect 42696 4324 42752 4380
rect 42752 4324 42756 4380
rect 42692 4320 42756 4324
rect 42772 4380 42836 4384
rect 42772 4324 42776 4380
rect 42776 4324 42832 4380
rect 42832 4324 42836 4380
rect 42772 4320 42836 4324
rect 42852 4380 42916 4384
rect 42852 4324 42856 4380
rect 42856 4324 42912 4380
rect 42912 4324 42916 4380
rect 42852 4320 42916 4324
rect 47612 4380 47676 4384
rect 47612 4324 47616 4380
rect 47616 4324 47672 4380
rect 47672 4324 47676 4380
rect 47612 4320 47676 4324
rect 47692 4380 47756 4384
rect 47692 4324 47696 4380
rect 47696 4324 47752 4380
rect 47752 4324 47756 4380
rect 47692 4320 47756 4324
rect 47772 4380 47836 4384
rect 47772 4324 47776 4380
rect 47776 4324 47832 4380
rect 47832 4324 47836 4380
rect 47772 4320 47836 4324
rect 47852 4380 47916 4384
rect 47852 4324 47856 4380
rect 47856 4324 47912 4380
rect 47912 4324 47916 4380
rect 47852 4320 47916 4324
rect 52612 4380 52676 4384
rect 52612 4324 52616 4380
rect 52616 4324 52672 4380
rect 52672 4324 52676 4380
rect 52612 4320 52676 4324
rect 52692 4380 52756 4384
rect 52692 4324 52696 4380
rect 52696 4324 52752 4380
rect 52752 4324 52756 4380
rect 52692 4320 52756 4324
rect 52772 4380 52836 4384
rect 52772 4324 52776 4380
rect 52776 4324 52832 4380
rect 52832 4324 52836 4380
rect 52772 4320 52836 4324
rect 52852 4380 52916 4384
rect 52852 4324 52856 4380
rect 52856 4324 52912 4380
rect 52912 4324 52916 4380
rect 52852 4320 52916 4324
rect 57612 4380 57676 4384
rect 57612 4324 57616 4380
rect 57616 4324 57672 4380
rect 57672 4324 57676 4380
rect 57612 4320 57676 4324
rect 57692 4380 57756 4384
rect 57692 4324 57696 4380
rect 57696 4324 57752 4380
rect 57752 4324 57756 4380
rect 57692 4320 57756 4324
rect 57772 4380 57836 4384
rect 57772 4324 57776 4380
rect 57776 4324 57832 4380
rect 57832 4324 57836 4380
rect 57772 4320 57836 4324
rect 57852 4380 57916 4384
rect 57852 4324 57856 4380
rect 57856 4324 57912 4380
rect 57912 4324 57916 4380
rect 57852 4320 57916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 21952 3836 22016 3840
rect 21952 3780 21956 3836
rect 21956 3780 22012 3836
rect 22012 3780 22016 3836
rect 21952 3776 22016 3780
rect 22032 3836 22096 3840
rect 22032 3780 22036 3836
rect 22036 3780 22092 3836
rect 22092 3780 22096 3836
rect 22032 3776 22096 3780
rect 22112 3836 22176 3840
rect 22112 3780 22116 3836
rect 22116 3780 22172 3836
rect 22172 3780 22176 3836
rect 22112 3776 22176 3780
rect 22192 3836 22256 3840
rect 22192 3780 22196 3836
rect 22196 3780 22252 3836
rect 22252 3780 22256 3836
rect 22192 3776 22256 3780
rect 26952 3836 27016 3840
rect 26952 3780 26956 3836
rect 26956 3780 27012 3836
rect 27012 3780 27016 3836
rect 26952 3776 27016 3780
rect 27032 3836 27096 3840
rect 27032 3780 27036 3836
rect 27036 3780 27092 3836
rect 27092 3780 27096 3836
rect 27032 3776 27096 3780
rect 27112 3836 27176 3840
rect 27112 3780 27116 3836
rect 27116 3780 27172 3836
rect 27172 3780 27176 3836
rect 27112 3776 27176 3780
rect 27192 3836 27256 3840
rect 27192 3780 27196 3836
rect 27196 3780 27252 3836
rect 27252 3780 27256 3836
rect 27192 3776 27256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 36952 3836 37016 3840
rect 36952 3780 36956 3836
rect 36956 3780 37012 3836
rect 37012 3780 37016 3836
rect 36952 3776 37016 3780
rect 37032 3836 37096 3840
rect 37032 3780 37036 3836
rect 37036 3780 37092 3836
rect 37092 3780 37096 3836
rect 37032 3776 37096 3780
rect 37112 3836 37176 3840
rect 37112 3780 37116 3836
rect 37116 3780 37172 3836
rect 37172 3780 37176 3836
rect 37112 3776 37176 3780
rect 37192 3836 37256 3840
rect 37192 3780 37196 3836
rect 37196 3780 37252 3836
rect 37252 3780 37256 3836
rect 37192 3776 37256 3780
rect 41952 3836 42016 3840
rect 41952 3780 41956 3836
rect 41956 3780 42012 3836
rect 42012 3780 42016 3836
rect 41952 3776 42016 3780
rect 42032 3836 42096 3840
rect 42032 3780 42036 3836
rect 42036 3780 42092 3836
rect 42092 3780 42096 3836
rect 42032 3776 42096 3780
rect 42112 3836 42176 3840
rect 42112 3780 42116 3836
rect 42116 3780 42172 3836
rect 42172 3780 42176 3836
rect 42112 3776 42176 3780
rect 42192 3836 42256 3840
rect 42192 3780 42196 3836
rect 42196 3780 42252 3836
rect 42252 3780 42256 3836
rect 42192 3776 42256 3780
rect 46952 3836 47016 3840
rect 46952 3780 46956 3836
rect 46956 3780 47012 3836
rect 47012 3780 47016 3836
rect 46952 3776 47016 3780
rect 47032 3836 47096 3840
rect 47032 3780 47036 3836
rect 47036 3780 47092 3836
rect 47092 3780 47096 3836
rect 47032 3776 47096 3780
rect 47112 3836 47176 3840
rect 47112 3780 47116 3836
rect 47116 3780 47172 3836
rect 47172 3780 47176 3836
rect 47112 3776 47176 3780
rect 47192 3836 47256 3840
rect 47192 3780 47196 3836
rect 47196 3780 47252 3836
rect 47252 3780 47256 3836
rect 47192 3776 47256 3780
rect 51952 3836 52016 3840
rect 51952 3780 51956 3836
rect 51956 3780 52012 3836
rect 52012 3780 52016 3836
rect 51952 3776 52016 3780
rect 52032 3836 52096 3840
rect 52032 3780 52036 3836
rect 52036 3780 52092 3836
rect 52092 3780 52096 3836
rect 52032 3776 52096 3780
rect 52112 3836 52176 3840
rect 52112 3780 52116 3836
rect 52116 3780 52172 3836
rect 52172 3780 52176 3836
rect 52112 3776 52176 3780
rect 52192 3836 52256 3840
rect 52192 3780 52196 3836
rect 52196 3780 52252 3836
rect 52252 3780 52256 3836
rect 52192 3776 52256 3780
rect 56952 3836 57016 3840
rect 56952 3780 56956 3836
rect 56956 3780 57012 3836
rect 57012 3780 57016 3836
rect 56952 3776 57016 3780
rect 57032 3836 57096 3840
rect 57032 3780 57036 3836
rect 57036 3780 57092 3836
rect 57092 3780 57096 3836
rect 57032 3776 57096 3780
rect 57112 3836 57176 3840
rect 57112 3780 57116 3836
rect 57116 3780 57172 3836
rect 57172 3780 57176 3836
rect 57112 3776 57176 3780
rect 57192 3836 57256 3840
rect 57192 3780 57196 3836
rect 57196 3780 57252 3836
rect 57252 3780 57256 3836
rect 57192 3776 57256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 22612 3292 22676 3296
rect 22612 3236 22616 3292
rect 22616 3236 22672 3292
rect 22672 3236 22676 3292
rect 22612 3232 22676 3236
rect 22692 3292 22756 3296
rect 22692 3236 22696 3292
rect 22696 3236 22752 3292
rect 22752 3236 22756 3292
rect 22692 3232 22756 3236
rect 22772 3292 22836 3296
rect 22772 3236 22776 3292
rect 22776 3236 22832 3292
rect 22832 3236 22836 3292
rect 22772 3232 22836 3236
rect 22852 3292 22916 3296
rect 22852 3236 22856 3292
rect 22856 3236 22912 3292
rect 22912 3236 22916 3292
rect 22852 3232 22916 3236
rect 27612 3292 27676 3296
rect 27612 3236 27616 3292
rect 27616 3236 27672 3292
rect 27672 3236 27676 3292
rect 27612 3232 27676 3236
rect 27692 3292 27756 3296
rect 27692 3236 27696 3292
rect 27696 3236 27752 3292
rect 27752 3236 27756 3292
rect 27692 3232 27756 3236
rect 27772 3292 27836 3296
rect 27772 3236 27776 3292
rect 27776 3236 27832 3292
rect 27832 3236 27836 3292
rect 27772 3232 27836 3236
rect 27852 3292 27916 3296
rect 27852 3236 27856 3292
rect 27856 3236 27912 3292
rect 27912 3236 27916 3292
rect 27852 3232 27916 3236
rect 32612 3292 32676 3296
rect 32612 3236 32616 3292
rect 32616 3236 32672 3292
rect 32672 3236 32676 3292
rect 32612 3232 32676 3236
rect 32692 3292 32756 3296
rect 32692 3236 32696 3292
rect 32696 3236 32752 3292
rect 32752 3236 32756 3292
rect 32692 3232 32756 3236
rect 32772 3292 32836 3296
rect 32772 3236 32776 3292
rect 32776 3236 32832 3292
rect 32832 3236 32836 3292
rect 32772 3232 32836 3236
rect 32852 3292 32916 3296
rect 32852 3236 32856 3292
rect 32856 3236 32912 3292
rect 32912 3236 32916 3292
rect 32852 3232 32916 3236
rect 37612 3292 37676 3296
rect 37612 3236 37616 3292
rect 37616 3236 37672 3292
rect 37672 3236 37676 3292
rect 37612 3232 37676 3236
rect 37692 3292 37756 3296
rect 37692 3236 37696 3292
rect 37696 3236 37752 3292
rect 37752 3236 37756 3292
rect 37692 3232 37756 3236
rect 37772 3292 37836 3296
rect 37772 3236 37776 3292
rect 37776 3236 37832 3292
rect 37832 3236 37836 3292
rect 37772 3232 37836 3236
rect 37852 3292 37916 3296
rect 37852 3236 37856 3292
rect 37856 3236 37912 3292
rect 37912 3236 37916 3292
rect 37852 3232 37916 3236
rect 42612 3292 42676 3296
rect 42612 3236 42616 3292
rect 42616 3236 42672 3292
rect 42672 3236 42676 3292
rect 42612 3232 42676 3236
rect 42692 3292 42756 3296
rect 42692 3236 42696 3292
rect 42696 3236 42752 3292
rect 42752 3236 42756 3292
rect 42692 3232 42756 3236
rect 42772 3292 42836 3296
rect 42772 3236 42776 3292
rect 42776 3236 42832 3292
rect 42832 3236 42836 3292
rect 42772 3232 42836 3236
rect 42852 3292 42916 3296
rect 42852 3236 42856 3292
rect 42856 3236 42912 3292
rect 42912 3236 42916 3292
rect 42852 3232 42916 3236
rect 47612 3292 47676 3296
rect 47612 3236 47616 3292
rect 47616 3236 47672 3292
rect 47672 3236 47676 3292
rect 47612 3232 47676 3236
rect 47692 3292 47756 3296
rect 47692 3236 47696 3292
rect 47696 3236 47752 3292
rect 47752 3236 47756 3292
rect 47692 3232 47756 3236
rect 47772 3292 47836 3296
rect 47772 3236 47776 3292
rect 47776 3236 47832 3292
rect 47832 3236 47836 3292
rect 47772 3232 47836 3236
rect 47852 3292 47916 3296
rect 47852 3236 47856 3292
rect 47856 3236 47912 3292
rect 47912 3236 47916 3292
rect 47852 3232 47916 3236
rect 52612 3292 52676 3296
rect 52612 3236 52616 3292
rect 52616 3236 52672 3292
rect 52672 3236 52676 3292
rect 52612 3232 52676 3236
rect 52692 3292 52756 3296
rect 52692 3236 52696 3292
rect 52696 3236 52752 3292
rect 52752 3236 52756 3292
rect 52692 3232 52756 3236
rect 52772 3292 52836 3296
rect 52772 3236 52776 3292
rect 52776 3236 52832 3292
rect 52832 3236 52836 3292
rect 52772 3232 52836 3236
rect 52852 3292 52916 3296
rect 52852 3236 52856 3292
rect 52856 3236 52912 3292
rect 52912 3236 52916 3292
rect 52852 3232 52916 3236
rect 57612 3292 57676 3296
rect 57612 3236 57616 3292
rect 57616 3236 57672 3292
rect 57672 3236 57676 3292
rect 57612 3232 57676 3236
rect 57692 3292 57756 3296
rect 57692 3236 57696 3292
rect 57696 3236 57752 3292
rect 57752 3236 57756 3292
rect 57692 3232 57756 3236
rect 57772 3292 57836 3296
rect 57772 3236 57776 3292
rect 57776 3236 57832 3292
rect 57832 3236 57836 3292
rect 57772 3232 57836 3236
rect 57852 3292 57916 3296
rect 57852 3236 57856 3292
rect 57856 3236 57912 3292
rect 57912 3236 57916 3292
rect 57852 3232 57916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 21952 2748 22016 2752
rect 21952 2692 21956 2748
rect 21956 2692 22012 2748
rect 22012 2692 22016 2748
rect 21952 2688 22016 2692
rect 22032 2748 22096 2752
rect 22032 2692 22036 2748
rect 22036 2692 22092 2748
rect 22092 2692 22096 2748
rect 22032 2688 22096 2692
rect 22112 2748 22176 2752
rect 22112 2692 22116 2748
rect 22116 2692 22172 2748
rect 22172 2692 22176 2748
rect 22112 2688 22176 2692
rect 22192 2748 22256 2752
rect 22192 2692 22196 2748
rect 22196 2692 22252 2748
rect 22252 2692 22256 2748
rect 22192 2688 22256 2692
rect 26952 2748 27016 2752
rect 26952 2692 26956 2748
rect 26956 2692 27012 2748
rect 27012 2692 27016 2748
rect 26952 2688 27016 2692
rect 27032 2748 27096 2752
rect 27032 2692 27036 2748
rect 27036 2692 27092 2748
rect 27092 2692 27096 2748
rect 27032 2688 27096 2692
rect 27112 2748 27176 2752
rect 27112 2692 27116 2748
rect 27116 2692 27172 2748
rect 27172 2692 27176 2748
rect 27112 2688 27176 2692
rect 27192 2748 27256 2752
rect 27192 2692 27196 2748
rect 27196 2692 27252 2748
rect 27252 2692 27256 2748
rect 27192 2688 27256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 36952 2748 37016 2752
rect 36952 2692 36956 2748
rect 36956 2692 37012 2748
rect 37012 2692 37016 2748
rect 36952 2688 37016 2692
rect 37032 2748 37096 2752
rect 37032 2692 37036 2748
rect 37036 2692 37092 2748
rect 37092 2692 37096 2748
rect 37032 2688 37096 2692
rect 37112 2748 37176 2752
rect 37112 2692 37116 2748
rect 37116 2692 37172 2748
rect 37172 2692 37176 2748
rect 37112 2688 37176 2692
rect 37192 2748 37256 2752
rect 37192 2692 37196 2748
rect 37196 2692 37252 2748
rect 37252 2692 37256 2748
rect 37192 2688 37256 2692
rect 41952 2748 42016 2752
rect 41952 2692 41956 2748
rect 41956 2692 42012 2748
rect 42012 2692 42016 2748
rect 41952 2688 42016 2692
rect 42032 2748 42096 2752
rect 42032 2692 42036 2748
rect 42036 2692 42092 2748
rect 42092 2692 42096 2748
rect 42032 2688 42096 2692
rect 42112 2748 42176 2752
rect 42112 2692 42116 2748
rect 42116 2692 42172 2748
rect 42172 2692 42176 2748
rect 42112 2688 42176 2692
rect 42192 2748 42256 2752
rect 42192 2692 42196 2748
rect 42196 2692 42252 2748
rect 42252 2692 42256 2748
rect 42192 2688 42256 2692
rect 46952 2748 47016 2752
rect 46952 2692 46956 2748
rect 46956 2692 47012 2748
rect 47012 2692 47016 2748
rect 46952 2688 47016 2692
rect 47032 2748 47096 2752
rect 47032 2692 47036 2748
rect 47036 2692 47092 2748
rect 47092 2692 47096 2748
rect 47032 2688 47096 2692
rect 47112 2748 47176 2752
rect 47112 2692 47116 2748
rect 47116 2692 47172 2748
rect 47172 2692 47176 2748
rect 47112 2688 47176 2692
rect 47192 2748 47256 2752
rect 47192 2692 47196 2748
rect 47196 2692 47252 2748
rect 47252 2692 47256 2748
rect 47192 2688 47256 2692
rect 51952 2748 52016 2752
rect 51952 2692 51956 2748
rect 51956 2692 52012 2748
rect 52012 2692 52016 2748
rect 51952 2688 52016 2692
rect 52032 2748 52096 2752
rect 52032 2692 52036 2748
rect 52036 2692 52092 2748
rect 52092 2692 52096 2748
rect 52032 2688 52096 2692
rect 52112 2748 52176 2752
rect 52112 2692 52116 2748
rect 52116 2692 52172 2748
rect 52172 2692 52176 2748
rect 52112 2688 52176 2692
rect 52192 2748 52256 2752
rect 52192 2692 52196 2748
rect 52196 2692 52252 2748
rect 52252 2692 52256 2748
rect 52192 2688 52256 2692
rect 56952 2748 57016 2752
rect 56952 2692 56956 2748
rect 56956 2692 57012 2748
rect 57012 2692 57016 2748
rect 56952 2688 57016 2692
rect 57032 2748 57096 2752
rect 57032 2692 57036 2748
rect 57036 2692 57092 2748
rect 57092 2692 57096 2748
rect 57032 2688 57096 2692
rect 57112 2748 57176 2752
rect 57112 2692 57116 2748
rect 57116 2692 57172 2748
rect 57172 2692 57176 2748
rect 57112 2688 57176 2692
rect 57192 2748 57256 2752
rect 57192 2692 57196 2748
rect 57196 2692 57252 2748
rect 57252 2692 57256 2748
rect 57192 2688 57256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
rect 22612 2204 22676 2208
rect 22612 2148 22616 2204
rect 22616 2148 22672 2204
rect 22672 2148 22676 2204
rect 22612 2144 22676 2148
rect 22692 2204 22756 2208
rect 22692 2148 22696 2204
rect 22696 2148 22752 2204
rect 22752 2148 22756 2204
rect 22692 2144 22756 2148
rect 22772 2204 22836 2208
rect 22772 2148 22776 2204
rect 22776 2148 22832 2204
rect 22832 2148 22836 2204
rect 22772 2144 22836 2148
rect 22852 2204 22916 2208
rect 22852 2148 22856 2204
rect 22856 2148 22912 2204
rect 22912 2148 22916 2204
rect 22852 2144 22916 2148
rect 27612 2204 27676 2208
rect 27612 2148 27616 2204
rect 27616 2148 27672 2204
rect 27672 2148 27676 2204
rect 27612 2144 27676 2148
rect 27692 2204 27756 2208
rect 27692 2148 27696 2204
rect 27696 2148 27752 2204
rect 27752 2148 27756 2204
rect 27692 2144 27756 2148
rect 27772 2204 27836 2208
rect 27772 2148 27776 2204
rect 27776 2148 27832 2204
rect 27832 2148 27836 2204
rect 27772 2144 27836 2148
rect 27852 2204 27916 2208
rect 27852 2148 27856 2204
rect 27856 2148 27912 2204
rect 27912 2148 27916 2204
rect 27852 2144 27916 2148
rect 32612 2204 32676 2208
rect 32612 2148 32616 2204
rect 32616 2148 32672 2204
rect 32672 2148 32676 2204
rect 32612 2144 32676 2148
rect 32692 2204 32756 2208
rect 32692 2148 32696 2204
rect 32696 2148 32752 2204
rect 32752 2148 32756 2204
rect 32692 2144 32756 2148
rect 32772 2204 32836 2208
rect 32772 2148 32776 2204
rect 32776 2148 32832 2204
rect 32832 2148 32836 2204
rect 32772 2144 32836 2148
rect 32852 2204 32916 2208
rect 32852 2148 32856 2204
rect 32856 2148 32912 2204
rect 32912 2148 32916 2204
rect 32852 2144 32916 2148
rect 37612 2204 37676 2208
rect 37612 2148 37616 2204
rect 37616 2148 37672 2204
rect 37672 2148 37676 2204
rect 37612 2144 37676 2148
rect 37692 2204 37756 2208
rect 37692 2148 37696 2204
rect 37696 2148 37752 2204
rect 37752 2148 37756 2204
rect 37692 2144 37756 2148
rect 37772 2204 37836 2208
rect 37772 2148 37776 2204
rect 37776 2148 37832 2204
rect 37832 2148 37836 2204
rect 37772 2144 37836 2148
rect 37852 2204 37916 2208
rect 37852 2148 37856 2204
rect 37856 2148 37912 2204
rect 37912 2148 37916 2204
rect 37852 2144 37916 2148
rect 42612 2204 42676 2208
rect 42612 2148 42616 2204
rect 42616 2148 42672 2204
rect 42672 2148 42676 2204
rect 42612 2144 42676 2148
rect 42692 2204 42756 2208
rect 42692 2148 42696 2204
rect 42696 2148 42752 2204
rect 42752 2148 42756 2204
rect 42692 2144 42756 2148
rect 42772 2204 42836 2208
rect 42772 2148 42776 2204
rect 42776 2148 42832 2204
rect 42832 2148 42836 2204
rect 42772 2144 42836 2148
rect 42852 2204 42916 2208
rect 42852 2148 42856 2204
rect 42856 2148 42912 2204
rect 42912 2148 42916 2204
rect 42852 2144 42916 2148
rect 47612 2204 47676 2208
rect 47612 2148 47616 2204
rect 47616 2148 47672 2204
rect 47672 2148 47676 2204
rect 47612 2144 47676 2148
rect 47692 2204 47756 2208
rect 47692 2148 47696 2204
rect 47696 2148 47752 2204
rect 47752 2148 47756 2204
rect 47692 2144 47756 2148
rect 47772 2204 47836 2208
rect 47772 2148 47776 2204
rect 47776 2148 47832 2204
rect 47832 2148 47836 2204
rect 47772 2144 47836 2148
rect 47852 2204 47916 2208
rect 47852 2148 47856 2204
rect 47856 2148 47912 2204
rect 47912 2148 47916 2204
rect 47852 2144 47916 2148
rect 52612 2204 52676 2208
rect 52612 2148 52616 2204
rect 52616 2148 52672 2204
rect 52672 2148 52676 2204
rect 52612 2144 52676 2148
rect 52692 2204 52756 2208
rect 52692 2148 52696 2204
rect 52696 2148 52752 2204
rect 52752 2148 52756 2204
rect 52692 2144 52756 2148
rect 52772 2204 52836 2208
rect 52772 2148 52776 2204
rect 52776 2148 52832 2204
rect 52832 2148 52836 2204
rect 52772 2144 52836 2148
rect 52852 2204 52916 2208
rect 52852 2148 52856 2204
rect 52856 2148 52912 2204
rect 52912 2148 52916 2204
rect 52852 2144 52916 2148
rect 57612 2204 57676 2208
rect 57612 2148 57616 2204
rect 57616 2148 57672 2204
rect 57672 2148 57676 2204
rect 57612 2144 57676 2148
rect 57692 2204 57756 2208
rect 57692 2148 57696 2204
rect 57696 2148 57752 2204
rect 57752 2148 57756 2204
rect 57692 2144 57756 2148
rect 57772 2204 57836 2208
rect 57772 2148 57776 2204
rect 57776 2148 57832 2204
rect 57832 2148 57836 2204
rect 57772 2144 57836 2148
rect 57852 2204 57916 2208
rect 57852 2148 57856 2204
rect 57856 2148 57912 2204
rect 57912 2148 57916 2204
rect 57852 2144 57916 2148
<< metal4 >>
rect 1944 57152 2264 57712
rect 1944 57088 1952 57152
rect 2016 57088 2032 57152
rect 2096 57088 2112 57152
rect 2176 57088 2192 57152
rect 2256 57088 2264 57152
rect 1944 56064 2264 57088
rect 1944 56000 1952 56064
rect 2016 56000 2032 56064
rect 2096 56000 2112 56064
rect 2176 56000 2192 56064
rect 2256 56000 2264 56064
rect 1944 54976 2264 56000
rect 1944 54912 1952 54976
rect 2016 54912 2032 54976
rect 2096 54912 2112 54976
rect 2176 54912 2192 54976
rect 2256 54912 2264 54976
rect 1944 53888 2264 54912
rect 1944 53824 1952 53888
rect 2016 53824 2032 53888
rect 2096 53824 2112 53888
rect 2176 53824 2192 53888
rect 2256 53824 2264 53888
rect 1944 53294 2264 53824
rect 1944 53058 1986 53294
rect 2222 53058 2264 53294
rect 1944 52800 2264 53058
rect 1944 52736 1952 52800
rect 2016 52736 2032 52800
rect 2096 52736 2112 52800
rect 2176 52736 2192 52800
rect 2256 52736 2264 52800
rect 1944 51712 2264 52736
rect 1944 51648 1952 51712
rect 2016 51648 2032 51712
rect 2096 51648 2112 51712
rect 2176 51648 2192 51712
rect 2256 51648 2264 51712
rect 1944 50624 2264 51648
rect 1944 50560 1952 50624
rect 2016 50560 2032 50624
rect 2096 50560 2112 50624
rect 2176 50560 2192 50624
rect 2256 50560 2264 50624
rect 1944 49536 2264 50560
rect 1944 49472 1952 49536
rect 2016 49472 2032 49536
rect 2096 49472 2112 49536
rect 2176 49472 2192 49536
rect 2256 49472 2264 49536
rect 1944 48448 2264 49472
rect 1944 48384 1952 48448
rect 2016 48384 2032 48448
rect 2096 48384 2112 48448
rect 2176 48384 2192 48448
rect 2256 48384 2264 48448
rect 1944 48294 2264 48384
rect 1944 48058 1986 48294
rect 2222 48058 2264 48294
rect 1944 47360 2264 48058
rect 1944 47296 1952 47360
rect 2016 47296 2032 47360
rect 2096 47296 2112 47360
rect 2176 47296 2192 47360
rect 2256 47296 2264 47360
rect 1944 46272 2264 47296
rect 1944 46208 1952 46272
rect 2016 46208 2032 46272
rect 2096 46208 2112 46272
rect 2176 46208 2192 46272
rect 2256 46208 2264 46272
rect 1944 45184 2264 46208
rect 1944 45120 1952 45184
rect 2016 45120 2032 45184
rect 2096 45120 2112 45184
rect 2176 45120 2192 45184
rect 2256 45120 2264 45184
rect 1944 44096 2264 45120
rect 1944 44032 1952 44096
rect 2016 44032 2032 44096
rect 2096 44032 2112 44096
rect 2176 44032 2192 44096
rect 2256 44032 2264 44096
rect 1944 43294 2264 44032
rect 1944 43058 1986 43294
rect 2222 43058 2264 43294
rect 1944 43008 2264 43058
rect 1944 42944 1952 43008
rect 2016 42944 2032 43008
rect 2096 42944 2112 43008
rect 2176 42944 2192 43008
rect 2256 42944 2264 43008
rect 1944 41920 2264 42944
rect 1944 41856 1952 41920
rect 2016 41856 2032 41920
rect 2096 41856 2112 41920
rect 2176 41856 2192 41920
rect 2256 41856 2264 41920
rect 1944 40832 2264 41856
rect 1944 40768 1952 40832
rect 2016 40768 2032 40832
rect 2096 40768 2112 40832
rect 2176 40768 2192 40832
rect 2256 40768 2264 40832
rect 1944 39744 2264 40768
rect 1944 39680 1952 39744
rect 2016 39680 2032 39744
rect 2096 39680 2112 39744
rect 2176 39680 2192 39744
rect 2256 39680 2264 39744
rect 1944 38656 2264 39680
rect 1944 38592 1952 38656
rect 2016 38592 2032 38656
rect 2096 38592 2112 38656
rect 2176 38592 2192 38656
rect 2256 38592 2264 38656
rect 1944 38294 2264 38592
rect 1944 38058 1986 38294
rect 2222 38058 2264 38294
rect 1944 37568 2264 38058
rect 1944 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2264 37568
rect 1944 36480 2264 37504
rect 1944 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2264 36480
rect 1944 35392 2264 36416
rect 1944 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2264 35392
rect 1944 34304 2264 35328
rect 1944 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2264 34304
rect 1944 33294 2264 34240
rect 1944 33216 1986 33294
rect 2222 33216 2264 33294
rect 1944 33152 1952 33216
rect 2256 33152 2264 33216
rect 1944 33058 1986 33152
rect 2222 33058 2264 33152
rect 1944 32128 2264 33058
rect 1944 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2264 32128
rect 1944 31040 2264 32064
rect 1944 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2264 31040
rect 1944 29952 2264 30976
rect 1944 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2264 29952
rect 1944 28864 2264 29888
rect 1944 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2264 28864
rect 1944 28294 2264 28800
rect 1944 28058 1986 28294
rect 2222 28058 2264 28294
rect 1944 27776 2264 28058
rect 1944 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2264 27776
rect 1944 26688 2264 27712
rect 1944 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2264 26688
rect 1944 25600 2264 26624
rect 1944 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2264 25600
rect 1944 24512 2264 25536
rect 1944 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2264 24512
rect 1944 23424 2264 24448
rect 1944 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2264 23424
rect 1944 23294 2264 23360
rect 1944 23058 1986 23294
rect 2222 23058 2264 23294
rect 1944 22336 2264 23058
rect 1944 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2264 22336
rect 1944 21248 2264 22272
rect 1944 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2264 21248
rect 1944 20160 2264 21184
rect 1944 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2264 20160
rect 1944 19072 2264 20096
rect 1944 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2264 19072
rect 1944 18294 2264 19008
rect 1944 18058 1986 18294
rect 2222 18058 2264 18294
rect 1944 17984 2264 18058
rect 1944 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2264 17984
rect 1944 16896 2264 17920
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 57696 2924 57712
rect 2604 57632 2612 57696
rect 2676 57632 2692 57696
rect 2756 57632 2772 57696
rect 2836 57632 2852 57696
rect 2916 57632 2924 57696
rect 2604 56608 2924 57632
rect 2604 56544 2612 56608
rect 2676 56544 2692 56608
rect 2756 56544 2772 56608
rect 2836 56544 2852 56608
rect 2916 56544 2924 56608
rect 2604 55520 2924 56544
rect 2604 55456 2612 55520
rect 2676 55456 2692 55520
rect 2756 55456 2772 55520
rect 2836 55456 2852 55520
rect 2916 55456 2924 55520
rect 2604 54432 2924 55456
rect 2604 54368 2612 54432
rect 2676 54368 2692 54432
rect 2756 54368 2772 54432
rect 2836 54368 2852 54432
rect 2916 54368 2924 54432
rect 2604 53954 2924 54368
rect 2604 53718 2646 53954
rect 2882 53718 2924 53954
rect 2604 53344 2924 53718
rect 2604 53280 2612 53344
rect 2676 53280 2692 53344
rect 2756 53280 2772 53344
rect 2836 53280 2852 53344
rect 2916 53280 2924 53344
rect 2604 52256 2924 53280
rect 2604 52192 2612 52256
rect 2676 52192 2692 52256
rect 2756 52192 2772 52256
rect 2836 52192 2852 52256
rect 2916 52192 2924 52256
rect 2604 51168 2924 52192
rect 2604 51104 2612 51168
rect 2676 51104 2692 51168
rect 2756 51104 2772 51168
rect 2836 51104 2852 51168
rect 2916 51104 2924 51168
rect 2604 50080 2924 51104
rect 2604 50016 2612 50080
rect 2676 50016 2692 50080
rect 2756 50016 2772 50080
rect 2836 50016 2852 50080
rect 2916 50016 2924 50080
rect 2604 48992 2924 50016
rect 2604 48928 2612 48992
rect 2676 48954 2692 48992
rect 2756 48954 2772 48992
rect 2836 48954 2852 48992
rect 2916 48928 2924 48992
rect 2604 48718 2646 48928
rect 2882 48718 2924 48928
rect 2604 47904 2924 48718
rect 2604 47840 2612 47904
rect 2676 47840 2692 47904
rect 2756 47840 2772 47904
rect 2836 47840 2852 47904
rect 2916 47840 2924 47904
rect 2604 46816 2924 47840
rect 2604 46752 2612 46816
rect 2676 46752 2692 46816
rect 2756 46752 2772 46816
rect 2836 46752 2852 46816
rect 2916 46752 2924 46816
rect 2604 45728 2924 46752
rect 2604 45664 2612 45728
rect 2676 45664 2692 45728
rect 2756 45664 2772 45728
rect 2836 45664 2852 45728
rect 2916 45664 2924 45728
rect 2604 44640 2924 45664
rect 2604 44576 2612 44640
rect 2676 44576 2692 44640
rect 2756 44576 2772 44640
rect 2836 44576 2852 44640
rect 2916 44576 2924 44640
rect 2604 43954 2924 44576
rect 2604 43718 2646 43954
rect 2882 43718 2924 43954
rect 2604 43552 2924 43718
rect 2604 43488 2612 43552
rect 2676 43488 2692 43552
rect 2756 43488 2772 43552
rect 2836 43488 2852 43552
rect 2916 43488 2924 43552
rect 2604 42464 2924 43488
rect 2604 42400 2612 42464
rect 2676 42400 2692 42464
rect 2756 42400 2772 42464
rect 2836 42400 2852 42464
rect 2916 42400 2924 42464
rect 2604 41376 2924 42400
rect 2604 41312 2612 41376
rect 2676 41312 2692 41376
rect 2756 41312 2772 41376
rect 2836 41312 2852 41376
rect 2916 41312 2924 41376
rect 2604 40288 2924 41312
rect 2604 40224 2612 40288
rect 2676 40224 2692 40288
rect 2756 40224 2772 40288
rect 2836 40224 2852 40288
rect 2916 40224 2924 40288
rect 2604 39200 2924 40224
rect 2604 39136 2612 39200
rect 2676 39136 2692 39200
rect 2756 39136 2772 39200
rect 2836 39136 2852 39200
rect 2916 39136 2924 39200
rect 2604 38954 2924 39136
rect 2604 38718 2646 38954
rect 2882 38718 2924 38954
rect 2604 38112 2924 38718
rect 2604 38048 2612 38112
rect 2676 38048 2692 38112
rect 2756 38048 2772 38112
rect 2836 38048 2852 38112
rect 2916 38048 2924 38112
rect 2604 37024 2924 38048
rect 2604 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2924 37024
rect 2604 35936 2924 36960
rect 2604 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2924 35936
rect 2604 34848 2924 35872
rect 2604 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2924 34848
rect 2604 33954 2924 34784
rect 2604 33760 2646 33954
rect 2882 33760 2924 33954
rect 2604 33696 2612 33760
rect 2676 33696 2692 33718
rect 2756 33696 2772 33718
rect 2836 33696 2852 33718
rect 2916 33696 2924 33760
rect 2604 32672 2924 33696
rect 2604 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2924 32672
rect 2604 31584 2924 32608
rect 2604 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2924 31584
rect 2604 30496 2924 31520
rect 2604 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2924 30496
rect 2604 29408 2924 30432
rect 2604 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2924 29408
rect 2604 28954 2924 29344
rect 2604 28718 2646 28954
rect 2882 28718 2924 28954
rect 2604 28320 2924 28718
rect 2604 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2924 28320
rect 2604 27232 2924 28256
rect 2604 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2924 27232
rect 2604 26144 2924 27168
rect 2604 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2924 26144
rect 2604 25056 2924 26080
rect 2604 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2924 25056
rect 2604 23968 2924 24992
rect 2604 23904 2612 23968
rect 2676 23954 2692 23968
rect 2756 23954 2772 23968
rect 2836 23954 2852 23968
rect 2916 23904 2924 23968
rect 2604 23718 2646 23904
rect 2882 23718 2924 23904
rect 2604 22880 2924 23718
rect 2604 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2924 22880
rect 2604 21792 2924 22816
rect 2604 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2924 21792
rect 2604 20704 2924 21728
rect 2604 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2924 20704
rect 2604 19616 2924 20640
rect 2604 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2924 19616
rect 2604 18954 2924 19552
rect 2604 18718 2646 18954
rect 2882 18718 2924 18954
rect 2604 18528 2924 18718
rect 2604 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2924 18528
rect 2604 17440 2924 18464
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 2604 13088 2924 13718
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 57152 7264 57712
rect 6944 57088 6952 57152
rect 7016 57088 7032 57152
rect 7096 57088 7112 57152
rect 7176 57088 7192 57152
rect 7256 57088 7264 57152
rect 6944 56064 7264 57088
rect 6944 56000 6952 56064
rect 7016 56000 7032 56064
rect 7096 56000 7112 56064
rect 7176 56000 7192 56064
rect 7256 56000 7264 56064
rect 6944 54976 7264 56000
rect 6944 54912 6952 54976
rect 7016 54912 7032 54976
rect 7096 54912 7112 54976
rect 7176 54912 7192 54976
rect 7256 54912 7264 54976
rect 6944 53888 7264 54912
rect 6944 53824 6952 53888
rect 7016 53824 7032 53888
rect 7096 53824 7112 53888
rect 7176 53824 7192 53888
rect 7256 53824 7264 53888
rect 6944 53294 7264 53824
rect 6944 53058 6986 53294
rect 7222 53058 7264 53294
rect 6944 52800 7264 53058
rect 6944 52736 6952 52800
rect 7016 52736 7032 52800
rect 7096 52736 7112 52800
rect 7176 52736 7192 52800
rect 7256 52736 7264 52800
rect 6944 51712 7264 52736
rect 6944 51648 6952 51712
rect 7016 51648 7032 51712
rect 7096 51648 7112 51712
rect 7176 51648 7192 51712
rect 7256 51648 7264 51712
rect 6944 50624 7264 51648
rect 6944 50560 6952 50624
rect 7016 50560 7032 50624
rect 7096 50560 7112 50624
rect 7176 50560 7192 50624
rect 7256 50560 7264 50624
rect 6944 49536 7264 50560
rect 6944 49472 6952 49536
rect 7016 49472 7032 49536
rect 7096 49472 7112 49536
rect 7176 49472 7192 49536
rect 7256 49472 7264 49536
rect 6944 48448 7264 49472
rect 6944 48384 6952 48448
rect 7016 48384 7032 48448
rect 7096 48384 7112 48448
rect 7176 48384 7192 48448
rect 7256 48384 7264 48448
rect 6944 48294 7264 48384
rect 6944 48058 6986 48294
rect 7222 48058 7264 48294
rect 6944 47360 7264 48058
rect 6944 47296 6952 47360
rect 7016 47296 7032 47360
rect 7096 47296 7112 47360
rect 7176 47296 7192 47360
rect 7256 47296 7264 47360
rect 6944 46272 7264 47296
rect 6944 46208 6952 46272
rect 7016 46208 7032 46272
rect 7096 46208 7112 46272
rect 7176 46208 7192 46272
rect 7256 46208 7264 46272
rect 6944 45184 7264 46208
rect 6944 45120 6952 45184
rect 7016 45120 7032 45184
rect 7096 45120 7112 45184
rect 7176 45120 7192 45184
rect 7256 45120 7264 45184
rect 6944 44096 7264 45120
rect 6944 44032 6952 44096
rect 7016 44032 7032 44096
rect 7096 44032 7112 44096
rect 7176 44032 7192 44096
rect 7256 44032 7264 44096
rect 6944 43294 7264 44032
rect 6944 43058 6986 43294
rect 7222 43058 7264 43294
rect 6944 43008 7264 43058
rect 6944 42944 6952 43008
rect 7016 42944 7032 43008
rect 7096 42944 7112 43008
rect 7176 42944 7192 43008
rect 7256 42944 7264 43008
rect 6944 41920 7264 42944
rect 6944 41856 6952 41920
rect 7016 41856 7032 41920
rect 7096 41856 7112 41920
rect 7176 41856 7192 41920
rect 7256 41856 7264 41920
rect 6944 40832 7264 41856
rect 6944 40768 6952 40832
rect 7016 40768 7032 40832
rect 7096 40768 7112 40832
rect 7176 40768 7192 40832
rect 7256 40768 7264 40832
rect 6944 39744 7264 40768
rect 6944 39680 6952 39744
rect 7016 39680 7032 39744
rect 7096 39680 7112 39744
rect 7176 39680 7192 39744
rect 7256 39680 7264 39744
rect 6944 38656 7264 39680
rect 6944 38592 6952 38656
rect 7016 38592 7032 38656
rect 7096 38592 7112 38656
rect 7176 38592 7192 38656
rect 7256 38592 7264 38656
rect 6944 38294 7264 38592
rect 6944 38058 6986 38294
rect 7222 38058 7264 38294
rect 6944 37568 7264 38058
rect 6944 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7264 37568
rect 6944 36480 7264 37504
rect 6944 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7264 36480
rect 6944 35392 7264 36416
rect 6944 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7264 35392
rect 6944 34304 7264 35328
rect 6944 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7264 34304
rect 6944 33294 7264 34240
rect 6944 33216 6986 33294
rect 7222 33216 7264 33294
rect 6944 33152 6952 33216
rect 7256 33152 7264 33216
rect 6944 33058 6986 33152
rect 7222 33058 7264 33152
rect 6944 32128 7264 33058
rect 6944 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7264 32128
rect 6944 31040 7264 32064
rect 6944 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7264 31040
rect 6944 29952 7264 30976
rect 6944 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7264 29952
rect 6944 28864 7264 29888
rect 6944 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7264 28864
rect 6944 28294 7264 28800
rect 6944 28058 6986 28294
rect 7222 28058 7264 28294
rect 6944 27776 7264 28058
rect 6944 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7264 27776
rect 6944 26688 7264 27712
rect 6944 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7264 26688
rect 6944 25600 7264 26624
rect 6944 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7264 25600
rect 6944 24512 7264 25536
rect 6944 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7264 24512
rect 6944 23424 7264 24448
rect 6944 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7264 23424
rect 6944 23294 7264 23360
rect 6944 23058 6986 23294
rect 7222 23058 7264 23294
rect 6944 22336 7264 23058
rect 6944 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7264 22336
rect 6944 21248 7264 22272
rect 6944 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7264 21248
rect 6944 20160 7264 21184
rect 6944 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7264 20160
rect 6944 19072 7264 20096
rect 6944 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7264 19072
rect 6944 18294 7264 19008
rect 6944 18058 6986 18294
rect 7222 18058 7264 18294
rect 6944 17984 7264 18058
rect 6944 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7264 17984
rect 6944 16896 7264 17920
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 57696 7924 57712
rect 7604 57632 7612 57696
rect 7676 57632 7692 57696
rect 7756 57632 7772 57696
rect 7836 57632 7852 57696
rect 7916 57632 7924 57696
rect 7604 56608 7924 57632
rect 7604 56544 7612 56608
rect 7676 56544 7692 56608
rect 7756 56544 7772 56608
rect 7836 56544 7852 56608
rect 7916 56544 7924 56608
rect 7604 55520 7924 56544
rect 7604 55456 7612 55520
rect 7676 55456 7692 55520
rect 7756 55456 7772 55520
rect 7836 55456 7852 55520
rect 7916 55456 7924 55520
rect 7604 54432 7924 55456
rect 7604 54368 7612 54432
rect 7676 54368 7692 54432
rect 7756 54368 7772 54432
rect 7836 54368 7852 54432
rect 7916 54368 7924 54432
rect 7604 53954 7924 54368
rect 7604 53718 7646 53954
rect 7882 53718 7924 53954
rect 7604 53344 7924 53718
rect 7604 53280 7612 53344
rect 7676 53280 7692 53344
rect 7756 53280 7772 53344
rect 7836 53280 7852 53344
rect 7916 53280 7924 53344
rect 7604 52256 7924 53280
rect 7604 52192 7612 52256
rect 7676 52192 7692 52256
rect 7756 52192 7772 52256
rect 7836 52192 7852 52256
rect 7916 52192 7924 52256
rect 7604 51168 7924 52192
rect 7604 51104 7612 51168
rect 7676 51104 7692 51168
rect 7756 51104 7772 51168
rect 7836 51104 7852 51168
rect 7916 51104 7924 51168
rect 7604 50080 7924 51104
rect 7604 50016 7612 50080
rect 7676 50016 7692 50080
rect 7756 50016 7772 50080
rect 7836 50016 7852 50080
rect 7916 50016 7924 50080
rect 7604 48992 7924 50016
rect 7604 48928 7612 48992
rect 7676 48954 7692 48992
rect 7756 48954 7772 48992
rect 7836 48954 7852 48992
rect 7916 48928 7924 48992
rect 7604 48718 7646 48928
rect 7882 48718 7924 48928
rect 7604 47904 7924 48718
rect 7604 47840 7612 47904
rect 7676 47840 7692 47904
rect 7756 47840 7772 47904
rect 7836 47840 7852 47904
rect 7916 47840 7924 47904
rect 7604 46816 7924 47840
rect 7604 46752 7612 46816
rect 7676 46752 7692 46816
rect 7756 46752 7772 46816
rect 7836 46752 7852 46816
rect 7916 46752 7924 46816
rect 7604 45728 7924 46752
rect 7604 45664 7612 45728
rect 7676 45664 7692 45728
rect 7756 45664 7772 45728
rect 7836 45664 7852 45728
rect 7916 45664 7924 45728
rect 7604 44640 7924 45664
rect 7604 44576 7612 44640
rect 7676 44576 7692 44640
rect 7756 44576 7772 44640
rect 7836 44576 7852 44640
rect 7916 44576 7924 44640
rect 7604 43954 7924 44576
rect 7604 43718 7646 43954
rect 7882 43718 7924 43954
rect 7604 43552 7924 43718
rect 7604 43488 7612 43552
rect 7676 43488 7692 43552
rect 7756 43488 7772 43552
rect 7836 43488 7852 43552
rect 7916 43488 7924 43552
rect 7604 42464 7924 43488
rect 7604 42400 7612 42464
rect 7676 42400 7692 42464
rect 7756 42400 7772 42464
rect 7836 42400 7852 42464
rect 7916 42400 7924 42464
rect 7604 41376 7924 42400
rect 7604 41312 7612 41376
rect 7676 41312 7692 41376
rect 7756 41312 7772 41376
rect 7836 41312 7852 41376
rect 7916 41312 7924 41376
rect 7604 40288 7924 41312
rect 7604 40224 7612 40288
rect 7676 40224 7692 40288
rect 7756 40224 7772 40288
rect 7836 40224 7852 40288
rect 7916 40224 7924 40288
rect 7604 39200 7924 40224
rect 7604 39136 7612 39200
rect 7676 39136 7692 39200
rect 7756 39136 7772 39200
rect 7836 39136 7852 39200
rect 7916 39136 7924 39200
rect 7604 38954 7924 39136
rect 7604 38718 7646 38954
rect 7882 38718 7924 38954
rect 7604 38112 7924 38718
rect 7604 38048 7612 38112
rect 7676 38048 7692 38112
rect 7756 38048 7772 38112
rect 7836 38048 7852 38112
rect 7916 38048 7924 38112
rect 7604 37024 7924 38048
rect 7604 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7924 37024
rect 7604 35936 7924 36960
rect 7604 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7924 35936
rect 7604 34848 7924 35872
rect 7604 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7924 34848
rect 7604 33954 7924 34784
rect 7604 33760 7646 33954
rect 7882 33760 7924 33954
rect 7604 33696 7612 33760
rect 7676 33696 7692 33718
rect 7756 33696 7772 33718
rect 7836 33696 7852 33718
rect 7916 33696 7924 33760
rect 7604 32672 7924 33696
rect 7604 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7924 32672
rect 7604 31584 7924 32608
rect 7604 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7924 31584
rect 7604 30496 7924 31520
rect 7604 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7924 30496
rect 7604 29408 7924 30432
rect 7604 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7924 29408
rect 7604 28954 7924 29344
rect 7604 28718 7646 28954
rect 7882 28718 7924 28954
rect 7604 28320 7924 28718
rect 7604 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7924 28320
rect 7604 27232 7924 28256
rect 7604 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7924 27232
rect 7604 26144 7924 27168
rect 7604 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7924 26144
rect 7604 25056 7924 26080
rect 7604 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7924 25056
rect 7604 23968 7924 24992
rect 7604 23904 7612 23968
rect 7676 23954 7692 23968
rect 7756 23954 7772 23968
rect 7836 23954 7852 23968
rect 7916 23904 7924 23968
rect 7604 23718 7646 23904
rect 7882 23718 7924 23904
rect 7604 22880 7924 23718
rect 7604 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7924 22880
rect 7604 21792 7924 22816
rect 7604 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7924 21792
rect 7604 20704 7924 21728
rect 7604 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7924 20704
rect 7604 19616 7924 20640
rect 7604 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7924 19616
rect 7604 18954 7924 19552
rect 7604 18718 7646 18954
rect 7882 18718 7924 18954
rect 7604 18528 7924 18718
rect 7604 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7924 18528
rect 7604 17440 7924 18464
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7604 7648 7924 8672
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11944 57152 12264 57712
rect 11944 57088 11952 57152
rect 12016 57088 12032 57152
rect 12096 57088 12112 57152
rect 12176 57088 12192 57152
rect 12256 57088 12264 57152
rect 11944 56064 12264 57088
rect 11944 56000 11952 56064
rect 12016 56000 12032 56064
rect 12096 56000 12112 56064
rect 12176 56000 12192 56064
rect 12256 56000 12264 56064
rect 11944 54976 12264 56000
rect 11944 54912 11952 54976
rect 12016 54912 12032 54976
rect 12096 54912 12112 54976
rect 12176 54912 12192 54976
rect 12256 54912 12264 54976
rect 11944 53888 12264 54912
rect 11944 53824 11952 53888
rect 12016 53824 12032 53888
rect 12096 53824 12112 53888
rect 12176 53824 12192 53888
rect 12256 53824 12264 53888
rect 11944 53294 12264 53824
rect 11944 53058 11986 53294
rect 12222 53058 12264 53294
rect 11944 52800 12264 53058
rect 11944 52736 11952 52800
rect 12016 52736 12032 52800
rect 12096 52736 12112 52800
rect 12176 52736 12192 52800
rect 12256 52736 12264 52800
rect 11944 51712 12264 52736
rect 11944 51648 11952 51712
rect 12016 51648 12032 51712
rect 12096 51648 12112 51712
rect 12176 51648 12192 51712
rect 12256 51648 12264 51712
rect 11944 50624 12264 51648
rect 11944 50560 11952 50624
rect 12016 50560 12032 50624
rect 12096 50560 12112 50624
rect 12176 50560 12192 50624
rect 12256 50560 12264 50624
rect 11944 49536 12264 50560
rect 11944 49472 11952 49536
rect 12016 49472 12032 49536
rect 12096 49472 12112 49536
rect 12176 49472 12192 49536
rect 12256 49472 12264 49536
rect 11944 48448 12264 49472
rect 11944 48384 11952 48448
rect 12016 48384 12032 48448
rect 12096 48384 12112 48448
rect 12176 48384 12192 48448
rect 12256 48384 12264 48448
rect 11944 48294 12264 48384
rect 11944 48058 11986 48294
rect 12222 48058 12264 48294
rect 11944 47360 12264 48058
rect 11944 47296 11952 47360
rect 12016 47296 12032 47360
rect 12096 47296 12112 47360
rect 12176 47296 12192 47360
rect 12256 47296 12264 47360
rect 11944 46272 12264 47296
rect 11944 46208 11952 46272
rect 12016 46208 12032 46272
rect 12096 46208 12112 46272
rect 12176 46208 12192 46272
rect 12256 46208 12264 46272
rect 11944 45184 12264 46208
rect 11944 45120 11952 45184
rect 12016 45120 12032 45184
rect 12096 45120 12112 45184
rect 12176 45120 12192 45184
rect 12256 45120 12264 45184
rect 11944 44096 12264 45120
rect 11944 44032 11952 44096
rect 12016 44032 12032 44096
rect 12096 44032 12112 44096
rect 12176 44032 12192 44096
rect 12256 44032 12264 44096
rect 11944 43294 12264 44032
rect 11944 43058 11986 43294
rect 12222 43058 12264 43294
rect 11944 43008 12264 43058
rect 11944 42944 11952 43008
rect 12016 42944 12032 43008
rect 12096 42944 12112 43008
rect 12176 42944 12192 43008
rect 12256 42944 12264 43008
rect 11944 41920 12264 42944
rect 11944 41856 11952 41920
rect 12016 41856 12032 41920
rect 12096 41856 12112 41920
rect 12176 41856 12192 41920
rect 12256 41856 12264 41920
rect 11944 40832 12264 41856
rect 11944 40768 11952 40832
rect 12016 40768 12032 40832
rect 12096 40768 12112 40832
rect 12176 40768 12192 40832
rect 12256 40768 12264 40832
rect 11944 39744 12264 40768
rect 11944 39680 11952 39744
rect 12016 39680 12032 39744
rect 12096 39680 12112 39744
rect 12176 39680 12192 39744
rect 12256 39680 12264 39744
rect 11944 38656 12264 39680
rect 11944 38592 11952 38656
rect 12016 38592 12032 38656
rect 12096 38592 12112 38656
rect 12176 38592 12192 38656
rect 12256 38592 12264 38656
rect 11944 38294 12264 38592
rect 11944 38058 11986 38294
rect 12222 38058 12264 38294
rect 11944 37568 12264 38058
rect 11944 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12264 37568
rect 11944 36480 12264 37504
rect 11944 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12264 36480
rect 11944 35392 12264 36416
rect 11944 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12264 35392
rect 11944 34304 12264 35328
rect 11944 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12264 34304
rect 11944 33294 12264 34240
rect 11944 33216 11986 33294
rect 12222 33216 12264 33294
rect 11944 33152 11952 33216
rect 12256 33152 12264 33216
rect 11944 33058 11986 33152
rect 12222 33058 12264 33152
rect 11944 32128 12264 33058
rect 11944 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12264 32128
rect 11944 31040 12264 32064
rect 11944 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12264 31040
rect 11944 29952 12264 30976
rect 11944 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12264 29952
rect 11944 28864 12264 29888
rect 11944 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12264 28864
rect 11944 28294 12264 28800
rect 11944 28058 11986 28294
rect 12222 28058 12264 28294
rect 11944 27776 12264 28058
rect 11944 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12264 27776
rect 11944 26688 12264 27712
rect 11944 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12264 26688
rect 11944 25600 12264 26624
rect 11944 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12264 25600
rect 11944 24512 12264 25536
rect 11944 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12264 24512
rect 11944 23424 12264 24448
rect 11944 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12264 23424
rect 11944 23294 12264 23360
rect 11944 23058 11986 23294
rect 12222 23058 12264 23294
rect 11944 22336 12264 23058
rect 11944 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12264 22336
rect 11944 21248 12264 22272
rect 11944 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12264 21248
rect 11944 20160 12264 21184
rect 11944 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12264 20160
rect 11944 19072 12264 20096
rect 11944 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12264 19072
rect 11944 18294 12264 19008
rect 11944 18058 11986 18294
rect 12222 18058 12264 18294
rect 11944 17984 12264 18058
rect 11944 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12264 17984
rect 11944 16896 12264 17920
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11944 13632 12264 14656
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11944 11456 12264 12480
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11944 4928 12264 5952
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11944 3294 12264 3776
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 11944 2128 12264 2688
rect 12604 57696 12924 57712
rect 12604 57632 12612 57696
rect 12676 57632 12692 57696
rect 12756 57632 12772 57696
rect 12836 57632 12852 57696
rect 12916 57632 12924 57696
rect 12604 56608 12924 57632
rect 12604 56544 12612 56608
rect 12676 56544 12692 56608
rect 12756 56544 12772 56608
rect 12836 56544 12852 56608
rect 12916 56544 12924 56608
rect 12604 55520 12924 56544
rect 12604 55456 12612 55520
rect 12676 55456 12692 55520
rect 12756 55456 12772 55520
rect 12836 55456 12852 55520
rect 12916 55456 12924 55520
rect 12604 54432 12924 55456
rect 12604 54368 12612 54432
rect 12676 54368 12692 54432
rect 12756 54368 12772 54432
rect 12836 54368 12852 54432
rect 12916 54368 12924 54432
rect 12604 53954 12924 54368
rect 12604 53718 12646 53954
rect 12882 53718 12924 53954
rect 12604 53344 12924 53718
rect 12604 53280 12612 53344
rect 12676 53280 12692 53344
rect 12756 53280 12772 53344
rect 12836 53280 12852 53344
rect 12916 53280 12924 53344
rect 12604 52256 12924 53280
rect 12604 52192 12612 52256
rect 12676 52192 12692 52256
rect 12756 52192 12772 52256
rect 12836 52192 12852 52256
rect 12916 52192 12924 52256
rect 12604 51168 12924 52192
rect 12604 51104 12612 51168
rect 12676 51104 12692 51168
rect 12756 51104 12772 51168
rect 12836 51104 12852 51168
rect 12916 51104 12924 51168
rect 12604 50080 12924 51104
rect 12604 50016 12612 50080
rect 12676 50016 12692 50080
rect 12756 50016 12772 50080
rect 12836 50016 12852 50080
rect 12916 50016 12924 50080
rect 12604 48992 12924 50016
rect 12604 48928 12612 48992
rect 12676 48954 12692 48992
rect 12756 48954 12772 48992
rect 12836 48954 12852 48992
rect 12916 48928 12924 48992
rect 12604 48718 12646 48928
rect 12882 48718 12924 48928
rect 12604 47904 12924 48718
rect 12604 47840 12612 47904
rect 12676 47840 12692 47904
rect 12756 47840 12772 47904
rect 12836 47840 12852 47904
rect 12916 47840 12924 47904
rect 12604 46816 12924 47840
rect 12604 46752 12612 46816
rect 12676 46752 12692 46816
rect 12756 46752 12772 46816
rect 12836 46752 12852 46816
rect 12916 46752 12924 46816
rect 12604 45728 12924 46752
rect 12604 45664 12612 45728
rect 12676 45664 12692 45728
rect 12756 45664 12772 45728
rect 12836 45664 12852 45728
rect 12916 45664 12924 45728
rect 12604 44640 12924 45664
rect 12604 44576 12612 44640
rect 12676 44576 12692 44640
rect 12756 44576 12772 44640
rect 12836 44576 12852 44640
rect 12916 44576 12924 44640
rect 12604 43954 12924 44576
rect 12604 43718 12646 43954
rect 12882 43718 12924 43954
rect 12604 43552 12924 43718
rect 12604 43488 12612 43552
rect 12676 43488 12692 43552
rect 12756 43488 12772 43552
rect 12836 43488 12852 43552
rect 12916 43488 12924 43552
rect 12604 42464 12924 43488
rect 12604 42400 12612 42464
rect 12676 42400 12692 42464
rect 12756 42400 12772 42464
rect 12836 42400 12852 42464
rect 12916 42400 12924 42464
rect 12604 41376 12924 42400
rect 12604 41312 12612 41376
rect 12676 41312 12692 41376
rect 12756 41312 12772 41376
rect 12836 41312 12852 41376
rect 12916 41312 12924 41376
rect 12604 40288 12924 41312
rect 12604 40224 12612 40288
rect 12676 40224 12692 40288
rect 12756 40224 12772 40288
rect 12836 40224 12852 40288
rect 12916 40224 12924 40288
rect 12604 39200 12924 40224
rect 12604 39136 12612 39200
rect 12676 39136 12692 39200
rect 12756 39136 12772 39200
rect 12836 39136 12852 39200
rect 12916 39136 12924 39200
rect 12604 38954 12924 39136
rect 12604 38718 12646 38954
rect 12882 38718 12924 38954
rect 12604 38112 12924 38718
rect 12604 38048 12612 38112
rect 12676 38048 12692 38112
rect 12756 38048 12772 38112
rect 12836 38048 12852 38112
rect 12916 38048 12924 38112
rect 12604 37024 12924 38048
rect 12604 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12924 37024
rect 12604 35936 12924 36960
rect 12604 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12924 35936
rect 12604 34848 12924 35872
rect 12604 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12924 34848
rect 12604 33954 12924 34784
rect 12604 33760 12646 33954
rect 12882 33760 12924 33954
rect 12604 33696 12612 33760
rect 12676 33696 12692 33718
rect 12756 33696 12772 33718
rect 12836 33696 12852 33718
rect 12916 33696 12924 33760
rect 12604 32672 12924 33696
rect 12604 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12924 32672
rect 12604 31584 12924 32608
rect 12604 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12924 31584
rect 12604 30496 12924 31520
rect 12604 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12924 30496
rect 12604 29408 12924 30432
rect 12604 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12924 29408
rect 12604 28954 12924 29344
rect 12604 28718 12646 28954
rect 12882 28718 12924 28954
rect 12604 28320 12924 28718
rect 12604 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12924 28320
rect 12604 27232 12924 28256
rect 12604 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12924 27232
rect 12604 26144 12924 27168
rect 12604 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12924 26144
rect 12604 25056 12924 26080
rect 12604 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12924 25056
rect 12604 23968 12924 24992
rect 12604 23904 12612 23968
rect 12676 23954 12692 23968
rect 12756 23954 12772 23968
rect 12836 23954 12852 23968
rect 12916 23904 12924 23968
rect 12604 23718 12646 23904
rect 12882 23718 12924 23904
rect 12604 22880 12924 23718
rect 12604 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12924 22880
rect 12604 21792 12924 22816
rect 12604 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12924 21792
rect 12604 20704 12924 21728
rect 12604 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12924 20704
rect 12604 19616 12924 20640
rect 12604 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12924 19616
rect 12604 18954 12924 19552
rect 12604 18718 12646 18954
rect 12882 18718 12924 18954
rect 12604 18528 12924 18718
rect 12604 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12924 18528
rect 12604 17440 12924 18464
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 16944 57152 17264 57712
rect 16944 57088 16952 57152
rect 17016 57088 17032 57152
rect 17096 57088 17112 57152
rect 17176 57088 17192 57152
rect 17256 57088 17264 57152
rect 16944 56064 17264 57088
rect 16944 56000 16952 56064
rect 17016 56000 17032 56064
rect 17096 56000 17112 56064
rect 17176 56000 17192 56064
rect 17256 56000 17264 56064
rect 16944 54976 17264 56000
rect 16944 54912 16952 54976
rect 17016 54912 17032 54976
rect 17096 54912 17112 54976
rect 17176 54912 17192 54976
rect 17256 54912 17264 54976
rect 16944 53888 17264 54912
rect 16944 53824 16952 53888
rect 17016 53824 17032 53888
rect 17096 53824 17112 53888
rect 17176 53824 17192 53888
rect 17256 53824 17264 53888
rect 16944 53294 17264 53824
rect 16944 53058 16986 53294
rect 17222 53058 17264 53294
rect 16944 52800 17264 53058
rect 16944 52736 16952 52800
rect 17016 52736 17032 52800
rect 17096 52736 17112 52800
rect 17176 52736 17192 52800
rect 17256 52736 17264 52800
rect 16944 51712 17264 52736
rect 16944 51648 16952 51712
rect 17016 51648 17032 51712
rect 17096 51648 17112 51712
rect 17176 51648 17192 51712
rect 17256 51648 17264 51712
rect 16944 50624 17264 51648
rect 16944 50560 16952 50624
rect 17016 50560 17032 50624
rect 17096 50560 17112 50624
rect 17176 50560 17192 50624
rect 17256 50560 17264 50624
rect 16944 49536 17264 50560
rect 16944 49472 16952 49536
rect 17016 49472 17032 49536
rect 17096 49472 17112 49536
rect 17176 49472 17192 49536
rect 17256 49472 17264 49536
rect 16944 48448 17264 49472
rect 16944 48384 16952 48448
rect 17016 48384 17032 48448
rect 17096 48384 17112 48448
rect 17176 48384 17192 48448
rect 17256 48384 17264 48448
rect 16944 48294 17264 48384
rect 16944 48058 16986 48294
rect 17222 48058 17264 48294
rect 16944 47360 17264 48058
rect 16944 47296 16952 47360
rect 17016 47296 17032 47360
rect 17096 47296 17112 47360
rect 17176 47296 17192 47360
rect 17256 47296 17264 47360
rect 16944 46272 17264 47296
rect 16944 46208 16952 46272
rect 17016 46208 17032 46272
rect 17096 46208 17112 46272
rect 17176 46208 17192 46272
rect 17256 46208 17264 46272
rect 16944 45184 17264 46208
rect 16944 45120 16952 45184
rect 17016 45120 17032 45184
rect 17096 45120 17112 45184
rect 17176 45120 17192 45184
rect 17256 45120 17264 45184
rect 16944 44096 17264 45120
rect 16944 44032 16952 44096
rect 17016 44032 17032 44096
rect 17096 44032 17112 44096
rect 17176 44032 17192 44096
rect 17256 44032 17264 44096
rect 16944 43294 17264 44032
rect 16944 43058 16986 43294
rect 17222 43058 17264 43294
rect 16944 43008 17264 43058
rect 16944 42944 16952 43008
rect 17016 42944 17032 43008
rect 17096 42944 17112 43008
rect 17176 42944 17192 43008
rect 17256 42944 17264 43008
rect 16944 41920 17264 42944
rect 16944 41856 16952 41920
rect 17016 41856 17032 41920
rect 17096 41856 17112 41920
rect 17176 41856 17192 41920
rect 17256 41856 17264 41920
rect 16944 40832 17264 41856
rect 16944 40768 16952 40832
rect 17016 40768 17032 40832
rect 17096 40768 17112 40832
rect 17176 40768 17192 40832
rect 17256 40768 17264 40832
rect 16944 39744 17264 40768
rect 16944 39680 16952 39744
rect 17016 39680 17032 39744
rect 17096 39680 17112 39744
rect 17176 39680 17192 39744
rect 17256 39680 17264 39744
rect 16944 38656 17264 39680
rect 16944 38592 16952 38656
rect 17016 38592 17032 38656
rect 17096 38592 17112 38656
rect 17176 38592 17192 38656
rect 17256 38592 17264 38656
rect 16944 38294 17264 38592
rect 16944 38058 16986 38294
rect 17222 38058 17264 38294
rect 16944 37568 17264 38058
rect 16944 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17264 37568
rect 16944 36480 17264 37504
rect 16944 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17264 36480
rect 16944 35392 17264 36416
rect 16944 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17264 35392
rect 16944 34304 17264 35328
rect 16944 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17264 34304
rect 16944 33294 17264 34240
rect 16944 33216 16986 33294
rect 17222 33216 17264 33294
rect 16944 33152 16952 33216
rect 17256 33152 17264 33216
rect 16944 33058 16986 33152
rect 17222 33058 17264 33152
rect 16944 32128 17264 33058
rect 16944 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17264 32128
rect 16944 31040 17264 32064
rect 16944 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17264 31040
rect 16944 29952 17264 30976
rect 16944 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17264 29952
rect 16944 28864 17264 29888
rect 16944 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17264 28864
rect 16944 28294 17264 28800
rect 16944 28058 16986 28294
rect 17222 28058 17264 28294
rect 16944 27776 17264 28058
rect 16944 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17264 27776
rect 16944 26688 17264 27712
rect 16944 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17264 26688
rect 16944 25600 17264 26624
rect 16944 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17264 25600
rect 16944 24512 17264 25536
rect 16944 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17264 24512
rect 16944 23424 17264 24448
rect 16944 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17264 23424
rect 16944 23294 17264 23360
rect 16944 23058 16986 23294
rect 17222 23058 17264 23294
rect 16944 22336 17264 23058
rect 16944 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17264 22336
rect 16944 21248 17264 22272
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 18294 17264 19008
rect 16944 18058 16986 18294
rect 17222 18058 17264 18294
rect 16944 17984 17264 18058
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16944 12544 17264 13058
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 17604 57696 17924 57712
rect 17604 57632 17612 57696
rect 17676 57632 17692 57696
rect 17756 57632 17772 57696
rect 17836 57632 17852 57696
rect 17916 57632 17924 57696
rect 17604 56608 17924 57632
rect 17604 56544 17612 56608
rect 17676 56544 17692 56608
rect 17756 56544 17772 56608
rect 17836 56544 17852 56608
rect 17916 56544 17924 56608
rect 17604 55520 17924 56544
rect 17604 55456 17612 55520
rect 17676 55456 17692 55520
rect 17756 55456 17772 55520
rect 17836 55456 17852 55520
rect 17916 55456 17924 55520
rect 17604 54432 17924 55456
rect 17604 54368 17612 54432
rect 17676 54368 17692 54432
rect 17756 54368 17772 54432
rect 17836 54368 17852 54432
rect 17916 54368 17924 54432
rect 17604 53954 17924 54368
rect 17604 53718 17646 53954
rect 17882 53718 17924 53954
rect 17604 53344 17924 53718
rect 17604 53280 17612 53344
rect 17676 53280 17692 53344
rect 17756 53280 17772 53344
rect 17836 53280 17852 53344
rect 17916 53280 17924 53344
rect 17604 52256 17924 53280
rect 17604 52192 17612 52256
rect 17676 52192 17692 52256
rect 17756 52192 17772 52256
rect 17836 52192 17852 52256
rect 17916 52192 17924 52256
rect 17604 51168 17924 52192
rect 17604 51104 17612 51168
rect 17676 51104 17692 51168
rect 17756 51104 17772 51168
rect 17836 51104 17852 51168
rect 17916 51104 17924 51168
rect 17604 50080 17924 51104
rect 17604 50016 17612 50080
rect 17676 50016 17692 50080
rect 17756 50016 17772 50080
rect 17836 50016 17852 50080
rect 17916 50016 17924 50080
rect 17604 48992 17924 50016
rect 17604 48928 17612 48992
rect 17676 48954 17692 48992
rect 17756 48954 17772 48992
rect 17836 48954 17852 48992
rect 17916 48928 17924 48992
rect 17604 48718 17646 48928
rect 17882 48718 17924 48928
rect 17604 47904 17924 48718
rect 17604 47840 17612 47904
rect 17676 47840 17692 47904
rect 17756 47840 17772 47904
rect 17836 47840 17852 47904
rect 17916 47840 17924 47904
rect 17604 46816 17924 47840
rect 17604 46752 17612 46816
rect 17676 46752 17692 46816
rect 17756 46752 17772 46816
rect 17836 46752 17852 46816
rect 17916 46752 17924 46816
rect 17604 45728 17924 46752
rect 17604 45664 17612 45728
rect 17676 45664 17692 45728
rect 17756 45664 17772 45728
rect 17836 45664 17852 45728
rect 17916 45664 17924 45728
rect 17604 44640 17924 45664
rect 17604 44576 17612 44640
rect 17676 44576 17692 44640
rect 17756 44576 17772 44640
rect 17836 44576 17852 44640
rect 17916 44576 17924 44640
rect 17604 43954 17924 44576
rect 17604 43718 17646 43954
rect 17882 43718 17924 43954
rect 17604 43552 17924 43718
rect 17604 43488 17612 43552
rect 17676 43488 17692 43552
rect 17756 43488 17772 43552
rect 17836 43488 17852 43552
rect 17916 43488 17924 43552
rect 17604 42464 17924 43488
rect 17604 42400 17612 42464
rect 17676 42400 17692 42464
rect 17756 42400 17772 42464
rect 17836 42400 17852 42464
rect 17916 42400 17924 42464
rect 17604 41376 17924 42400
rect 17604 41312 17612 41376
rect 17676 41312 17692 41376
rect 17756 41312 17772 41376
rect 17836 41312 17852 41376
rect 17916 41312 17924 41376
rect 17604 40288 17924 41312
rect 17604 40224 17612 40288
rect 17676 40224 17692 40288
rect 17756 40224 17772 40288
rect 17836 40224 17852 40288
rect 17916 40224 17924 40288
rect 17604 39200 17924 40224
rect 17604 39136 17612 39200
rect 17676 39136 17692 39200
rect 17756 39136 17772 39200
rect 17836 39136 17852 39200
rect 17916 39136 17924 39200
rect 17604 38954 17924 39136
rect 17604 38718 17646 38954
rect 17882 38718 17924 38954
rect 17604 38112 17924 38718
rect 17604 38048 17612 38112
rect 17676 38048 17692 38112
rect 17756 38048 17772 38112
rect 17836 38048 17852 38112
rect 17916 38048 17924 38112
rect 17604 37024 17924 38048
rect 17604 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17924 37024
rect 17604 35936 17924 36960
rect 17604 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17924 35936
rect 17604 34848 17924 35872
rect 17604 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17924 34848
rect 17604 33954 17924 34784
rect 17604 33760 17646 33954
rect 17882 33760 17924 33954
rect 17604 33696 17612 33760
rect 17676 33696 17692 33718
rect 17756 33696 17772 33718
rect 17836 33696 17852 33718
rect 17916 33696 17924 33760
rect 17604 32672 17924 33696
rect 17604 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17924 32672
rect 17604 31584 17924 32608
rect 17604 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17924 31584
rect 17604 30496 17924 31520
rect 17604 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17924 30496
rect 17604 29408 17924 30432
rect 17604 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17924 29408
rect 17604 28954 17924 29344
rect 17604 28718 17646 28954
rect 17882 28718 17924 28954
rect 17604 28320 17924 28718
rect 17604 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17924 28320
rect 17604 27232 17924 28256
rect 17604 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17924 27232
rect 17604 26144 17924 27168
rect 17604 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17924 26144
rect 17604 25056 17924 26080
rect 17604 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17924 25056
rect 17604 23968 17924 24992
rect 17604 23904 17612 23968
rect 17676 23954 17692 23968
rect 17756 23954 17772 23968
rect 17836 23954 17852 23968
rect 17916 23904 17924 23968
rect 17604 23718 17646 23904
rect 17882 23718 17924 23904
rect 17604 22880 17924 23718
rect 17604 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17924 22880
rect 17604 21792 17924 22816
rect 17604 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17924 21792
rect 17604 20704 17924 21728
rect 17604 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17924 20704
rect 17604 19616 17924 20640
rect 17604 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17924 19616
rect 17604 18954 17924 19552
rect 17604 18718 17646 18954
rect 17882 18718 17924 18954
rect 17604 18528 17924 18718
rect 17604 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17924 18528
rect 17604 17440 17924 18464
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17604 12000 17924 13024
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
rect 21944 57152 22264 57712
rect 21944 57088 21952 57152
rect 22016 57088 22032 57152
rect 22096 57088 22112 57152
rect 22176 57088 22192 57152
rect 22256 57088 22264 57152
rect 21944 56064 22264 57088
rect 21944 56000 21952 56064
rect 22016 56000 22032 56064
rect 22096 56000 22112 56064
rect 22176 56000 22192 56064
rect 22256 56000 22264 56064
rect 21944 54976 22264 56000
rect 21944 54912 21952 54976
rect 22016 54912 22032 54976
rect 22096 54912 22112 54976
rect 22176 54912 22192 54976
rect 22256 54912 22264 54976
rect 21944 53888 22264 54912
rect 21944 53824 21952 53888
rect 22016 53824 22032 53888
rect 22096 53824 22112 53888
rect 22176 53824 22192 53888
rect 22256 53824 22264 53888
rect 21944 53294 22264 53824
rect 21944 53058 21986 53294
rect 22222 53058 22264 53294
rect 21944 52800 22264 53058
rect 21944 52736 21952 52800
rect 22016 52736 22032 52800
rect 22096 52736 22112 52800
rect 22176 52736 22192 52800
rect 22256 52736 22264 52800
rect 21944 51712 22264 52736
rect 21944 51648 21952 51712
rect 22016 51648 22032 51712
rect 22096 51648 22112 51712
rect 22176 51648 22192 51712
rect 22256 51648 22264 51712
rect 21944 50624 22264 51648
rect 21944 50560 21952 50624
rect 22016 50560 22032 50624
rect 22096 50560 22112 50624
rect 22176 50560 22192 50624
rect 22256 50560 22264 50624
rect 21944 49536 22264 50560
rect 21944 49472 21952 49536
rect 22016 49472 22032 49536
rect 22096 49472 22112 49536
rect 22176 49472 22192 49536
rect 22256 49472 22264 49536
rect 21944 48448 22264 49472
rect 21944 48384 21952 48448
rect 22016 48384 22032 48448
rect 22096 48384 22112 48448
rect 22176 48384 22192 48448
rect 22256 48384 22264 48448
rect 21944 48294 22264 48384
rect 21944 48058 21986 48294
rect 22222 48058 22264 48294
rect 21944 47360 22264 48058
rect 21944 47296 21952 47360
rect 22016 47296 22032 47360
rect 22096 47296 22112 47360
rect 22176 47296 22192 47360
rect 22256 47296 22264 47360
rect 21944 46272 22264 47296
rect 21944 46208 21952 46272
rect 22016 46208 22032 46272
rect 22096 46208 22112 46272
rect 22176 46208 22192 46272
rect 22256 46208 22264 46272
rect 21944 45184 22264 46208
rect 21944 45120 21952 45184
rect 22016 45120 22032 45184
rect 22096 45120 22112 45184
rect 22176 45120 22192 45184
rect 22256 45120 22264 45184
rect 21944 44096 22264 45120
rect 21944 44032 21952 44096
rect 22016 44032 22032 44096
rect 22096 44032 22112 44096
rect 22176 44032 22192 44096
rect 22256 44032 22264 44096
rect 21944 43294 22264 44032
rect 21944 43058 21986 43294
rect 22222 43058 22264 43294
rect 21944 43008 22264 43058
rect 21944 42944 21952 43008
rect 22016 42944 22032 43008
rect 22096 42944 22112 43008
rect 22176 42944 22192 43008
rect 22256 42944 22264 43008
rect 21944 41920 22264 42944
rect 21944 41856 21952 41920
rect 22016 41856 22032 41920
rect 22096 41856 22112 41920
rect 22176 41856 22192 41920
rect 22256 41856 22264 41920
rect 21944 40832 22264 41856
rect 21944 40768 21952 40832
rect 22016 40768 22032 40832
rect 22096 40768 22112 40832
rect 22176 40768 22192 40832
rect 22256 40768 22264 40832
rect 21944 39744 22264 40768
rect 21944 39680 21952 39744
rect 22016 39680 22032 39744
rect 22096 39680 22112 39744
rect 22176 39680 22192 39744
rect 22256 39680 22264 39744
rect 21944 38656 22264 39680
rect 21944 38592 21952 38656
rect 22016 38592 22032 38656
rect 22096 38592 22112 38656
rect 22176 38592 22192 38656
rect 22256 38592 22264 38656
rect 21944 38294 22264 38592
rect 21944 38058 21986 38294
rect 22222 38058 22264 38294
rect 21944 37568 22264 38058
rect 21944 37504 21952 37568
rect 22016 37504 22032 37568
rect 22096 37504 22112 37568
rect 22176 37504 22192 37568
rect 22256 37504 22264 37568
rect 21944 36480 22264 37504
rect 21944 36416 21952 36480
rect 22016 36416 22032 36480
rect 22096 36416 22112 36480
rect 22176 36416 22192 36480
rect 22256 36416 22264 36480
rect 21944 35392 22264 36416
rect 21944 35328 21952 35392
rect 22016 35328 22032 35392
rect 22096 35328 22112 35392
rect 22176 35328 22192 35392
rect 22256 35328 22264 35392
rect 21944 34304 22264 35328
rect 21944 34240 21952 34304
rect 22016 34240 22032 34304
rect 22096 34240 22112 34304
rect 22176 34240 22192 34304
rect 22256 34240 22264 34304
rect 21944 33294 22264 34240
rect 21944 33216 21986 33294
rect 22222 33216 22264 33294
rect 21944 33152 21952 33216
rect 22256 33152 22264 33216
rect 21944 33058 21986 33152
rect 22222 33058 22264 33152
rect 21944 32128 22264 33058
rect 21944 32064 21952 32128
rect 22016 32064 22032 32128
rect 22096 32064 22112 32128
rect 22176 32064 22192 32128
rect 22256 32064 22264 32128
rect 21944 31040 22264 32064
rect 21944 30976 21952 31040
rect 22016 30976 22032 31040
rect 22096 30976 22112 31040
rect 22176 30976 22192 31040
rect 22256 30976 22264 31040
rect 21944 29952 22264 30976
rect 21944 29888 21952 29952
rect 22016 29888 22032 29952
rect 22096 29888 22112 29952
rect 22176 29888 22192 29952
rect 22256 29888 22264 29952
rect 21944 28864 22264 29888
rect 21944 28800 21952 28864
rect 22016 28800 22032 28864
rect 22096 28800 22112 28864
rect 22176 28800 22192 28864
rect 22256 28800 22264 28864
rect 21944 28294 22264 28800
rect 21944 28058 21986 28294
rect 22222 28058 22264 28294
rect 21944 27776 22264 28058
rect 21944 27712 21952 27776
rect 22016 27712 22032 27776
rect 22096 27712 22112 27776
rect 22176 27712 22192 27776
rect 22256 27712 22264 27776
rect 21944 26688 22264 27712
rect 21944 26624 21952 26688
rect 22016 26624 22032 26688
rect 22096 26624 22112 26688
rect 22176 26624 22192 26688
rect 22256 26624 22264 26688
rect 21944 25600 22264 26624
rect 21944 25536 21952 25600
rect 22016 25536 22032 25600
rect 22096 25536 22112 25600
rect 22176 25536 22192 25600
rect 22256 25536 22264 25600
rect 21944 24512 22264 25536
rect 21944 24448 21952 24512
rect 22016 24448 22032 24512
rect 22096 24448 22112 24512
rect 22176 24448 22192 24512
rect 22256 24448 22264 24512
rect 21944 23424 22264 24448
rect 21944 23360 21952 23424
rect 22016 23360 22032 23424
rect 22096 23360 22112 23424
rect 22176 23360 22192 23424
rect 22256 23360 22264 23424
rect 21944 23294 22264 23360
rect 21944 23058 21986 23294
rect 22222 23058 22264 23294
rect 21944 22336 22264 23058
rect 21944 22272 21952 22336
rect 22016 22272 22032 22336
rect 22096 22272 22112 22336
rect 22176 22272 22192 22336
rect 22256 22272 22264 22336
rect 21944 21248 22264 22272
rect 21944 21184 21952 21248
rect 22016 21184 22032 21248
rect 22096 21184 22112 21248
rect 22176 21184 22192 21248
rect 22256 21184 22264 21248
rect 21944 20160 22264 21184
rect 21944 20096 21952 20160
rect 22016 20096 22032 20160
rect 22096 20096 22112 20160
rect 22176 20096 22192 20160
rect 22256 20096 22264 20160
rect 21944 19072 22264 20096
rect 21944 19008 21952 19072
rect 22016 19008 22032 19072
rect 22096 19008 22112 19072
rect 22176 19008 22192 19072
rect 22256 19008 22264 19072
rect 21944 18294 22264 19008
rect 21944 18058 21986 18294
rect 22222 18058 22264 18294
rect 21944 17984 22264 18058
rect 21944 17920 21952 17984
rect 22016 17920 22032 17984
rect 22096 17920 22112 17984
rect 22176 17920 22192 17984
rect 22256 17920 22264 17984
rect 21944 16896 22264 17920
rect 21944 16832 21952 16896
rect 22016 16832 22032 16896
rect 22096 16832 22112 16896
rect 22176 16832 22192 16896
rect 22256 16832 22264 16896
rect 21944 15808 22264 16832
rect 21944 15744 21952 15808
rect 22016 15744 22032 15808
rect 22096 15744 22112 15808
rect 22176 15744 22192 15808
rect 22256 15744 22264 15808
rect 21944 14720 22264 15744
rect 21944 14656 21952 14720
rect 22016 14656 22032 14720
rect 22096 14656 22112 14720
rect 22176 14656 22192 14720
rect 22256 14656 22264 14720
rect 21944 13632 22264 14656
rect 21944 13568 21952 13632
rect 22016 13568 22032 13632
rect 22096 13568 22112 13632
rect 22176 13568 22192 13632
rect 22256 13568 22264 13632
rect 21944 13294 22264 13568
rect 21944 13058 21986 13294
rect 22222 13058 22264 13294
rect 21944 12544 22264 13058
rect 21944 12480 21952 12544
rect 22016 12480 22032 12544
rect 22096 12480 22112 12544
rect 22176 12480 22192 12544
rect 22256 12480 22264 12544
rect 21944 11456 22264 12480
rect 21944 11392 21952 11456
rect 22016 11392 22032 11456
rect 22096 11392 22112 11456
rect 22176 11392 22192 11456
rect 22256 11392 22264 11456
rect 21944 10368 22264 11392
rect 21944 10304 21952 10368
rect 22016 10304 22032 10368
rect 22096 10304 22112 10368
rect 22176 10304 22192 10368
rect 22256 10304 22264 10368
rect 21944 9280 22264 10304
rect 21944 9216 21952 9280
rect 22016 9216 22032 9280
rect 22096 9216 22112 9280
rect 22176 9216 22192 9280
rect 22256 9216 22264 9280
rect 21944 8294 22264 9216
rect 21944 8192 21986 8294
rect 22222 8192 22264 8294
rect 21944 8128 21952 8192
rect 22256 8128 22264 8192
rect 21944 8058 21986 8128
rect 22222 8058 22264 8128
rect 21944 7104 22264 8058
rect 21944 7040 21952 7104
rect 22016 7040 22032 7104
rect 22096 7040 22112 7104
rect 22176 7040 22192 7104
rect 22256 7040 22264 7104
rect 21944 6016 22264 7040
rect 21944 5952 21952 6016
rect 22016 5952 22032 6016
rect 22096 5952 22112 6016
rect 22176 5952 22192 6016
rect 22256 5952 22264 6016
rect 21944 4928 22264 5952
rect 21944 4864 21952 4928
rect 22016 4864 22032 4928
rect 22096 4864 22112 4928
rect 22176 4864 22192 4928
rect 22256 4864 22264 4928
rect 21944 3840 22264 4864
rect 21944 3776 21952 3840
rect 22016 3776 22032 3840
rect 22096 3776 22112 3840
rect 22176 3776 22192 3840
rect 22256 3776 22264 3840
rect 21944 3294 22264 3776
rect 21944 3058 21986 3294
rect 22222 3058 22264 3294
rect 21944 2752 22264 3058
rect 21944 2688 21952 2752
rect 22016 2688 22032 2752
rect 22096 2688 22112 2752
rect 22176 2688 22192 2752
rect 22256 2688 22264 2752
rect 21944 2128 22264 2688
rect 22604 57696 22924 57712
rect 22604 57632 22612 57696
rect 22676 57632 22692 57696
rect 22756 57632 22772 57696
rect 22836 57632 22852 57696
rect 22916 57632 22924 57696
rect 22604 56608 22924 57632
rect 22604 56544 22612 56608
rect 22676 56544 22692 56608
rect 22756 56544 22772 56608
rect 22836 56544 22852 56608
rect 22916 56544 22924 56608
rect 22604 55520 22924 56544
rect 22604 55456 22612 55520
rect 22676 55456 22692 55520
rect 22756 55456 22772 55520
rect 22836 55456 22852 55520
rect 22916 55456 22924 55520
rect 22604 54432 22924 55456
rect 22604 54368 22612 54432
rect 22676 54368 22692 54432
rect 22756 54368 22772 54432
rect 22836 54368 22852 54432
rect 22916 54368 22924 54432
rect 22604 53954 22924 54368
rect 22604 53718 22646 53954
rect 22882 53718 22924 53954
rect 22604 53344 22924 53718
rect 22604 53280 22612 53344
rect 22676 53280 22692 53344
rect 22756 53280 22772 53344
rect 22836 53280 22852 53344
rect 22916 53280 22924 53344
rect 22604 52256 22924 53280
rect 22604 52192 22612 52256
rect 22676 52192 22692 52256
rect 22756 52192 22772 52256
rect 22836 52192 22852 52256
rect 22916 52192 22924 52256
rect 22604 51168 22924 52192
rect 22604 51104 22612 51168
rect 22676 51104 22692 51168
rect 22756 51104 22772 51168
rect 22836 51104 22852 51168
rect 22916 51104 22924 51168
rect 22604 50080 22924 51104
rect 22604 50016 22612 50080
rect 22676 50016 22692 50080
rect 22756 50016 22772 50080
rect 22836 50016 22852 50080
rect 22916 50016 22924 50080
rect 22604 48992 22924 50016
rect 22604 48928 22612 48992
rect 22676 48954 22692 48992
rect 22756 48954 22772 48992
rect 22836 48954 22852 48992
rect 22916 48928 22924 48992
rect 22604 48718 22646 48928
rect 22882 48718 22924 48928
rect 22604 47904 22924 48718
rect 22604 47840 22612 47904
rect 22676 47840 22692 47904
rect 22756 47840 22772 47904
rect 22836 47840 22852 47904
rect 22916 47840 22924 47904
rect 22604 46816 22924 47840
rect 22604 46752 22612 46816
rect 22676 46752 22692 46816
rect 22756 46752 22772 46816
rect 22836 46752 22852 46816
rect 22916 46752 22924 46816
rect 22604 45728 22924 46752
rect 22604 45664 22612 45728
rect 22676 45664 22692 45728
rect 22756 45664 22772 45728
rect 22836 45664 22852 45728
rect 22916 45664 22924 45728
rect 22604 44640 22924 45664
rect 22604 44576 22612 44640
rect 22676 44576 22692 44640
rect 22756 44576 22772 44640
rect 22836 44576 22852 44640
rect 22916 44576 22924 44640
rect 22604 43954 22924 44576
rect 22604 43718 22646 43954
rect 22882 43718 22924 43954
rect 22604 43552 22924 43718
rect 22604 43488 22612 43552
rect 22676 43488 22692 43552
rect 22756 43488 22772 43552
rect 22836 43488 22852 43552
rect 22916 43488 22924 43552
rect 22604 42464 22924 43488
rect 22604 42400 22612 42464
rect 22676 42400 22692 42464
rect 22756 42400 22772 42464
rect 22836 42400 22852 42464
rect 22916 42400 22924 42464
rect 22604 41376 22924 42400
rect 22604 41312 22612 41376
rect 22676 41312 22692 41376
rect 22756 41312 22772 41376
rect 22836 41312 22852 41376
rect 22916 41312 22924 41376
rect 22604 40288 22924 41312
rect 22604 40224 22612 40288
rect 22676 40224 22692 40288
rect 22756 40224 22772 40288
rect 22836 40224 22852 40288
rect 22916 40224 22924 40288
rect 22604 39200 22924 40224
rect 22604 39136 22612 39200
rect 22676 39136 22692 39200
rect 22756 39136 22772 39200
rect 22836 39136 22852 39200
rect 22916 39136 22924 39200
rect 22604 38954 22924 39136
rect 22604 38718 22646 38954
rect 22882 38718 22924 38954
rect 22604 38112 22924 38718
rect 22604 38048 22612 38112
rect 22676 38048 22692 38112
rect 22756 38048 22772 38112
rect 22836 38048 22852 38112
rect 22916 38048 22924 38112
rect 22604 37024 22924 38048
rect 22604 36960 22612 37024
rect 22676 36960 22692 37024
rect 22756 36960 22772 37024
rect 22836 36960 22852 37024
rect 22916 36960 22924 37024
rect 22604 35936 22924 36960
rect 22604 35872 22612 35936
rect 22676 35872 22692 35936
rect 22756 35872 22772 35936
rect 22836 35872 22852 35936
rect 22916 35872 22924 35936
rect 22604 34848 22924 35872
rect 22604 34784 22612 34848
rect 22676 34784 22692 34848
rect 22756 34784 22772 34848
rect 22836 34784 22852 34848
rect 22916 34784 22924 34848
rect 22604 33954 22924 34784
rect 22604 33760 22646 33954
rect 22882 33760 22924 33954
rect 22604 33696 22612 33760
rect 22676 33696 22692 33718
rect 22756 33696 22772 33718
rect 22836 33696 22852 33718
rect 22916 33696 22924 33760
rect 22604 32672 22924 33696
rect 22604 32608 22612 32672
rect 22676 32608 22692 32672
rect 22756 32608 22772 32672
rect 22836 32608 22852 32672
rect 22916 32608 22924 32672
rect 22604 31584 22924 32608
rect 22604 31520 22612 31584
rect 22676 31520 22692 31584
rect 22756 31520 22772 31584
rect 22836 31520 22852 31584
rect 22916 31520 22924 31584
rect 22604 30496 22924 31520
rect 22604 30432 22612 30496
rect 22676 30432 22692 30496
rect 22756 30432 22772 30496
rect 22836 30432 22852 30496
rect 22916 30432 22924 30496
rect 22604 29408 22924 30432
rect 22604 29344 22612 29408
rect 22676 29344 22692 29408
rect 22756 29344 22772 29408
rect 22836 29344 22852 29408
rect 22916 29344 22924 29408
rect 22604 28954 22924 29344
rect 22604 28718 22646 28954
rect 22882 28718 22924 28954
rect 22604 28320 22924 28718
rect 22604 28256 22612 28320
rect 22676 28256 22692 28320
rect 22756 28256 22772 28320
rect 22836 28256 22852 28320
rect 22916 28256 22924 28320
rect 22604 27232 22924 28256
rect 22604 27168 22612 27232
rect 22676 27168 22692 27232
rect 22756 27168 22772 27232
rect 22836 27168 22852 27232
rect 22916 27168 22924 27232
rect 22604 26144 22924 27168
rect 22604 26080 22612 26144
rect 22676 26080 22692 26144
rect 22756 26080 22772 26144
rect 22836 26080 22852 26144
rect 22916 26080 22924 26144
rect 22604 25056 22924 26080
rect 22604 24992 22612 25056
rect 22676 24992 22692 25056
rect 22756 24992 22772 25056
rect 22836 24992 22852 25056
rect 22916 24992 22924 25056
rect 22604 23968 22924 24992
rect 22604 23904 22612 23968
rect 22676 23954 22692 23968
rect 22756 23954 22772 23968
rect 22836 23954 22852 23968
rect 22916 23904 22924 23968
rect 22604 23718 22646 23904
rect 22882 23718 22924 23904
rect 22604 22880 22924 23718
rect 22604 22816 22612 22880
rect 22676 22816 22692 22880
rect 22756 22816 22772 22880
rect 22836 22816 22852 22880
rect 22916 22816 22924 22880
rect 22604 21792 22924 22816
rect 22604 21728 22612 21792
rect 22676 21728 22692 21792
rect 22756 21728 22772 21792
rect 22836 21728 22852 21792
rect 22916 21728 22924 21792
rect 22604 20704 22924 21728
rect 22604 20640 22612 20704
rect 22676 20640 22692 20704
rect 22756 20640 22772 20704
rect 22836 20640 22852 20704
rect 22916 20640 22924 20704
rect 22604 19616 22924 20640
rect 22604 19552 22612 19616
rect 22676 19552 22692 19616
rect 22756 19552 22772 19616
rect 22836 19552 22852 19616
rect 22916 19552 22924 19616
rect 22604 18954 22924 19552
rect 22604 18718 22646 18954
rect 22882 18718 22924 18954
rect 22604 18528 22924 18718
rect 22604 18464 22612 18528
rect 22676 18464 22692 18528
rect 22756 18464 22772 18528
rect 22836 18464 22852 18528
rect 22916 18464 22924 18528
rect 22604 17440 22924 18464
rect 22604 17376 22612 17440
rect 22676 17376 22692 17440
rect 22756 17376 22772 17440
rect 22836 17376 22852 17440
rect 22916 17376 22924 17440
rect 22604 16352 22924 17376
rect 22604 16288 22612 16352
rect 22676 16288 22692 16352
rect 22756 16288 22772 16352
rect 22836 16288 22852 16352
rect 22916 16288 22924 16352
rect 22604 15264 22924 16288
rect 22604 15200 22612 15264
rect 22676 15200 22692 15264
rect 22756 15200 22772 15264
rect 22836 15200 22852 15264
rect 22916 15200 22924 15264
rect 22604 14176 22924 15200
rect 22604 14112 22612 14176
rect 22676 14112 22692 14176
rect 22756 14112 22772 14176
rect 22836 14112 22852 14176
rect 22916 14112 22924 14176
rect 22604 13954 22924 14112
rect 22604 13718 22646 13954
rect 22882 13718 22924 13954
rect 22604 13088 22924 13718
rect 22604 13024 22612 13088
rect 22676 13024 22692 13088
rect 22756 13024 22772 13088
rect 22836 13024 22852 13088
rect 22916 13024 22924 13088
rect 22604 12000 22924 13024
rect 22604 11936 22612 12000
rect 22676 11936 22692 12000
rect 22756 11936 22772 12000
rect 22836 11936 22852 12000
rect 22916 11936 22924 12000
rect 22604 10912 22924 11936
rect 22604 10848 22612 10912
rect 22676 10848 22692 10912
rect 22756 10848 22772 10912
rect 22836 10848 22852 10912
rect 22916 10848 22924 10912
rect 22604 9824 22924 10848
rect 22604 9760 22612 9824
rect 22676 9760 22692 9824
rect 22756 9760 22772 9824
rect 22836 9760 22852 9824
rect 22916 9760 22924 9824
rect 22604 8954 22924 9760
rect 22604 8736 22646 8954
rect 22882 8736 22924 8954
rect 22604 8672 22612 8736
rect 22676 8672 22692 8718
rect 22756 8672 22772 8718
rect 22836 8672 22852 8718
rect 22916 8672 22924 8736
rect 22604 7648 22924 8672
rect 22604 7584 22612 7648
rect 22676 7584 22692 7648
rect 22756 7584 22772 7648
rect 22836 7584 22852 7648
rect 22916 7584 22924 7648
rect 22604 6560 22924 7584
rect 22604 6496 22612 6560
rect 22676 6496 22692 6560
rect 22756 6496 22772 6560
rect 22836 6496 22852 6560
rect 22916 6496 22924 6560
rect 22604 5472 22924 6496
rect 22604 5408 22612 5472
rect 22676 5408 22692 5472
rect 22756 5408 22772 5472
rect 22836 5408 22852 5472
rect 22916 5408 22924 5472
rect 22604 4384 22924 5408
rect 22604 4320 22612 4384
rect 22676 4320 22692 4384
rect 22756 4320 22772 4384
rect 22836 4320 22852 4384
rect 22916 4320 22924 4384
rect 22604 3954 22924 4320
rect 22604 3718 22646 3954
rect 22882 3718 22924 3954
rect 22604 3296 22924 3718
rect 22604 3232 22612 3296
rect 22676 3232 22692 3296
rect 22756 3232 22772 3296
rect 22836 3232 22852 3296
rect 22916 3232 22924 3296
rect 22604 2208 22924 3232
rect 22604 2144 22612 2208
rect 22676 2144 22692 2208
rect 22756 2144 22772 2208
rect 22836 2144 22852 2208
rect 22916 2144 22924 2208
rect 22604 2128 22924 2144
rect 26944 57152 27264 57712
rect 26944 57088 26952 57152
rect 27016 57088 27032 57152
rect 27096 57088 27112 57152
rect 27176 57088 27192 57152
rect 27256 57088 27264 57152
rect 26944 56064 27264 57088
rect 26944 56000 26952 56064
rect 27016 56000 27032 56064
rect 27096 56000 27112 56064
rect 27176 56000 27192 56064
rect 27256 56000 27264 56064
rect 26944 54976 27264 56000
rect 26944 54912 26952 54976
rect 27016 54912 27032 54976
rect 27096 54912 27112 54976
rect 27176 54912 27192 54976
rect 27256 54912 27264 54976
rect 26944 53888 27264 54912
rect 26944 53824 26952 53888
rect 27016 53824 27032 53888
rect 27096 53824 27112 53888
rect 27176 53824 27192 53888
rect 27256 53824 27264 53888
rect 26944 53294 27264 53824
rect 26944 53058 26986 53294
rect 27222 53058 27264 53294
rect 26944 52800 27264 53058
rect 26944 52736 26952 52800
rect 27016 52736 27032 52800
rect 27096 52736 27112 52800
rect 27176 52736 27192 52800
rect 27256 52736 27264 52800
rect 26944 51712 27264 52736
rect 26944 51648 26952 51712
rect 27016 51648 27032 51712
rect 27096 51648 27112 51712
rect 27176 51648 27192 51712
rect 27256 51648 27264 51712
rect 26944 50624 27264 51648
rect 26944 50560 26952 50624
rect 27016 50560 27032 50624
rect 27096 50560 27112 50624
rect 27176 50560 27192 50624
rect 27256 50560 27264 50624
rect 26944 49536 27264 50560
rect 26944 49472 26952 49536
rect 27016 49472 27032 49536
rect 27096 49472 27112 49536
rect 27176 49472 27192 49536
rect 27256 49472 27264 49536
rect 26944 48448 27264 49472
rect 26944 48384 26952 48448
rect 27016 48384 27032 48448
rect 27096 48384 27112 48448
rect 27176 48384 27192 48448
rect 27256 48384 27264 48448
rect 26944 48294 27264 48384
rect 26944 48058 26986 48294
rect 27222 48058 27264 48294
rect 26944 47360 27264 48058
rect 26944 47296 26952 47360
rect 27016 47296 27032 47360
rect 27096 47296 27112 47360
rect 27176 47296 27192 47360
rect 27256 47296 27264 47360
rect 26944 46272 27264 47296
rect 26944 46208 26952 46272
rect 27016 46208 27032 46272
rect 27096 46208 27112 46272
rect 27176 46208 27192 46272
rect 27256 46208 27264 46272
rect 26944 45184 27264 46208
rect 26944 45120 26952 45184
rect 27016 45120 27032 45184
rect 27096 45120 27112 45184
rect 27176 45120 27192 45184
rect 27256 45120 27264 45184
rect 26944 44096 27264 45120
rect 26944 44032 26952 44096
rect 27016 44032 27032 44096
rect 27096 44032 27112 44096
rect 27176 44032 27192 44096
rect 27256 44032 27264 44096
rect 26944 43294 27264 44032
rect 26944 43058 26986 43294
rect 27222 43058 27264 43294
rect 26944 43008 27264 43058
rect 26944 42944 26952 43008
rect 27016 42944 27032 43008
rect 27096 42944 27112 43008
rect 27176 42944 27192 43008
rect 27256 42944 27264 43008
rect 26944 41920 27264 42944
rect 26944 41856 26952 41920
rect 27016 41856 27032 41920
rect 27096 41856 27112 41920
rect 27176 41856 27192 41920
rect 27256 41856 27264 41920
rect 26944 40832 27264 41856
rect 26944 40768 26952 40832
rect 27016 40768 27032 40832
rect 27096 40768 27112 40832
rect 27176 40768 27192 40832
rect 27256 40768 27264 40832
rect 26944 39744 27264 40768
rect 26944 39680 26952 39744
rect 27016 39680 27032 39744
rect 27096 39680 27112 39744
rect 27176 39680 27192 39744
rect 27256 39680 27264 39744
rect 26944 38656 27264 39680
rect 26944 38592 26952 38656
rect 27016 38592 27032 38656
rect 27096 38592 27112 38656
rect 27176 38592 27192 38656
rect 27256 38592 27264 38656
rect 26944 38294 27264 38592
rect 26944 38058 26986 38294
rect 27222 38058 27264 38294
rect 26944 37568 27264 38058
rect 26944 37504 26952 37568
rect 27016 37504 27032 37568
rect 27096 37504 27112 37568
rect 27176 37504 27192 37568
rect 27256 37504 27264 37568
rect 26944 36480 27264 37504
rect 26944 36416 26952 36480
rect 27016 36416 27032 36480
rect 27096 36416 27112 36480
rect 27176 36416 27192 36480
rect 27256 36416 27264 36480
rect 26944 35392 27264 36416
rect 26944 35328 26952 35392
rect 27016 35328 27032 35392
rect 27096 35328 27112 35392
rect 27176 35328 27192 35392
rect 27256 35328 27264 35392
rect 26944 34304 27264 35328
rect 26944 34240 26952 34304
rect 27016 34240 27032 34304
rect 27096 34240 27112 34304
rect 27176 34240 27192 34304
rect 27256 34240 27264 34304
rect 26944 33294 27264 34240
rect 26944 33216 26986 33294
rect 27222 33216 27264 33294
rect 26944 33152 26952 33216
rect 27256 33152 27264 33216
rect 26944 33058 26986 33152
rect 27222 33058 27264 33152
rect 26944 32128 27264 33058
rect 26944 32064 26952 32128
rect 27016 32064 27032 32128
rect 27096 32064 27112 32128
rect 27176 32064 27192 32128
rect 27256 32064 27264 32128
rect 26944 31040 27264 32064
rect 26944 30976 26952 31040
rect 27016 30976 27032 31040
rect 27096 30976 27112 31040
rect 27176 30976 27192 31040
rect 27256 30976 27264 31040
rect 26944 29952 27264 30976
rect 26944 29888 26952 29952
rect 27016 29888 27032 29952
rect 27096 29888 27112 29952
rect 27176 29888 27192 29952
rect 27256 29888 27264 29952
rect 26944 28864 27264 29888
rect 26944 28800 26952 28864
rect 27016 28800 27032 28864
rect 27096 28800 27112 28864
rect 27176 28800 27192 28864
rect 27256 28800 27264 28864
rect 26944 28294 27264 28800
rect 26944 28058 26986 28294
rect 27222 28058 27264 28294
rect 26944 27776 27264 28058
rect 26944 27712 26952 27776
rect 27016 27712 27032 27776
rect 27096 27712 27112 27776
rect 27176 27712 27192 27776
rect 27256 27712 27264 27776
rect 26944 26688 27264 27712
rect 26944 26624 26952 26688
rect 27016 26624 27032 26688
rect 27096 26624 27112 26688
rect 27176 26624 27192 26688
rect 27256 26624 27264 26688
rect 26944 25600 27264 26624
rect 26944 25536 26952 25600
rect 27016 25536 27032 25600
rect 27096 25536 27112 25600
rect 27176 25536 27192 25600
rect 27256 25536 27264 25600
rect 26944 24512 27264 25536
rect 26944 24448 26952 24512
rect 27016 24448 27032 24512
rect 27096 24448 27112 24512
rect 27176 24448 27192 24512
rect 27256 24448 27264 24512
rect 26944 23424 27264 24448
rect 26944 23360 26952 23424
rect 27016 23360 27032 23424
rect 27096 23360 27112 23424
rect 27176 23360 27192 23424
rect 27256 23360 27264 23424
rect 26944 23294 27264 23360
rect 26944 23058 26986 23294
rect 27222 23058 27264 23294
rect 26944 22336 27264 23058
rect 26944 22272 26952 22336
rect 27016 22272 27032 22336
rect 27096 22272 27112 22336
rect 27176 22272 27192 22336
rect 27256 22272 27264 22336
rect 26944 21248 27264 22272
rect 26944 21184 26952 21248
rect 27016 21184 27032 21248
rect 27096 21184 27112 21248
rect 27176 21184 27192 21248
rect 27256 21184 27264 21248
rect 26944 20160 27264 21184
rect 26944 20096 26952 20160
rect 27016 20096 27032 20160
rect 27096 20096 27112 20160
rect 27176 20096 27192 20160
rect 27256 20096 27264 20160
rect 26944 19072 27264 20096
rect 26944 19008 26952 19072
rect 27016 19008 27032 19072
rect 27096 19008 27112 19072
rect 27176 19008 27192 19072
rect 27256 19008 27264 19072
rect 26944 18294 27264 19008
rect 26944 18058 26986 18294
rect 27222 18058 27264 18294
rect 26944 17984 27264 18058
rect 26944 17920 26952 17984
rect 27016 17920 27032 17984
rect 27096 17920 27112 17984
rect 27176 17920 27192 17984
rect 27256 17920 27264 17984
rect 26944 16896 27264 17920
rect 26944 16832 26952 16896
rect 27016 16832 27032 16896
rect 27096 16832 27112 16896
rect 27176 16832 27192 16896
rect 27256 16832 27264 16896
rect 26944 15808 27264 16832
rect 26944 15744 26952 15808
rect 27016 15744 27032 15808
rect 27096 15744 27112 15808
rect 27176 15744 27192 15808
rect 27256 15744 27264 15808
rect 26944 14720 27264 15744
rect 26944 14656 26952 14720
rect 27016 14656 27032 14720
rect 27096 14656 27112 14720
rect 27176 14656 27192 14720
rect 27256 14656 27264 14720
rect 26944 13632 27264 14656
rect 26944 13568 26952 13632
rect 27016 13568 27032 13632
rect 27096 13568 27112 13632
rect 27176 13568 27192 13632
rect 27256 13568 27264 13632
rect 26944 13294 27264 13568
rect 26944 13058 26986 13294
rect 27222 13058 27264 13294
rect 26944 12544 27264 13058
rect 26944 12480 26952 12544
rect 27016 12480 27032 12544
rect 27096 12480 27112 12544
rect 27176 12480 27192 12544
rect 27256 12480 27264 12544
rect 26944 11456 27264 12480
rect 26944 11392 26952 11456
rect 27016 11392 27032 11456
rect 27096 11392 27112 11456
rect 27176 11392 27192 11456
rect 27256 11392 27264 11456
rect 26944 10368 27264 11392
rect 26944 10304 26952 10368
rect 27016 10304 27032 10368
rect 27096 10304 27112 10368
rect 27176 10304 27192 10368
rect 27256 10304 27264 10368
rect 26944 9280 27264 10304
rect 26944 9216 26952 9280
rect 27016 9216 27032 9280
rect 27096 9216 27112 9280
rect 27176 9216 27192 9280
rect 27256 9216 27264 9280
rect 26944 8294 27264 9216
rect 26944 8192 26986 8294
rect 27222 8192 27264 8294
rect 26944 8128 26952 8192
rect 27256 8128 27264 8192
rect 26944 8058 26986 8128
rect 27222 8058 27264 8128
rect 26944 7104 27264 8058
rect 26944 7040 26952 7104
rect 27016 7040 27032 7104
rect 27096 7040 27112 7104
rect 27176 7040 27192 7104
rect 27256 7040 27264 7104
rect 26944 6016 27264 7040
rect 26944 5952 26952 6016
rect 27016 5952 27032 6016
rect 27096 5952 27112 6016
rect 27176 5952 27192 6016
rect 27256 5952 27264 6016
rect 26944 4928 27264 5952
rect 26944 4864 26952 4928
rect 27016 4864 27032 4928
rect 27096 4864 27112 4928
rect 27176 4864 27192 4928
rect 27256 4864 27264 4928
rect 26944 3840 27264 4864
rect 26944 3776 26952 3840
rect 27016 3776 27032 3840
rect 27096 3776 27112 3840
rect 27176 3776 27192 3840
rect 27256 3776 27264 3840
rect 26944 3294 27264 3776
rect 26944 3058 26986 3294
rect 27222 3058 27264 3294
rect 26944 2752 27264 3058
rect 26944 2688 26952 2752
rect 27016 2688 27032 2752
rect 27096 2688 27112 2752
rect 27176 2688 27192 2752
rect 27256 2688 27264 2752
rect 26944 2128 27264 2688
rect 27604 57696 27924 57712
rect 27604 57632 27612 57696
rect 27676 57632 27692 57696
rect 27756 57632 27772 57696
rect 27836 57632 27852 57696
rect 27916 57632 27924 57696
rect 27604 56608 27924 57632
rect 27604 56544 27612 56608
rect 27676 56544 27692 56608
rect 27756 56544 27772 56608
rect 27836 56544 27852 56608
rect 27916 56544 27924 56608
rect 27604 55520 27924 56544
rect 27604 55456 27612 55520
rect 27676 55456 27692 55520
rect 27756 55456 27772 55520
rect 27836 55456 27852 55520
rect 27916 55456 27924 55520
rect 27604 54432 27924 55456
rect 27604 54368 27612 54432
rect 27676 54368 27692 54432
rect 27756 54368 27772 54432
rect 27836 54368 27852 54432
rect 27916 54368 27924 54432
rect 27604 53954 27924 54368
rect 27604 53718 27646 53954
rect 27882 53718 27924 53954
rect 27604 53344 27924 53718
rect 27604 53280 27612 53344
rect 27676 53280 27692 53344
rect 27756 53280 27772 53344
rect 27836 53280 27852 53344
rect 27916 53280 27924 53344
rect 27604 52256 27924 53280
rect 27604 52192 27612 52256
rect 27676 52192 27692 52256
rect 27756 52192 27772 52256
rect 27836 52192 27852 52256
rect 27916 52192 27924 52256
rect 27604 51168 27924 52192
rect 27604 51104 27612 51168
rect 27676 51104 27692 51168
rect 27756 51104 27772 51168
rect 27836 51104 27852 51168
rect 27916 51104 27924 51168
rect 27604 50080 27924 51104
rect 27604 50016 27612 50080
rect 27676 50016 27692 50080
rect 27756 50016 27772 50080
rect 27836 50016 27852 50080
rect 27916 50016 27924 50080
rect 27604 48992 27924 50016
rect 27604 48928 27612 48992
rect 27676 48954 27692 48992
rect 27756 48954 27772 48992
rect 27836 48954 27852 48992
rect 27916 48928 27924 48992
rect 27604 48718 27646 48928
rect 27882 48718 27924 48928
rect 27604 47904 27924 48718
rect 27604 47840 27612 47904
rect 27676 47840 27692 47904
rect 27756 47840 27772 47904
rect 27836 47840 27852 47904
rect 27916 47840 27924 47904
rect 27604 46816 27924 47840
rect 27604 46752 27612 46816
rect 27676 46752 27692 46816
rect 27756 46752 27772 46816
rect 27836 46752 27852 46816
rect 27916 46752 27924 46816
rect 27604 45728 27924 46752
rect 27604 45664 27612 45728
rect 27676 45664 27692 45728
rect 27756 45664 27772 45728
rect 27836 45664 27852 45728
rect 27916 45664 27924 45728
rect 27604 44640 27924 45664
rect 27604 44576 27612 44640
rect 27676 44576 27692 44640
rect 27756 44576 27772 44640
rect 27836 44576 27852 44640
rect 27916 44576 27924 44640
rect 27604 43954 27924 44576
rect 27604 43718 27646 43954
rect 27882 43718 27924 43954
rect 27604 43552 27924 43718
rect 27604 43488 27612 43552
rect 27676 43488 27692 43552
rect 27756 43488 27772 43552
rect 27836 43488 27852 43552
rect 27916 43488 27924 43552
rect 27604 42464 27924 43488
rect 27604 42400 27612 42464
rect 27676 42400 27692 42464
rect 27756 42400 27772 42464
rect 27836 42400 27852 42464
rect 27916 42400 27924 42464
rect 27604 41376 27924 42400
rect 27604 41312 27612 41376
rect 27676 41312 27692 41376
rect 27756 41312 27772 41376
rect 27836 41312 27852 41376
rect 27916 41312 27924 41376
rect 27604 40288 27924 41312
rect 27604 40224 27612 40288
rect 27676 40224 27692 40288
rect 27756 40224 27772 40288
rect 27836 40224 27852 40288
rect 27916 40224 27924 40288
rect 27604 39200 27924 40224
rect 27604 39136 27612 39200
rect 27676 39136 27692 39200
rect 27756 39136 27772 39200
rect 27836 39136 27852 39200
rect 27916 39136 27924 39200
rect 27604 38954 27924 39136
rect 27604 38718 27646 38954
rect 27882 38718 27924 38954
rect 27604 38112 27924 38718
rect 27604 38048 27612 38112
rect 27676 38048 27692 38112
rect 27756 38048 27772 38112
rect 27836 38048 27852 38112
rect 27916 38048 27924 38112
rect 27604 37024 27924 38048
rect 27604 36960 27612 37024
rect 27676 36960 27692 37024
rect 27756 36960 27772 37024
rect 27836 36960 27852 37024
rect 27916 36960 27924 37024
rect 27604 35936 27924 36960
rect 27604 35872 27612 35936
rect 27676 35872 27692 35936
rect 27756 35872 27772 35936
rect 27836 35872 27852 35936
rect 27916 35872 27924 35936
rect 27604 34848 27924 35872
rect 27604 34784 27612 34848
rect 27676 34784 27692 34848
rect 27756 34784 27772 34848
rect 27836 34784 27852 34848
rect 27916 34784 27924 34848
rect 27604 33954 27924 34784
rect 27604 33760 27646 33954
rect 27882 33760 27924 33954
rect 27604 33696 27612 33760
rect 27676 33696 27692 33718
rect 27756 33696 27772 33718
rect 27836 33696 27852 33718
rect 27916 33696 27924 33760
rect 27604 32672 27924 33696
rect 27604 32608 27612 32672
rect 27676 32608 27692 32672
rect 27756 32608 27772 32672
rect 27836 32608 27852 32672
rect 27916 32608 27924 32672
rect 27604 31584 27924 32608
rect 27604 31520 27612 31584
rect 27676 31520 27692 31584
rect 27756 31520 27772 31584
rect 27836 31520 27852 31584
rect 27916 31520 27924 31584
rect 27604 30496 27924 31520
rect 27604 30432 27612 30496
rect 27676 30432 27692 30496
rect 27756 30432 27772 30496
rect 27836 30432 27852 30496
rect 27916 30432 27924 30496
rect 27604 29408 27924 30432
rect 27604 29344 27612 29408
rect 27676 29344 27692 29408
rect 27756 29344 27772 29408
rect 27836 29344 27852 29408
rect 27916 29344 27924 29408
rect 27604 28954 27924 29344
rect 27604 28718 27646 28954
rect 27882 28718 27924 28954
rect 27604 28320 27924 28718
rect 27604 28256 27612 28320
rect 27676 28256 27692 28320
rect 27756 28256 27772 28320
rect 27836 28256 27852 28320
rect 27916 28256 27924 28320
rect 27604 27232 27924 28256
rect 27604 27168 27612 27232
rect 27676 27168 27692 27232
rect 27756 27168 27772 27232
rect 27836 27168 27852 27232
rect 27916 27168 27924 27232
rect 27604 26144 27924 27168
rect 27604 26080 27612 26144
rect 27676 26080 27692 26144
rect 27756 26080 27772 26144
rect 27836 26080 27852 26144
rect 27916 26080 27924 26144
rect 27604 25056 27924 26080
rect 27604 24992 27612 25056
rect 27676 24992 27692 25056
rect 27756 24992 27772 25056
rect 27836 24992 27852 25056
rect 27916 24992 27924 25056
rect 27604 23968 27924 24992
rect 27604 23904 27612 23968
rect 27676 23954 27692 23968
rect 27756 23954 27772 23968
rect 27836 23954 27852 23968
rect 27916 23904 27924 23968
rect 27604 23718 27646 23904
rect 27882 23718 27924 23904
rect 27604 22880 27924 23718
rect 27604 22816 27612 22880
rect 27676 22816 27692 22880
rect 27756 22816 27772 22880
rect 27836 22816 27852 22880
rect 27916 22816 27924 22880
rect 27604 21792 27924 22816
rect 27604 21728 27612 21792
rect 27676 21728 27692 21792
rect 27756 21728 27772 21792
rect 27836 21728 27852 21792
rect 27916 21728 27924 21792
rect 27604 20704 27924 21728
rect 27604 20640 27612 20704
rect 27676 20640 27692 20704
rect 27756 20640 27772 20704
rect 27836 20640 27852 20704
rect 27916 20640 27924 20704
rect 27604 19616 27924 20640
rect 27604 19552 27612 19616
rect 27676 19552 27692 19616
rect 27756 19552 27772 19616
rect 27836 19552 27852 19616
rect 27916 19552 27924 19616
rect 27604 18954 27924 19552
rect 27604 18718 27646 18954
rect 27882 18718 27924 18954
rect 27604 18528 27924 18718
rect 27604 18464 27612 18528
rect 27676 18464 27692 18528
rect 27756 18464 27772 18528
rect 27836 18464 27852 18528
rect 27916 18464 27924 18528
rect 27604 17440 27924 18464
rect 27604 17376 27612 17440
rect 27676 17376 27692 17440
rect 27756 17376 27772 17440
rect 27836 17376 27852 17440
rect 27916 17376 27924 17440
rect 27604 16352 27924 17376
rect 27604 16288 27612 16352
rect 27676 16288 27692 16352
rect 27756 16288 27772 16352
rect 27836 16288 27852 16352
rect 27916 16288 27924 16352
rect 27604 15264 27924 16288
rect 27604 15200 27612 15264
rect 27676 15200 27692 15264
rect 27756 15200 27772 15264
rect 27836 15200 27852 15264
rect 27916 15200 27924 15264
rect 27604 14176 27924 15200
rect 27604 14112 27612 14176
rect 27676 14112 27692 14176
rect 27756 14112 27772 14176
rect 27836 14112 27852 14176
rect 27916 14112 27924 14176
rect 27604 13954 27924 14112
rect 27604 13718 27646 13954
rect 27882 13718 27924 13954
rect 27604 13088 27924 13718
rect 27604 13024 27612 13088
rect 27676 13024 27692 13088
rect 27756 13024 27772 13088
rect 27836 13024 27852 13088
rect 27916 13024 27924 13088
rect 27604 12000 27924 13024
rect 27604 11936 27612 12000
rect 27676 11936 27692 12000
rect 27756 11936 27772 12000
rect 27836 11936 27852 12000
rect 27916 11936 27924 12000
rect 27604 10912 27924 11936
rect 27604 10848 27612 10912
rect 27676 10848 27692 10912
rect 27756 10848 27772 10912
rect 27836 10848 27852 10912
rect 27916 10848 27924 10912
rect 27604 9824 27924 10848
rect 27604 9760 27612 9824
rect 27676 9760 27692 9824
rect 27756 9760 27772 9824
rect 27836 9760 27852 9824
rect 27916 9760 27924 9824
rect 27604 8954 27924 9760
rect 27604 8736 27646 8954
rect 27882 8736 27924 8954
rect 27604 8672 27612 8736
rect 27676 8672 27692 8718
rect 27756 8672 27772 8718
rect 27836 8672 27852 8718
rect 27916 8672 27924 8736
rect 27604 7648 27924 8672
rect 27604 7584 27612 7648
rect 27676 7584 27692 7648
rect 27756 7584 27772 7648
rect 27836 7584 27852 7648
rect 27916 7584 27924 7648
rect 27604 6560 27924 7584
rect 27604 6496 27612 6560
rect 27676 6496 27692 6560
rect 27756 6496 27772 6560
rect 27836 6496 27852 6560
rect 27916 6496 27924 6560
rect 27604 5472 27924 6496
rect 27604 5408 27612 5472
rect 27676 5408 27692 5472
rect 27756 5408 27772 5472
rect 27836 5408 27852 5472
rect 27916 5408 27924 5472
rect 27604 4384 27924 5408
rect 27604 4320 27612 4384
rect 27676 4320 27692 4384
rect 27756 4320 27772 4384
rect 27836 4320 27852 4384
rect 27916 4320 27924 4384
rect 27604 3954 27924 4320
rect 27604 3718 27646 3954
rect 27882 3718 27924 3954
rect 27604 3296 27924 3718
rect 27604 3232 27612 3296
rect 27676 3232 27692 3296
rect 27756 3232 27772 3296
rect 27836 3232 27852 3296
rect 27916 3232 27924 3296
rect 27604 2208 27924 3232
rect 27604 2144 27612 2208
rect 27676 2144 27692 2208
rect 27756 2144 27772 2208
rect 27836 2144 27852 2208
rect 27916 2144 27924 2208
rect 27604 2128 27924 2144
rect 31944 57152 32264 57712
rect 31944 57088 31952 57152
rect 32016 57088 32032 57152
rect 32096 57088 32112 57152
rect 32176 57088 32192 57152
rect 32256 57088 32264 57152
rect 31944 56064 32264 57088
rect 31944 56000 31952 56064
rect 32016 56000 32032 56064
rect 32096 56000 32112 56064
rect 32176 56000 32192 56064
rect 32256 56000 32264 56064
rect 31944 54976 32264 56000
rect 31944 54912 31952 54976
rect 32016 54912 32032 54976
rect 32096 54912 32112 54976
rect 32176 54912 32192 54976
rect 32256 54912 32264 54976
rect 31944 53888 32264 54912
rect 31944 53824 31952 53888
rect 32016 53824 32032 53888
rect 32096 53824 32112 53888
rect 32176 53824 32192 53888
rect 32256 53824 32264 53888
rect 31944 53294 32264 53824
rect 31944 53058 31986 53294
rect 32222 53058 32264 53294
rect 31944 52800 32264 53058
rect 31944 52736 31952 52800
rect 32016 52736 32032 52800
rect 32096 52736 32112 52800
rect 32176 52736 32192 52800
rect 32256 52736 32264 52800
rect 31944 51712 32264 52736
rect 31944 51648 31952 51712
rect 32016 51648 32032 51712
rect 32096 51648 32112 51712
rect 32176 51648 32192 51712
rect 32256 51648 32264 51712
rect 31944 50624 32264 51648
rect 31944 50560 31952 50624
rect 32016 50560 32032 50624
rect 32096 50560 32112 50624
rect 32176 50560 32192 50624
rect 32256 50560 32264 50624
rect 31944 49536 32264 50560
rect 31944 49472 31952 49536
rect 32016 49472 32032 49536
rect 32096 49472 32112 49536
rect 32176 49472 32192 49536
rect 32256 49472 32264 49536
rect 31944 48448 32264 49472
rect 31944 48384 31952 48448
rect 32016 48384 32032 48448
rect 32096 48384 32112 48448
rect 32176 48384 32192 48448
rect 32256 48384 32264 48448
rect 31944 48294 32264 48384
rect 31944 48058 31986 48294
rect 32222 48058 32264 48294
rect 31944 47360 32264 48058
rect 31944 47296 31952 47360
rect 32016 47296 32032 47360
rect 32096 47296 32112 47360
rect 32176 47296 32192 47360
rect 32256 47296 32264 47360
rect 31944 46272 32264 47296
rect 31944 46208 31952 46272
rect 32016 46208 32032 46272
rect 32096 46208 32112 46272
rect 32176 46208 32192 46272
rect 32256 46208 32264 46272
rect 31944 45184 32264 46208
rect 31944 45120 31952 45184
rect 32016 45120 32032 45184
rect 32096 45120 32112 45184
rect 32176 45120 32192 45184
rect 32256 45120 32264 45184
rect 31944 44096 32264 45120
rect 31944 44032 31952 44096
rect 32016 44032 32032 44096
rect 32096 44032 32112 44096
rect 32176 44032 32192 44096
rect 32256 44032 32264 44096
rect 31944 43294 32264 44032
rect 31944 43058 31986 43294
rect 32222 43058 32264 43294
rect 31944 43008 32264 43058
rect 31944 42944 31952 43008
rect 32016 42944 32032 43008
rect 32096 42944 32112 43008
rect 32176 42944 32192 43008
rect 32256 42944 32264 43008
rect 31944 41920 32264 42944
rect 31944 41856 31952 41920
rect 32016 41856 32032 41920
rect 32096 41856 32112 41920
rect 32176 41856 32192 41920
rect 32256 41856 32264 41920
rect 31944 40832 32264 41856
rect 31944 40768 31952 40832
rect 32016 40768 32032 40832
rect 32096 40768 32112 40832
rect 32176 40768 32192 40832
rect 32256 40768 32264 40832
rect 31944 39744 32264 40768
rect 31944 39680 31952 39744
rect 32016 39680 32032 39744
rect 32096 39680 32112 39744
rect 32176 39680 32192 39744
rect 32256 39680 32264 39744
rect 31944 38656 32264 39680
rect 31944 38592 31952 38656
rect 32016 38592 32032 38656
rect 32096 38592 32112 38656
rect 32176 38592 32192 38656
rect 32256 38592 32264 38656
rect 31944 38294 32264 38592
rect 31944 38058 31986 38294
rect 32222 38058 32264 38294
rect 31944 37568 32264 38058
rect 31944 37504 31952 37568
rect 32016 37504 32032 37568
rect 32096 37504 32112 37568
rect 32176 37504 32192 37568
rect 32256 37504 32264 37568
rect 31944 36480 32264 37504
rect 31944 36416 31952 36480
rect 32016 36416 32032 36480
rect 32096 36416 32112 36480
rect 32176 36416 32192 36480
rect 32256 36416 32264 36480
rect 31944 35392 32264 36416
rect 31944 35328 31952 35392
rect 32016 35328 32032 35392
rect 32096 35328 32112 35392
rect 32176 35328 32192 35392
rect 32256 35328 32264 35392
rect 31944 34304 32264 35328
rect 31944 34240 31952 34304
rect 32016 34240 32032 34304
rect 32096 34240 32112 34304
rect 32176 34240 32192 34304
rect 32256 34240 32264 34304
rect 31944 33294 32264 34240
rect 31944 33216 31986 33294
rect 32222 33216 32264 33294
rect 31944 33152 31952 33216
rect 32256 33152 32264 33216
rect 31944 33058 31986 33152
rect 32222 33058 32264 33152
rect 31944 32128 32264 33058
rect 31944 32064 31952 32128
rect 32016 32064 32032 32128
rect 32096 32064 32112 32128
rect 32176 32064 32192 32128
rect 32256 32064 32264 32128
rect 31944 31040 32264 32064
rect 31944 30976 31952 31040
rect 32016 30976 32032 31040
rect 32096 30976 32112 31040
rect 32176 30976 32192 31040
rect 32256 30976 32264 31040
rect 31944 29952 32264 30976
rect 31944 29888 31952 29952
rect 32016 29888 32032 29952
rect 32096 29888 32112 29952
rect 32176 29888 32192 29952
rect 32256 29888 32264 29952
rect 31944 28864 32264 29888
rect 31944 28800 31952 28864
rect 32016 28800 32032 28864
rect 32096 28800 32112 28864
rect 32176 28800 32192 28864
rect 32256 28800 32264 28864
rect 31944 28294 32264 28800
rect 31944 28058 31986 28294
rect 32222 28058 32264 28294
rect 31944 27776 32264 28058
rect 31944 27712 31952 27776
rect 32016 27712 32032 27776
rect 32096 27712 32112 27776
rect 32176 27712 32192 27776
rect 32256 27712 32264 27776
rect 31944 26688 32264 27712
rect 31944 26624 31952 26688
rect 32016 26624 32032 26688
rect 32096 26624 32112 26688
rect 32176 26624 32192 26688
rect 32256 26624 32264 26688
rect 31944 25600 32264 26624
rect 31944 25536 31952 25600
rect 32016 25536 32032 25600
rect 32096 25536 32112 25600
rect 32176 25536 32192 25600
rect 32256 25536 32264 25600
rect 31944 24512 32264 25536
rect 31944 24448 31952 24512
rect 32016 24448 32032 24512
rect 32096 24448 32112 24512
rect 32176 24448 32192 24512
rect 32256 24448 32264 24512
rect 31944 23424 32264 24448
rect 31944 23360 31952 23424
rect 32016 23360 32032 23424
rect 32096 23360 32112 23424
rect 32176 23360 32192 23424
rect 32256 23360 32264 23424
rect 31944 23294 32264 23360
rect 31944 23058 31986 23294
rect 32222 23058 32264 23294
rect 31944 22336 32264 23058
rect 31944 22272 31952 22336
rect 32016 22272 32032 22336
rect 32096 22272 32112 22336
rect 32176 22272 32192 22336
rect 32256 22272 32264 22336
rect 31944 21248 32264 22272
rect 31944 21184 31952 21248
rect 32016 21184 32032 21248
rect 32096 21184 32112 21248
rect 32176 21184 32192 21248
rect 32256 21184 32264 21248
rect 31944 20160 32264 21184
rect 31944 20096 31952 20160
rect 32016 20096 32032 20160
rect 32096 20096 32112 20160
rect 32176 20096 32192 20160
rect 32256 20096 32264 20160
rect 31944 19072 32264 20096
rect 31944 19008 31952 19072
rect 32016 19008 32032 19072
rect 32096 19008 32112 19072
rect 32176 19008 32192 19072
rect 32256 19008 32264 19072
rect 31944 18294 32264 19008
rect 31944 18058 31986 18294
rect 32222 18058 32264 18294
rect 31944 17984 32264 18058
rect 31944 17920 31952 17984
rect 32016 17920 32032 17984
rect 32096 17920 32112 17984
rect 32176 17920 32192 17984
rect 32256 17920 32264 17984
rect 31944 16896 32264 17920
rect 31944 16832 31952 16896
rect 32016 16832 32032 16896
rect 32096 16832 32112 16896
rect 32176 16832 32192 16896
rect 32256 16832 32264 16896
rect 31944 15808 32264 16832
rect 31944 15744 31952 15808
rect 32016 15744 32032 15808
rect 32096 15744 32112 15808
rect 32176 15744 32192 15808
rect 32256 15744 32264 15808
rect 31944 14720 32264 15744
rect 31944 14656 31952 14720
rect 32016 14656 32032 14720
rect 32096 14656 32112 14720
rect 32176 14656 32192 14720
rect 32256 14656 32264 14720
rect 31944 13632 32264 14656
rect 31944 13568 31952 13632
rect 32016 13568 32032 13632
rect 32096 13568 32112 13632
rect 32176 13568 32192 13632
rect 32256 13568 32264 13632
rect 31944 13294 32264 13568
rect 31944 13058 31986 13294
rect 32222 13058 32264 13294
rect 31944 12544 32264 13058
rect 31944 12480 31952 12544
rect 32016 12480 32032 12544
rect 32096 12480 32112 12544
rect 32176 12480 32192 12544
rect 32256 12480 32264 12544
rect 31944 11456 32264 12480
rect 31944 11392 31952 11456
rect 32016 11392 32032 11456
rect 32096 11392 32112 11456
rect 32176 11392 32192 11456
rect 32256 11392 32264 11456
rect 31944 10368 32264 11392
rect 31944 10304 31952 10368
rect 32016 10304 32032 10368
rect 32096 10304 32112 10368
rect 32176 10304 32192 10368
rect 32256 10304 32264 10368
rect 31944 9280 32264 10304
rect 31944 9216 31952 9280
rect 32016 9216 32032 9280
rect 32096 9216 32112 9280
rect 32176 9216 32192 9280
rect 32256 9216 32264 9280
rect 31944 8294 32264 9216
rect 31944 8192 31986 8294
rect 32222 8192 32264 8294
rect 31944 8128 31952 8192
rect 32256 8128 32264 8192
rect 31944 8058 31986 8128
rect 32222 8058 32264 8128
rect 31944 7104 32264 8058
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 3294 32264 3776
rect 31944 3058 31986 3294
rect 32222 3058 32264 3294
rect 31944 2752 32264 3058
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 2128 32264 2688
rect 32604 57696 32924 57712
rect 32604 57632 32612 57696
rect 32676 57632 32692 57696
rect 32756 57632 32772 57696
rect 32836 57632 32852 57696
rect 32916 57632 32924 57696
rect 32604 56608 32924 57632
rect 32604 56544 32612 56608
rect 32676 56544 32692 56608
rect 32756 56544 32772 56608
rect 32836 56544 32852 56608
rect 32916 56544 32924 56608
rect 32604 55520 32924 56544
rect 32604 55456 32612 55520
rect 32676 55456 32692 55520
rect 32756 55456 32772 55520
rect 32836 55456 32852 55520
rect 32916 55456 32924 55520
rect 32604 54432 32924 55456
rect 32604 54368 32612 54432
rect 32676 54368 32692 54432
rect 32756 54368 32772 54432
rect 32836 54368 32852 54432
rect 32916 54368 32924 54432
rect 32604 53954 32924 54368
rect 32604 53718 32646 53954
rect 32882 53718 32924 53954
rect 32604 53344 32924 53718
rect 32604 53280 32612 53344
rect 32676 53280 32692 53344
rect 32756 53280 32772 53344
rect 32836 53280 32852 53344
rect 32916 53280 32924 53344
rect 32604 52256 32924 53280
rect 32604 52192 32612 52256
rect 32676 52192 32692 52256
rect 32756 52192 32772 52256
rect 32836 52192 32852 52256
rect 32916 52192 32924 52256
rect 32604 51168 32924 52192
rect 32604 51104 32612 51168
rect 32676 51104 32692 51168
rect 32756 51104 32772 51168
rect 32836 51104 32852 51168
rect 32916 51104 32924 51168
rect 32604 50080 32924 51104
rect 32604 50016 32612 50080
rect 32676 50016 32692 50080
rect 32756 50016 32772 50080
rect 32836 50016 32852 50080
rect 32916 50016 32924 50080
rect 32604 48992 32924 50016
rect 32604 48928 32612 48992
rect 32676 48954 32692 48992
rect 32756 48954 32772 48992
rect 32836 48954 32852 48992
rect 32916 48928 32924 48992
rect 32604 48718 32646 48928
rect 32882 48718 32924 48928
rect 32604 47904 32924 48718
rect 32604 47840 32612 47904
rect 32676 47840 32692 47904
rect 32756 47840 32772 47904
rect 32836 47840 32852 47904
rect 32916 47840 32924 47904
rect 32604 46816 32924 47840
rect 32604 46752 32612 46816
rect 32676 46752 32692 46816
rect 32756 46752 32772 46816
rect 32836 46752 32852 46816
rect 32916 46752 32924 46816
rect 32604 45728 32924 46752
rect 32604 45664 32612 45728
rect 32676 45664 32692 45728
rect 32756 45664 32772 45728
rect 32836 45664 32852 45728
rect 32916 45664 32924 45728
rect 32604 44640 32924 45664
rect 32604 44576 32612 44640
rect 32676 44576 32692 44640
rect 32756 44576 32772 44640
rect 32836 44576 32852 44640
rect 32916 44576 32924 44640
rect 32604 43954 32924 44576
rect 32604 43718 32646 43954
rect 32882 43718 32924 43954
rect 32604 43552 32924 43718
rect 32604 43488 32612 43552
rect 32676 43488 32692 43552
rect 32756 43488 32772 43552
rect 32836 43488 32852 43552
rect 32916 43488 32924 43552
rect 32604 42464 32924 43488
rect 32604 42400 32612 42464
rect 32676 42400 32692 42464
rect 32756 42400 32772 42464
rect 32836 42400 32852 42464
rect 32916 42400 32924 42464
rect 32604 41376 32924 42400
rect 32604 41312 32612 41376
rect 32676 41312 32692 41376
rect 32756 41312 32772 41376
rect 32836 41312 32852 41376
rect 32916 41312 32924 41376
rect 32604 40288 32924 41312
rect 32604 40224 32612 40288
rect 32676 40224 32692 40288
rect 32756 40224 32772 40288
rect 32836 40224 32852 40288
rect 32916 40224 32924 40288
rect 32604 39200 32924 40224
rect 32604 39136 32612 39200
rect 32676 39136 32692 39200
rect 32756 39136 32772 39200
rect 32836 39136 32852 39200
rect 32916 39136 32924 39200
rect 32604 38954 32924 39136
rect 32604 38718 32646 38954
rect 32882 38718 32924 38954
rect 32604 38112 32924 38718
rect 32604 38048 32612 38112
rect 32676 38048 32692 38112
rect 32756 38048 32772 38112
rect 32836 38048 32852 38112
rect 32916 38048 32924 38112
rect 32604 37024 32924 38048
rect 32604 36960 32612 37024
rect 32676 36960 32692 37024
rect 32756 36960 32772 37024
rect 32836 36960 32852 37024
rect 32916 36960 32924 37024
rect 32604 35936 32924 36960
rect 32604 35872 32612 35936
rect 32676 35872 32692 35936
rect 32756 35872 32772 35936
rect 32836 35872 32852 35936
rect 32916 35872 32924 35936
rect 32604 34848 32924 35872
rect 32604 34784 32612 34848
rect 32676 34784 32692 34848
rect 32756 34784 32772 34848
rect 32836 34784 32852 34848
rect 32916 34784 32924 34848
rect 32604 33954 32924 34784
rect 32604 33760 32646 33954
rect 32882 33760 32924 33954
rect 32604 33696 32612 33760
rect 32676 33696 32692 33718
rect 32756 33696 32772 33718
rect 32836 33696 32852 33718
rect 32916 33696 32924 33760
rect 32604 32672 32924 33696
rect 32604 32608 32612 32672
rect 32676 32608 32692 32672
rect 32756 32608 32772 32672
rect 32836 32608 32852 32672
rect 32916 32608 32924 32672
rect 32604 31584 32924 32608
rect 32604 31520 32612 31584
rect 32676 31520 32692 31584
rect 32756 31520 32772 31584
rect 32836 31520 32852 31584
rect 32916 31520 32924 31584
rect 32604 30496 32924 31520
rect 32604 30432 32612 30496
rect 32676 30432 32692 30496
rect 32756 30432 32772 30496
rect 32836 30432 32852 30496
rect 32916 30432 32924 30496
rect 32604 29408 32924 30432
rect 32604 29344 32612 29408
rect 32676 29344 32692 29408
rect 32756 29344 32772 29408
rect 32836 29344 32852 29408
rect 32916 29344 32924 29408
rect 32604 28954 32924 29344
rect 32604 28718 32646 28954
rect 32882 28718 32924 28954
rect 32604 28320 32924 28718
rect 32604 28256 32612 28320
rect 32676 28256 32692 28320
rect 32756 28256 32772 28320
rect 32836 28256 32852 28320
rect 32916 28256 32924 28320
rect 32604 27232 32924 28256
rect 32604 27168 32612 27232
rect 32676 27168 32692 27232
rect 32756 27168 32772 27232
rect 32836 27168 32852 27232
rect 32916 27168 32924 27232
rect 32604 26144 32924 27168
rect 32604 26080 32612 26144
rect 32676 26080 32692 26144
rect 32756 26080 32772 26144
rect 32836 26080 32852 26144
rect 32916 26080 32924 26144
rect 32604 25056 32924 26080
rect 32604 24992 32612 25056
rect 32676 24992 32692 25056
rect 32756 24992 32772 25056
rect 32836 24992 32852 25056
rect 32916 24992 32924 25056
rect 32604 23968 32924 24992
rect 32604 23904 32612 23968
rect 32676 23954 32692 23968
rect 32756 23954 32772 23968
rect 32836 23954 32852 23968
rect 32916 23904 32924 23968
rect 32604 23718 32646 23904
rect 32882 23718 32924 23904
rect 32604 22880 32924 23718
rect 32604 22816 32612 22880
rect 32676 22816 32692 22880
rect 32756 22816 32772 22880
rect 32836 22816 32852 22880
rect 32916 22816 32924 22880
rect 32604 21792 32924 22816
rect 32604 21728 32612 21792
rect 32676 21728 32692 21792
rect 32756 21728 32772 21792
rect 32836 21728 32852 21792
rect 32916 21728 32924 21792
rect 32604 20704 32924 21728
rect 32604 20640 32612 20704
rect 32676 20640 32692 20704
rect 32756 20640 32772 20704
rect 32836 20640 32852 20704
rect 32916 20640 32924 20704
rect 32604 19616 32924 20640
rect 32604 19552 32612 19616
rect 32676 19552 32692 19616
rect 32756 19552 32772 19616
rect 32836 19552 32852 19616
rect 32916 19552 32924 19616
rect 32604 18954 32924 19552
rect 32604 18718 32646 18954
rect 32882 18718 32924 18954
rect 32604 18528 32924 18718
rect 32604 18464 32612 18528
rect 32676 18464 32692 18528
rect 32756 18464 32772 18528
rect 32836 18464 32852 18528
rect 32916 18464 32924 18528
rect 32604 17440 32924 18464
rect 32604 17376 32612 17440
rect 32676 17376 32692 17440
rect 32756 17376 32772 17440
rect 32836 17376 32852 17440
rect 32916 17376 32924 17440
rect 32604 16352 32924 17376
rect 32604 16288 32612 16352
rect 32676 16288 32692 16352
rect 32756 16288 32772 16352
rect 32836 16288 32852 16352
rect 32916 16288 32924 16352
rect 32604 15264 32924 16288
rect 32604 15200 32612 15264
rect 32676 15200 32692 15264
rect 32756 15200 32772 15264
rect 32836 15200 32852 15264
rect 32916 15200 32924 15264
rect 32604 14176 32924 15200
rect 32604 14112 32612 14176
rect 32676 14112 32692 14176
rect 32756 14112 32772 14176
rect 32836 14112 32852 14176
rect 32916 14112 32924 14176
rect 32604 13954 32924 14112
rect 32604 13718 32646 13954
rect 32882 13718 32924 13954
rect 32604 13088 32924 13718
rect 32604 13024 32612 13088
rect 32676 13024 32692 13088
rect 32756 13024 32772 13088
rect 32836 13024 32852 13088
rect 32916 13024 32924 13088
rect 32604 12000 32924 13024
rect 32604 11936 32612 12000
rect 32676 11936 32692 12000
rect 32756 11936 32772 12000
rect 32836 11936 32852 12000
rect 32916 11936 32924 12000
rect 32604 10912 32924 11936
rect 32604 10848 32612 10912
rect 32676 10848 32692 10912
rect 32756 10848 32772 10912
rect 32836 10848 32852 10912
rect 32916 10848 32924 10912
rect 32604 9824 32924 10848
rect 32604 9760 32612 9824
rect 32676 9760 32692 9824
rect 32756 9760 32772 9824
rect 32836 9760 32852 9824
rect 32916 9760 32924 9824
rect 32604 8954 32924 9760
rect 32604 8736 32646 8954
rect 32882 8736 32924 8954
rect 32604 8672 32612 8736
rect 32676 8672 32692 8718
rect 32756 8672 32772 8718
rect 32836 8672 32852 8718
rect 32916 8672 32924 8736
rect 32604 7648 32924 8672
rect 32604 7584 32612 7648
rect 32676 7584 32692 7648
rect 32756 7584 32772 7648
rect 32836 7584 32852 7648
rect 32916 7584 32924 7648
rect 32604 6560 32924 7584
rect 32604 6496 32612 6560
rect 32676 6496 32692 6560
rect 32756 6496 32772 6560
rect 32836 6496 32852 6560
rect 32916 6496 32924 6560
rect 32604 5472 32924 6496
rect 32604 5408 32612 5472
rect 32676 5408 32692 5472
rect 32756 5408 32772 5472
rect 32836 5408 32852 5472
rect 32916 5408 32924 5472
rect 32604 4384 32924 5408
rect 32604 4320 32612 4384
rect 32676 4320 32692 4384
rect 32756 4320 32772 4384
rect 32836 4320 32852 4384
rect 32916 4320 32924 4384
rect 32604 3954 32924 4320
rect 32604 3718 32646 3954
rect 32882 3718 32924 3954
rect 32604 3296 32924 3718
rect 32604 3232 32612 3296
rect 32676 3232 32692 3296
rect 32756 3232 32772 3296
rect 32836 3232 32852 3296
rect 32916 3232 32924 3296
rect 32604 2208 32924 3232
rect 32604 2144 32612 2208
rect 32676 2144 32692 2208
rect 32756 2144 32772 2208
rect 32836 2144 32852 2208
rect 32916 2144 32924 2208
rect 32604 2128 32924 2144
rect 36944 57152 37264 57712
rect 36944 57088 36952 57152
rect 37016 57088 37032 57152
rect 37096 57088 37112 57152
rect 37176 57088 37192 57152
rect 37256 57088 37264 57152
rect 36944 56064 37264 57088
rect 36944 56000 36952 56064
rect 37016 56000 37032 56064
rect 37096 56000 37112 56064
rect 37176 56000 37192 56064
rect 37256 56000 37264 56064
rect 36944 54976 37264 56000
rect 36944 54912 36952 54976
rect 37016 54912 37032 54976
rect 37096 54912 37112 54976
rect 37176 54912 37192 54976
rect 37256 54912 37264 54976
rect 36944 53888 37264 54912
rect 36944 53824 36952 53888
rect 37016 53824 37032 53888
rect 37096 53824 37112 53888
rect 37176 53824 37192 53888
rect 37256 53824 37264 53888
rect 36944 53294 37264 53824
rect 36944 53058 36986 53294
rect 37222 53058 37264 53294
rect 36944 52800 37264 53058
rect 36944 52736 36952 52800
rect 37016 52736 37032 52800
rect 37096 52736 37112 52800
rect 37176 52736 37192 52800
rect 37256 52736 37264 52800
rect 36944 51712 37264 52736
rect 36944 51648 36952 51712
rect 37016 51648 37032 51712
rect 37096 51648 37112 51712
rect 37176 51648 37192 51712
rect 37256 51648 37264 51712
rect 36944 50624 37264 51648
rect 36944 50560 36952 50624
rect 37016 50560 37032 50624
rect 37096 50560 37112 50624
rect 37176 50560 37192 50624
rect 37256 50560 37264 50624
rect 36944 49536 37264 50560
rect 36944 49472 36952 49536
rect 37016 49472 37032 49536
rect 37096 49472 37112 49536
rect 37176 49472 37192 49536
rect 37256 49472 37264 49536
rect 36944 48448 37264 49472
rect 36944 48384 36952 48448
rect 37016 48384 37032 48448
rect 37096 48384 37112 48448
rect 37176 48384 37192 48448
rect 37256 48384 37264 48448
rect 36944 48294 37264 48384
rect 36944 48058 36986 48294
rect 37222 48058 37264 48294
rect 36944 47360 37264 48058
rect 36944 47296 36952 47360
rect 37016 47296 37032 47360
rect 37096 47296 37112 47360
rect 37176 47296 37192 47360
rect 37256 47296 37264 47360
rect 36944 46272 37264 47296
rect 36944 46208 36952 46272
rect 37016 46208 37032 46272
rect 37096 46208 37112 46272
rect 37176 46208 37192 46272
rect 37256 46208 37264 46272
rect 36944 45184 37264 46208
rect 36944 45120 36952 45184
rect 37016 45120 37032 45184
rect 37096 45120 37112 45184
rect 37176 45120 37192 45184
rect 37256 45120 37264 45184
rect 36944 44096 37264 45120
rect 36944 44032 36952 44096
rect 37016 44032 37032 44096
rect 37096 44032 37112 44096
rect 37176 44032 37192 44096
rect 37256 44032 37264 44096
rect 36944 43294 37264 44032
rect 36944 43058 36986 43294
rect 37222 43058 37264 43294
rect 36944 43008 37264 43058
rect 36944 42944 36952 43008
rect 37016 42944 37032 43008
rect 37096 42944 37112 43008
rect 37176 42944 37192 43008
rect 37256 42944 37264 43008
rect 36944 41920 37264 42944
rect 36944 41856 36952 41920
rect 37016 41856 37032 41920
rect 37096 41856 37112 41920
rect 37176 41856 37192 41920
rect 37256 41856 37264 41920
rect 36944 40832 37264 41856
rect 36944 40768 36952 40832
rect 37016 40768 37032 40832
rect 37096 40768 37112 40832
rect 37176 40768 37192 40832
rect 37256 40768 37264 40832
rect 36944 39744 37264 40768
rect 36944 39680 36952 39744
rect 37016 39680 37032 39744
rect 37096 39680 37112 39744
rect 37176 39680 37192 39744
rect 37256 39680 37264 39744
rect 36944 38656 37264 39680
rect 36944 38592 36952 38656
rect 37016 38592 37032 38656
rect 37096 38592 37112 38656
rect 37176 38592 37192 38656
rect 37256 38592 37264 38656
rect 36944 38294 37264 38592
rect 36944 38058 36986 38294
rect 37222 38058 37264 38294
rect 36944 37568 37264 38058
rect 36944 37504 36952 37568
rect 37016 37504 37032 37568
rect 37096 37504 37112 37568
rect 37176 37504 37192 37568
rect 37256 37504 37264 37568
rect 36944 36480 37264 37504
rect 36944 36416 36952 36480
rect 37016 36416 37032 36480
rect 37096 36416 37112 36480
rect 37176 36416 37192 36480
rect 37256 36416 37264 36480
rect 36944 35392 37264 36416
rect 36944 35328 36952 35392
rect 37016 35328 37032 35392
rect 37096 35328 37112 35392
rect 37176 35328 37192 35392
rect 37256 35328 37264 35392
rect 36944 34304 37264 35328
rect 36944 34240 36952 34304
rect 37016 34240 37032 34304
rect 37096 34240 37112 34304
rect 37176 34240 37192 34304
rect 37256 34240 37264 34304
rect 36944 33294 37264 34240
rect 36944 33216 36986 33294
rect 37222 33216 37264 33294
rect 36944 33152 36952 33216
rect 37256 33152 37264 33216
rect 36944 33058 36986 33152
rect 37222 33058 37264 33152
rect 36944 32128 37264 33058
rect 36944 32064 36952 32128
rect 37016 32064 37032 32128
rect 37096 32064 37112 32128
rect 37176 32064 37192 32128
rect 37256 32064 37264 32128
rect 36944 31040 37264 32064
rect 36944 30976 36952 31040
rect 37016 30976 37032 31040
rect 37096 30976 37112 31040
rect 37176 30976 37192 31040
rect 37256 30976 37264 31040
rect 36944 29952 37264 30976
rect 36944 29888 36952 29952
rect 37016 29888 37032 29952
rect 37096 29888 37112 29952
rect 37176 29888 37192 29952
rect 37256 29888 37264 29952
rect 36944 28864 37264 29888
rect 36944 28800 36952 28864
rect 37016 28800 37032 28864
rect 37096 28800 37112 28864
rect 37176 28800 37192 28864
rect 37256 28800 37264 28864
rect 36944 28294 37264 28800
rect 36944 28058 36986 28294
rect 37222 28058 37264 28294
rect 36944 27776 37264 28058
rect 36944 27712 36952 27776
rect 37016 27712 37032 27776
rect 37096 27712 37112 27776
rect 37176 27712 37192 27776
rect 37256 27712 37264 27776
rect 36944 26688 37264 27712
rect 36944 26624 36952 26688
rect 37016 26624 37032 26688
rect 37096 26624 37112 26688
rect 37176 26624 37192 26688
rect 37256 26624 37264 26688
rect 36944 25600 37264 26624
rect 36944 25536 36952 25600
rect 37016 25536 37032 25600
rect 37096 25536 37112 25600
rect 37176 25536 37192 25600
rect 37256 25536 37264 25600
rect 36944 24512 37264 25536
rect 36944 24448 36952 24512
rect 37016 24448 37032 24512
rect 37096 24448 37112 24512
rect 37176 24448 37192 24512
rect 37256 24448 37264 24512
rect 36944 23424 37264 24448
rect 36944 23360 36952 23424
rect 37016 23360 37032 23424
rect 37096 23360 37112 23424
rect 37176 23360 37192 23424
rect 37256 23360 37264 23424
rect 36944 23294 37264 23360
rect 36944 23058 36986 23294
rect 37222 23058 37264 23294
rect 36944 22336 37264 23058
rect 36944 22272 36952 22336
rect 37016 22272 37032 22336
rect 37096 22272 37112 22336
rect 37176 22272 37192 22336
rect 37256 22272 37264 22336
rect 36944 21248 37264 22272
rect 36944 21184 36952 21248
rect 37016 21184 37032 21248
rect 37096 21184 37112 21248
rect 37176 21184 37192 21248
rect 37256 21184 37264 21248
rect 36944 20160 37264 21184
rect 36944 20096 36952 20160
rect 37016 20096 37032 20160
rect 37096 20096 37112 20160
rect 37176 20096 37192 20160
rect 37256 20096 37264 20160
rect 36944 19072 37264 20096
rect 36944 19008 36952 19072
rect 37016 19008 37032 19072
rect 37096 19008 37112 19072
rect 37176 19008 37192 19072
rect 37256 19008 37264 19072
rect 36944 18294 37264 19008
rect 36944 18058 36986 18294
rect 37222 18058 37264 18294
rect 36944 17984 37264 18058
rect 36944 17920 36952 17984
rect 37016 17920 37032 17984
rect 37096 17920 37112 17984
rect 37176 17920 37192 17984
rect 37256 17920 37264 17984
rect 36944 16896 37264 17920
rect 36944 16832 36952 16896
rect 37016 16832 37032 16896
rect 37096 16832 37112 16896
rect 37176 16832 37192 16896
rect 37256 16832 37264 16896
rect 36944 15808 37264 16832
rect 36944 15744 36952 15808
rect 37016 15744 37032 15808
rect 37096 15744 37112 15808
rect 37176 15744 37192 15808
rect 37256 15744 37264 15808
rect 36944 14720 37264 15744
rect 36944 14656 36952 14720
rect 37016 14656 37032 14720
rect 37096 14656 37112 14720
rect 37176 14656 37192 14720
rect 37256 14656 37264 14720
rect 36944 13632 37264 14656
rect 36944 13568 36952 13632
rect 37016 13568 37032 13632
rect 37096 13568 37112 13632
rect 37176 13568 37192 13632
rect 37256 13568 37264 13632
rect 36944 13294 37264 13568
rect 36944 13058 36986 13294
rect 37222 13058 37264 13294
rect 36944 12544 37264 13058
rect 36944 12480 36952 12544
rect 37016 12480 37032 12544
rect 37096 12480 37112 12544
rect 37176 12480 37192 12544
rect 37256 12480 37264 12544
rect 36944 11456 37264 12480
rect 36944 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37264 11456
rect 36944 10368 37264 11392
rect 36944 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37264 10368
rect 36944 9280 37264 10304
rect 36944 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37264 9280
rect 36944 8294 37264 9216
rect 36944 8192 36986 8294
rect 37222 8192 37264 8294
rect 36944 8128 36952 8192
rect 37256 8128 37264 8192
rect 36944 8058 36986 8128
rect 37222 8058 37264 8128
rect 36944 7104 37264 8058
rect 36944 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37264 7104
rect 36944 6016 37264 7040
rect 36944 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37264 6016
rect 36944 4928 37264 5952
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 3840 37264 4864
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 3294 37264 3776
rect 36944 3058 36986 3294
rect 37222 3058 37264 3294
rect 36944 2752 37264 3058
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 2128 37264 2688
rect 37604 57696 37924 57712
rect 37604 57632 37612 57696
rect 37676 57632 37692 57696
rect 37756 57632 37772 57696
rect 37836 57632 37852 57696
rect 37916 57632 37924 57696
rect 37604 56608 37924 57632
rect 37604 56544 37612 56608
rect 37676 56544 37692 56608
rect 37756 56544 37772 56608
rect 37836 56544 37852 56608
rect 37916 56544 37924 56608
rect 37604 55520 37924 56544
rect 37604 55456 37612 55520
rect 37676 55456 37692 55520
rect 37756 55456 37772 55520
rect 37836 55456 37852 55520
rect 37916 55456 37924 55520
rect 37604 54432 37924 55456
rect 37604 54368 37612 54432
rect 37676 54368 37692 54432
rect 37756 54368 37772 54432
rect 37836 54368 37852 54432
rect 37916 54368 37924 54432
rect 37604 53954 37924 54368
rect 37604 53718 37646 53954
rect 37882 53718 37924 53954
rect 37604 53344 37924 53718
rect 37604 53280 37612 53344
rect 37676 53280 37692 53344
rect 37756 53280 37772 53344
rect 37836 53280 37852 53344
rect 37916 53280 37924 53344
rect 37604 52256 37924 53280
rect 37604 52192 37612 52256
rect 37676 52192 37692 52256
rect 37756 52192 37772 52256
rect 37836 52192 37852 52256
rect 37916 52192 37924 52256
rect 37604 51168 37924 52192
rect 37604 51104 37612 51168
rect 37676 51104 37692 51168
rect 37756 51104 37772 51168
rect 37836 51104 37852 51168
rect 37916 51104 37924 51168
rect 37604 50080 37924 51104
rect 37604 50016 37612 50080
rect 37676 50016 37692 50080
rect 37756 50016 37772 50080
rect 37836 50016 37852 50080
rect 37916 50016 37924 50080
rect 37604 48992 37924 50016
rect 37604 48928 37612 48992
rect 37676 48954 37692 48992
rect 37756 48954 37772 48992
rect 37836 48954 37852 48992
rect 37916 48928 37924 48992
rect 37604 48718 37646 48928
rect 37882 48718 37924 48928
rect 37604 47904 37924 48718
rect 37604 47840 37612 47904
rect 37676 47840 37692 47904
rect 37756 47840 37772 47904
rect 37836 47840 37852 47904
rect 37916 47840 37924 47904
rect 37604 46816 37924 47840
rect 37604 46752 37612 46816
rect 37676 46752 37692 46816
rect 37756 46752 37772 46816
rect 37836 46752 37852 46816
rect 37916 46752 37924 46816
rect 37604 45728 37924 46752
rect 37604 45664 37612 45728
rect 37676 45664 37692 45728
rect 37756 45664 37772 45728
rect 37836 45664 37852 45728
rect 37916 45664 37924 45728
rect 37604 44640 37924 45664
rect 37604 44576 37612 44640
rect 37676 44576 37692 44640
rect 37756 44576 37772 44640
rect 37836 44576 37852 44640
rect 37916 44576 37924 44640
rect 37604 43954 37924 44576
rect 37604 43718 37646 43954
rect 37882 43718 37924 43954
rect 37604 43552 37924 43718
rect 37604 43488 37612 43552
rect 37676 43488 37692 43552
rect 37756 43488 37772 43552
rect 37836 43488 37852 43552
rect 37916 43488 37924 43552
rect 37604 42464 37924 43488
rect 37604 42400 37612 42464
rect 37676 42400 37692 42464
rect 37756 42400 37772 42464
rect 37836 42400 37852 42464
rect 37916 42400 37924 42464
rect 37604 41376 37924 42400
rect 37604 41312 37612 41376
rect 37676 41312 37692 41376
rect 37756 41312 37772 41376
rect 37836 41312 37852 41376
rect 37916 41312 37924 41376
rect 37604 40288 37924 41312
rect 37604 40224 37612 40288
rect 37676 40224 37692 40288
rect 37756 40224 37772 40288
rect 37836 40224 37852 40288
rect 37916 40224 37924 40288
rect 37604 39200 37924 40224
rect 37604 39136 37612 39200
rect 37676 39136 37692 39200
rect 37756 39136 37772 39200
rect 37836 39136 37852 39200
rect 37916 39136 37924 39200
rect 37604 38954 37924 39136
rect 37604 38718 37646 38954
rect 37882 38718 37924 38954
rect 37604 38112 37924 38718
rect 37604 38048 37612 38112
rect 37676 38048 37692 38112
rect 37756 38048 37772 38112
rect 37836 38048 37852 38112
rect 37916 38048 37924 38112
rect 37604 37024 37924 38048
rect 37604 36960 37612 37024
rect 37676 36960 37692 37024
rect 37756 36960 37772 37024
rect 37836 36960 37852 37024
rect 37916 36960 37924 37024
rect 37604 35936 37924 36960
rect 37604 35872 37612 35936
rect 37676 35872 37692 35936
rect 37756 35872 37772 35936
rect 37836 35872 37852 35936
rect 37916 35872 37924 35936
rect 37604 34848 37924 35872
rect 37604 34784 37612 34848
rect 37676 34784 37692 34848
rect 37756 34784 37772 34848
rect 37836 34784 37852 34848
rect 37916 34784 37924 34848
rect 37604 33954 37924 34784
rect 37604 33760 37646 33954
rect 37882 33760 37924 33954
rect 37604 33696 37612 33760
rect 37676 33696 37692 33718
rect 37756 33696 37772 33718
rect 37836 33696 37852 33718
rect 37916 33696 37924 33760
rect 37604 32672 37924 33696
rect 37604 32608 37612 32672
rect 37676 32608 37692 32672
rect 37756 32608 37772 32672
rect 37836 32608 37852 32672
rect 37916 32608 37924 32672
rect 37604 31584 37924 32608
rect 37604 31520 37612 31584
rect 37676 31520 37692 31584
rect 37756 31520 37772 31584
rect 37836 31520 37852 31584
rect 37916 31520 37924 31584
rect 37604 30496 37924 31520
rect 37604 30432 37612 30496
rect 37676 30432 37692 30496
rect 37756 30432 37772 30496
rect 37836 30432 37852 30496
rect 37916 30432 37924 30496
rect 37604 29408 37924 30432
rect 37604 29344 37612 29408
rect 37676 29344 37692 29408
rect 37756 29344 37772 29408
rect 37836 29344 37852 29408
rect 37916 29344 37924 29408
rect 37604 28954 37924 29344
rect 37604 28718 37646 28954
rect 37882 28718 37924 28954
rect 37604 28320 37924 28718
rect 37604 28256 37612 28320
rect 37676 28256 37692 28320
rect 37756 28256 37772 28320
rect 37836 28256 37852 28320
rect 37916 28256 37924 28320
rect 37604 27232 37924 28256
rect 37604 27168 37612 27232
rect 37676 27168 37692 27232
rect 37756 27168 37772 27232
rect 37836 27168 37852 27232
rect 37916 27168 37924 27232
rect 37604 26144 37924 27168
rect 37604 26080 37612 26144
rect 37676 26080 37692 26144
rect 37756 26080 37772 26144
rect 37836 26080 37852 26144
rect 37916 26080 37924 26144
rect 37604 25056 37924 26080
rect 37604 24992 37612 25056
rect 37676 24992 37692 25056
rect 37756 24992 37772 25056
rect 37836 24992 37852 25056
rect 37916 24992 37924 25056
rect 37604 23968 37924 24992
rect 37604 23904 37612 23968
rect 37676 23954 37692 23968
rect 37756 23954 37772 23968
rect 37836 23954 37852 23968
rect 37916 23904 37924 23968
rect 37604 23718 37646 23904
rect 37882 23718 37924 23904
rect 37604 22880 37924 23718
rect 37604 22816 37612 22880
rect 37676 22816 37692 22880
rect 37756 22816 37772 22880
rect 37836 22816 37852 22880
rect 37916 22816 37924 22880
rect 37604 21792 37924 22816
rect 37604 21728 37612 21792
rect 37676 21728 37692 21792
rect 37756 21728 37772 21792
rect 37836 21728 37852 21792
rect 37916 21728 37924 21792
rect 37604 20704 37924 21728
rect 37604 20640 37612 20704
rect 37676 20640 37692 20704
rect 37756 20640 37772 20704
rect 37836 20640 37852 20704
rect 37916 20640 37924 20704
rect 37604 19616 37924 20640
rect 37604 19552 37612 19616
rect 37676 19552 37692 19616
rect 37756 19552 37772 19616
rect 37836 19552 37852 19616
rect 37916 19552 37924 19616
rect 37604 18954 37924 19552
rect 37604 18718 37646 18954
rect 37882 18718 37924 18954
rect 37604 18528 37924 18718
rect 37604 18464 37612 18528
rect 37676 18464 37692 18528
rect 37756 18464 37772 18528
rect 37836 18464 37852 18528
rect 37916 18464 37924 18528
rect 37604 17440 37924 18464
rect 37604 17376 37612 17440
rect 37676 17376 37692 17440
rect 37756 17376 37772 17440
rect 37836 17376 37852 17440
rect 37916 17376 37924 17440
rect 37604 16352 37924 17376
rect 37604 16288 37612 16352
rect 37676 16288 37692 16352
rect 37756 16288 37772 16352
rect 37836 16288 37852 16352
rect 37916 16288 37924 16352
rect 37604 15264 37924 16288
rect 37604 15200 37612 15264
rect 37676 15200 37692 15264
rect 37756 15200 37772 15264
rect 37836 15200 37852 15264
rect 37916 15200 37924 15264
rect 37604 14176 37924 15200
rect 37604 14112 37612 14176
rect 37676 14112 37692 14176
rect 37756 14112 37772 14176
rect 37836 14112 37852 14176
rect 37916 14112 37924 14176
rect 37604 13954 37924 14112
rect 37604 13718 37646 13954
rect 37882 13718 37924 13954
rect 37604 13088 37924 13718
rect 37604 13024 37612 13088
rect 37676 13024 37692 13088
rect 37756 13024 37772 13088
rect 37836 13024 37852 13088
rect 37916 13024 37924 13088
rect 37604 12000 37924 13024
rect 37604 11936 37612 12000
rect 37676 11936 37692 12000
rect 37756 11936 37772 12000
rect 37836 11936 37852 12000
rect 37916 11936 37924 12000
rect 37604 10912 37924 11936
rect 37604 10848 37612 10912
rect 37676 10848 37692 10912
rect 37756 10848 37772 10912
rect 37836 10848 37852 10912
rect 37916 10848 37924 10912
rect 37604 9824 37924 10848
rect 37604 9760 37612 9824
rect 37676 9760 37692 9824
rect 37756 9760 37772 9824
rect 37836 9760 37852 9824
rect 37916 9760 37924 9824
rect 37604 8954 37924 9760
rect 37604 8736 37646 8954
rect 37882 8736 37924 8954
rect 37604 8672 37612 8736
rect 37676 8672 37692 8718
rect 37756 8672 37772 8718
rect 37836 8672 37852 8718
rect 37916 8672 37924 8736
rect 37604 7648 37924 8672
rect 37604 7584 37612 7648
rect 37676 7584 37692 7648
rect 37756 7584 37772 7648
rect 37836 7584 37852 7648
rect 37916 7584 37924 7648
rect 37604 6560 37924 7584
rect 37604 6496 37612 6560
rect 37676 6496 37692 6560
rect 37756 6496 37772 6560
rect 37836 6496 37852 6560
rect 37916 6496 37924 6560
rect 37604 5472 37924 6496
rect 37604 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37924 5472
rect 37604 4384 37924 5408
rect 37604 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37924 4384
rect 37604 3954 37924 4320
rect 37604 3718 37646 3954
rect 37882 3718 37924 3954
rect 37604 3296 37924 3718
rect 37604 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37924 3296
rect 37604 2208 37924 3232
rect 37604 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37924 2208
rect 37604 2128 37924 2144
rect 41944 57152 42264 57712
rect 41944 57088 41952 57152
rect 42016 57088 42032 57152
rect 42096 57088 42112 57152
rect 42176 57088 42192 57152
rect 42256 57088 42264 57152
rect 41944 56064 42264 57088
rect 41944 56000 41952 56064
rect 42016 56000 42032 56064
rect 42096 56000 42112 56064
rect 42176 56000 42192 56064
rect 42256 56000 42264 56064
rect 41944 54976 42264 56000
rect 41944 54912 41952 54976
rect 42016 54912 42032 54976
rect 42096 54912 42112 54976
rect 42176 54912 42192 54976
rect 42256 54912 42264 54976
rect 41944 53888 42264 54912
rect 41944 53824 41952 53888
rect 42016 53824 42032 53888
rect 42096 53824 42112 53888
rect 42176 53824 42192 53888
rect 42256 53824 42264 53888
rect 41944 53294 42264 53824
rect 41944 53058 41986 53294
rect 42222 53058 42264 53294
rect 41944 52800 42264 53058
rect 41944 52736 41952 52800
rect 42016 52736 42032 52800
rect 42096 52736 42112 52800
rect 42176 52736 42192 52800
rect 42256 52736 42264 52800
rect 41944 51712 42264 52736
rect 41944 51648 41952 51712
rect 42016 51648 42032 51712
rect 42096 51648 42112 51712
rect 42176 51648 42192 51712
rect 42256 51648 42264 51712
rect 41944 50624 42264 51648
rect 41944 50560 41952 50624
rect 42016 50560 42032 50624
rect 42096 50560 42112 50624
rect 42176 50560 42192 50624
rect 42256 50560 42264 50624
rect 41944 49536 42264 50560
rect 41944 49472 41952 49536
rect 42016 49472 42032 49536
rect 42096 49472 42112 49536
rect 42176 49472 42192 49536
rect 42256 49472 42264 49536
rect 41944 48448 42264 49472
rect 41944 48384 41952 48448
rect 42016 48384 42032 48448
rect 42096 48384 42112 48448
rect 42176 48384 42192 48448
rect 42256 48384 42264 48448
rect 41944 48294 42264 48384
rect 41944 48058 41986 48294
rect 42222 48058 42264 48294
rect 41944 47360 42264 48058
rect 41944 47296 41952 47360
rect 42016 47296 42032 47360
rect 42096 47296 42112 47360
rect 42176 47296 42192 47360
rect 42256 47296 42264 47360
rect 41944 46272 42264 47296
rect 41944 46208 41952 46272
rect 42016 46208 42032 46272
rect 42096 46208 42112 46272
rect 42176 46208 42192 46272
rect 42256 46208 42264 46272
rect 41944 45184 42264 46208
rect 41944 45120 41952 45184
rect 42016 45120 42032 45184
rect 42096 45120 42112 45184
rect 42176 45120 42192 45184
rect 42256 45120 42264 45184
rect 41944 44096 42264 45120
rect 41944 44032 41952 44096
rect 42016 44032 42032 44096
rect 42096 44032 42112 44096
rect 42176 44032 42192 44096
rect 42256 44032 42264 44096
rect 41944 43294 42264 44032
rect 41944 43058 41986 43294
rect 42222 43058 42264 43294
rect 41944 43008 42264 43058
rect 41944 42944 41952 43008
rect 42016 42944 42032 43008
rect 42096 42944 42112 43008
rect 42176 42944 42192 43008
rect 42256 42944 42264 43008
rect 41944 41920 42264 42944
rect 41944 41856 41952 41920
rect 42016 41856 42032 41920
rect 42096 41856 42112 41920
rect 42176 41856 42192 41920
rect 42256 41856 42264 41920
rect 41944 40832 42264 41856
rect 41944 40768 41952 40832
rect 42016 40768 42032 40832
rect 42096 40768 42112 40832
rect 42176 40768 42192 40832
rect 42256 40768 42264 40832
rect 41944 39744 42264 40768
rect 41944 39680 41952 39744
rect 42016 39680 42032 39744
rect 42096 39680 42112 39744
rect 42176 39680 42192 39744
rect 42256 39680 42264 39744
rect 41944 38656 42264 39680
rect 41944 38592 41952 38656
rect 42016 38592 42032 38656
rect 42096 38592 42112 38656
rect 42176 38592 42192 38656
rect 42256 38592 42264 38656
rect 41944 38294 42264 38592
rect 41944 38058 41986 38294
rect 42222 38058 42264 38294
rect 41944 37568 42264 38058
rect 41944 37504 41952 37568
rect 42016 37504 42032 37568
rect 42096 37504 42112 37568
rect 42176 37504 42192 37568
rect 42256 37504 42264 37568
rect 41944 36480 42264 37504
rect 41944 36416 41952 36480
rect 42016 36416 42032 36480
rect 42096 36416 42112 36480
rect 42176 36416 42192 36480
rect 42256 36416 42264 36480
rect 41944 35392 42264 36416
rect 41944 35328 41952 35392
rect 42016 35328 42032 35392
rect 42096 35328 42112 35392
rect 42176 35328 42192 35392
rect 42256 35328 42264 35392
rect 41944 34304 42264 35328
rect 41944 34240 41952 34304
rect 42016 34240 42032 34304
rect 42096 34240 42112 34304
rect 42176 34240 42192 34304
rect 42256 34240 42264 34304
rect 41944 33294 42264 34240
rect 41944 33216 41986 33294
rect 42222 33216 42264 33294
rect 41944 33152 41952 33216
rect 42256 33152 42264 33216
rect 41944 33058 41986 33152
rect 42222 33058 42264 33152
rect 41944 32128 42264 33058
rect 41944 32064 41952 32128
rect 42016 32064 42032 32128
rect 42096 32064 42112 32128
rect 42176 32064 42192 32128
rect 42256 32064 42264 32128
rect 41944 31040 42264 32064
rect 41944 30976 41952 31040
rect 42016 30976 42032 31040
rect 42096 30976 42112 31040
rect 42176 30976 42192 31040
rect 42256 30976 42264 31040
rect 41944 29952 42264 30976
rect 41944 29888 41952 29952
rect 42016 29888 42032 29952
rect 42096 29888 42112 29952
rect 42176 29888 42192 29952
rect 42256 29888 42264 29952
rect 41944 28864 42264 29888
rect 41944 28800 41952 28864
rect 42016 28800 42032 28864
rect 42096 28800 42112 28864
rect 42176 28800 42192 28864
rect 42256 28800 42264 28864
rect 41944 28294 42264 28800
rect 41944 28058 41986 28294
rect 42222 28058 42264 28294
rect 41944 27776 42264 28058
rect 41944 27712 41952 27776
rect 42016 27712 42032 27776
rect 42096 27712 42112 27776
rect 42176 27712 42192 27776
rect 42256 27712 42264 27776
rect 41944 26688 42264 27712
rect 41944 26624 41952 26688
rect 42016 26624 42032 26688
rect 42096 26624 42112 26688
rect 42176 26624 42192 26688
rect 42256 26624 42264 26688
rect 41944 25600 42264 26624
rect 41944 25536 41952 25600
rect 42016 25536 42032 25600
rect 42096 25536 42112 25600
rect 42176 25536 42192 25600
rect 42256 25536 42264 25600
rect 41944 24512 42264 25536
rect 41944 24448 41952 24512
rect 42016 24448 42032 24512
rect 42096 24448 42112 24512
rect 42176 24448 42192 24512
rect 42256 24448 42264 24512
rect 41944 23424 42264 24448
rect 41944 23360 41952 23424
rect 42016 23360 42032 23424
rect 42096 23360 42112 23424
rect 42176 23360 42192 23424
rect 42256 23360 42264 23424
rect 41944 23294 42264 23360
rect 41944 23058 41986 23294
rect 42222 23058 42264 23294
rect 41944 22336 42264 23058
rect 41944 22272 41952 22336
rect 42016 22272 42032 22336
rect 42096 22272 42112 22336
rect 42176 22272 42192 22336
rect 42256 22272 42264 22336
rect 41944 21248 42264 22272
rect 41944 21184 41952 21248
rect 42016 21184 42032 21248
rect 42096 21184 42112 21248
rect 42176 21184 42192 21248
rect 42256 21184 42264 21248
rect 41944 20160 42264 21184
rect 41944 20096 41952 20160
rect 42016 20096 42032 20160
rect 42096 20096 42112 20160
rect 42176 20096 42192 20160
rect 42256 20096 42264 20160
rect 41944 19072 42264 20096
rect 41944 19008 41952 19072
rect 42016 19008 42032 19072
rect 42096 19008 42112 19072
rect 42176 19008 42192 19072
rect 42256 19008 42264 19072
rect 41944 18294 42264 19008
rect 41944 18058 41986 18294
rect 42222 18058 42264 18294
rect 41944 17984 42264 18058
rect 41944 17920 41952 17984
rect 42016 17920 42032 17984
rect 42096 17920 42112 17984
rect 42176 17920 42192 17984
rect 42256 17920 42264 17984
rect 41944 16896 42264 17920
rect 41944 16832 41952 16896
rect 42016 16832 42032 16896
rect 42096 16832 42112 16896
rect 42176 16832 42192 16896
rect 42256 16832 42264 16896
rect 41944 15808 42264 16832
rect 41944 15744 41952 15808
rect 42016 15744 42032 15808
rect 42096 15744 42112 15808
rect 42176 15744 42192 15808
rect 42256 15744 42264 15808
rect 41944 14720 42264 15744
rect 41944 14656 41952 14720
rect 42016 14656 42032 14720
rect 42096 14656 42112 14720
rect 42176 14656 42192 14720
rect 42256 14656 42264 14720
rect 41944 13632 42264 14656
rect 41944 13568 41952 13632
rect 42016 13568 42032 13632
rect 42096 13568 42112 13632
rect 42176 13568 42192 13632
rect 42256 13568 42264 13632
rect 41944 13294 42264 13568
rect 41944 13058 41986 13294
rect 42222 13058 42264 13294
rect 41944 12544 42264 13058
rect 41944 12480 41952 12544
rect 42016 12480 42032 12544
rect 42096 12480 42112 12544
rect 42176 12480 42192 12544
rect 42256 12480 42264 12544
rect 41944 11456 42264 12480
rect 41944 11392 41952 11456
rect 42016 11392 42032 11456
rect 42096 11392 42112 11456
rect 42176 11392 42192 11456
rect 42256 11392 42264 11456
rect 41944 10368 42264 11392
rect 41944 10304 41952 10368
rect 42016 10304 42032 10368
rect 42096 10304 42112 10368
rect 42176 10304 42192 10368
rect 42256 10304 42264 10368
rect 41944 9280 42264 10304
rect 41944 9216 41952 9280
rect 42016 9216 42032 9280
rect 42096 9216 42112 9280
rect 42176 9216 42192 9280
rect 42256 9216 42264 9280
rect 41944 8294 42264 9216
rect 41944 8192 41986 8294
rect 42222 8192 42264 8294
rect 41944 8128 41952 8192
rect 42256 8128 42264 8192
rect 41944 8058 41986 8128
rect 42222 8058 42264 8128
rect 41944 7104 42264 8058
rect 41944 7040 41952 7104
rect 42016 7040 42032 7104
rect 42096 7040 42112 7104
rect 42176 7040 42192 7104
rect 42256 7040 42264 7104
rect 41944 6016 42264 7040
rect 41944 5952 41952 6016
rect 42016 5952 42032 6016
rect 42096 5952 42112 6016
rect 42176 5952 42192 6016
rect 42256 5952 42264 6016
rect 41944 4928 42264 5952
rect 41944 4864 41952 4928
rect 42016 4864 42032 4928
rect 42096 4864 42112 4928
rect 42176 4864 42192 4928
rect 42256 4864 42264 4928
rect 41944 3840 42264 4864
rect 41944 3776 41952 3840
rect 42016 3776 42032 3840
rect 42096 3776 42112 3840
rect 42176 3776 42192 3840
rect 42256 3776 42264 3840
rect 41944 3294 42264 3776
rect 41944 3058 41986 3294
rect 42222 3058 42264 3294
rect 41944 2752 42264 3058
rect 41944 2688 41952 2752
rect 42016 2688 42032 2752
rect 42096 2688 42112 2752
rect 42176 2688 42192 2752
rect 42256 2688 42264 2752
rect 41944 2128 42264 2688
rect 42604 57696 42924 57712
rect 42604 57632 42612 57696
rect 42676 57632 42692 57696
rect 42756 57632 42772 57696
rect 42836 57632 42852 57696
rect 42916 57632 42924 57696
rect 42604 56608 42924 57632
rect 42604 56544 42612 56608
rect 42676 56544 42692 56608
rect 42756 56544 42772 56608
rect 42836 56544 42852 56608
rect 42916 56544 42924 56608
rect 42604 55520 42924 56544
rect 42604 55456 42612 55520
rect 42676 55456 42692 55520
rect 42756 55456 42772 55520
rect 42836 55456 42852 55520
rect 42916 55456 42924 55520
rect 42604 54432 42924 55456
rect 42604 54368 42612 54432
rect 42676 54368 42692 54432
rect 42756 54368 42772 54432
rect 42836 54368 42852 54432
rect 42916 54368 42924 54432
rect 42604 53954 42924 54368
rect 42604 53718 42646 53954
rect 42882 53718 42924 53954
rect 42604 53344 42924 53718
rect 42604 53280 42612 53344
rect 42676 53280 42692 53344
rect 42756 53280 42772 53344
rect 42836 53280 42852 53344
rect 42916 53280 42924 53344
rect 42604 52256 42924 53280
rect 42604 52192 42612 52256
rect 42676 52192 42692 52256
rect 42756 52192 42772 52256
rect 42836 52192 42852 52256
rect 42916 52192 42924 52256
rect 42604 51168 42924 52192
rect 42604 51104 42612 51168
rect 42676 51104 42692 51168
rect 42756 51104 42772 51168
rect 42836 51104 42852 51168
rect 42916 51104 42924 51168
rect 42604 50080 42924 51104
rect 42604 50016 42612 50080
rect 42676 50016 42692 50080
rect 42756 50016 42772 50080
rect 42836 50016 42852 50080
rect 42916 50016 42924 50080
rect 42604 48992 42924 50016
rect 42604 48928 42612 48992
rect 42676 48954 42692 48992
rect 42756 48954 42772 48992
rect 42836 48954 42852 48992
rect 42916 48928 42924 48992
rect 42604 48718 42646 48928
rect 42882 48718 42924 48928
rect 42604 47904 42924 48718
rect 42604 47840 42612 47904
rect 42676 47840 42692 47904
rect 42756 47840 42772 47904
rect 42836 47840 42852 47904
rect 42916 47840 42924 47904
rect 42604 46816 42924 47840
rect 42604 46752 42612 46816
rect 42676 46752 42692 46816
rect 42756 46752 42772 46816
rect 42836 46752 42852 46816
rect 42916 46752 42924 46816
rect 42604 45728 42924 46752
rect 42604 45664 42612 45728
rect 42676 45664 42692 45728
rect 42756 45664 42772 45728
rect 42836 45664 42852 45728
rect 42916 45664 42924 45728
rect 42604 44640 42924 45664
rect 42604 44576 42612 44640
rect 42676 44576 42692 44640
rect 42756 44576 42772 44640
rect 42836 44576 42852 44640
rect 42916 44576 42924 44640
rect 42604 43954 42924 44576
rect 42604 43718 42646 43954
rect 42882 43718 42924 43954
rect 42604 43552 42924 43718
rect 42604 43488 42612 43552
rect 42676 43488 42692 43552
rect 42756 43488 42772 43552
rect 42836 43488 42852 43552
rect 42916 43488 42924 43552
rect 42604 42464 42924 43488
rect 42604 42400 42612 42464
rect 42676 42400 42692 42464
rect 42756 42400 42772 42464
rect 42836 42400 42852 42464
rect 42916 42400 42924 42464
rect 42604 41376 42924 42400
rect 42604 41312 42612 41376
rect 42676 41312 42692 41376
rect 42756 41312 42772 41376
rect 42836 41312 42852 41376
rect 42916 41312 42924 41376
rect 42604 40288 42924 41312
rect 42604 40224 42612 40288
rect 42676 40224 42692 40288
rect 42756 40224 42772 40288
rect 42836 40224 42852 40288
rect 42916 40224 42924 40288
rect 42604 39200 42924 40224
rect 42604 39136 42612 39200
rect 42676 39136 42692 39200
rect 42756 39136 42772 39200
rect 42836 39136 42852 39200
rect 42916 39136 42924 39200
rect 42604 38954 42924 39136
rect 42604 38718 42646 38954
rect 42882 38718 42924 38954
rect 42604 38112 42924 38718
rect 42604 38048 42612 38112
rect 42676 38048 42692 38112
rect 42756 38048 42772 38112
rect 42836 38048 42852 38112
rect 42916 38048 42924 38112
rect 42604 37024 42924 38048
rect 42604 36960 42612 37024
rect 42676 36960 42692 37024
rect 42756 36960 42772 37024
rect 42836 36960 42852 37024
rect 42916 36960 42924 37024
rect 42604 35936 42924 36960
rect 42604 35872 42612 35936
rect 42676 35872 42692 35936
rect 42756 35872 42772 35936
rect 42836 35872 42852 35936
rect 42916 35872 42924 35936
rect 42604 34848 42924 35872
rect 42604 34784 42612 34848
rect 42676 34784 42692 34848
rect 42756 34784 42772 34848
rect 42836 34784 42852 34848
rect 42916 34784 42924 34848
rect 42604 33954 42924 34784
rect 42604 33760 42646 33954
rect 42882 33760 42924 33954
rect 42604 33696 42612 33760
rect 42676 33696 42692 33718
rect 42756 33696 42772 33718
rect 42836 33696 42852 33718
rect 42916 33696 42924 33760
rect 42604 32672 42924 33696
rect 42604 32608 42612 32672
rect 42676 32608 42692 32672
rect 42756 32608 42772 32672
rect 42836 32608 42852 32672
rect 42916 32608 42924 32672
rect 42604 31584 42924 32608
rect 42604 31520 42612 31584
rect 42676 31520 42692 31584
rect 42756 31520 42772 31584
rect 42836 31520 42852 31584
rect 42916 31520 42924 31584
rect 42604 30496 42924 31520
rect 42604 30432 42612 30496
rect 42676 30432 42692 30496
rect 42756 30432 42772 30496
rect 42836 30432 42852 30496
rect 42916 30432 42924 30496
rect 42604 29408 42924 30432
rect 42604 29344 42612 29408
rect 42676 29344 42692 29408
rect 42756 29344 42772 29408
rect 42836 29344 42852 29408
rect 42916 29344 42924 29408
rect 42604 28954 42924 29344
rect 42604 28718 42646 28954
rect 42882 28718 42924 28954
rect 42604 28320 42924 28718
rect 42604 28256 42612 28320
rect 42676 28256 42692 28320
rect 42756 28256 42772 28320
rect 42836 28256 42852 28320
rect 42916 28256 42924 28320
rect 42604 27232 42924 28256
rect 42604 27168 42612 27232
rect 42676 27168 42692 27232
rect 42756 27168 42772 27232
rect 42836 27168 42852 27232
rect 42916 27168 42924 27232
rect 42604 26144 42924 27168
rect 42604 26080 42612 26144
rect 42676 26080 42692 26144
rect 42756 26080 42772 26144
rect 42836 26080 42852 26144
rect 42916 26080 42924 26144
rect 42604 25056 42924 26080
rect 42604 24992 42612 25056
rect 42676 24992 42692 25056
rect 42756 24992 42772 25056
rect 42836 24992 42852 25056
rect 42916 24992 42924 25056
rect 42604 23968 42924 24992
rect 42604 23904 42612 23968
rect 42676 23954 42692 23968
rect 42756 23954 42772 23968
rect 42836 23954 42852 23968
rect 42916 23904 42924 23968
rect 42604 23718 42646 23904
rect 42882 23718 42924 23904
rect 42604 22880 42924 23718
rect 42604 22816 42612 22880
rect 42676 22816 42692 22880
rect 42756 22816 42772 22880
rect 42836 22816 42852 22880
rect 42916 22816 42924 22880
rect 42604 21792 42924 22816
rect 42604 21728 42612 21792
rect 42676 21728 42692 21792
rect 42756 21728 42772 21792
rect 42836 21728 42852 21792
rect 42916 21728 42924 21792
rect 42604 20704 42924 21728
rect 42604 20640 42612 20704
rect 42676 20640 42692 20704
rect 42756 20640 42772 20704
rect 42836 20640 42852 20704
rect 42916 20640 42924 20704
rect 42604 19616 42924 20640
rect 42604 19552 42612 19616
rect 42676 19552 42692 19616
rect 42756 19552 42772 19616
rect 42836 19552 42852 19616
rect 42916 19552 42924 19616
rect 42604 18954 42924 19552
rect 42604 18718 42646 18954
rect 42882 18718 42924 18954
rect 42604 18528 42924 18718
rect 42604 18464 42612 18528
rect 42676 18464 42692 18528
rect 42756 18464 42772 18528
rect 42836 18464 42852 18528
rect 42916 18464 42924 18528
rect 42604 17440 42924 18464
rect 42604 17376 42612 17440
rect 42676 17376 42692 17440
rect 42756 17376 42772 17440
rect 42836 17376 42852 17440
rect 42916 17376 42924 17440
rect 42604 16352 42924 17376
rect 42604 16288 42612 16352
rect 42676 16288 42692 16352
rect 42756 16288 42772 16352
rect 42836 16288 42852 16352
rect 42916 16288 42924 16352
rect 42604 15264 42924 16288
rect 42604 15200 42612 15264
rect 42676 15200 42692 15264
rect 42756 15200 42772 15264
rect 42836 15200 42852 15264
rect 42916 15200 42924 15264
rect 42604 14176 42924 15200
rect 42604 14112 42612 14176
rect 42676 14112 42692 14176
rect 42756 14112 42772 14176
rect 42836 14112 42852 14176
rect 42916 14112 42924 14176
rect 42604 13954 42924 14112
rect 42604 13718 42646 13954
rect 42882 13718 42924 13954
rect 42604 13088 42924 13718
rect 42604 13024 42612 13088
rect 42676 13024 42692 13088
rect 42756 13024 42772 13088
rect 42836 13024 42852 13088
rect 42916 13024 42924 13088
rect 42604 12000 42924 13024
rect 42604 11936 42612 12000
rect 42676 11936 42692 12000
rect 42756 11936 42772 12000
rect 42836 11936 42852 12000
rect 42916 11936 42924 12000
rect 42604 10912 42924 11936
rect 42604 10848 42612 10912
rect 42676 10848 42692 10912
rect 42756 10848 42772 10912
rect 42836 10848 42852 10912
rect 42916 10848 42924 10912
rect 42604 9824 42924 10848
rect 42604 9760 42612 9824
rect 42676 9760 42692 9824
rect 42756 9760 42772 9824
rect 42836 9760 42852 9824
rect 42916 9760 42924 9824
rect 42604 8954 42924 9760
rect 42604 8736 42646 8954
rect 42882 8736 42924 8954
rect 42604 8672 42612 8736
rect 42676 8672 42692 8718
rect 42756 8672 42772 8718
rect 42836 8672 42852 8718
rect 42916 8672 42924 8736
rect 42604 7648 42924 8672
rect 42604 7584 42612 7648
rect 42676 7584 42692 7648
rect 42756 7584 42772 7648
rect 42836 7584 42852 7648
rect 42916 7584 42924 7648
rect 42604 6560 42924 7584
rect 42604 6496 42612 6560
rect 42676 6496 42692 6560
rect 42756 6496 42772 6560
rect 42836 6496 42852 6560
rect 42916 6496 42924 6560
rect 42604 5472 42924 6496
rect 42604 5408 42612 5472
rect 42676 5408 42692 5472
rect 42756 5408 42772 5472
rect 42836 5408 42852 5472
rect 42916 5408 42924 5472
rect 42604 4384 42924 5408
rect 42604 4320 42612 4384
rect 42676 4320 42692 4384
rect 42756 4320 42772 4384
rect 42836 4320 42852 4384
rect 42916 4320 42924 4384
rect 42604 3954 42924 4320
rect 42604 3718 42646 3954
rect 42882 3718 42924 3954
rect 42604 3296 42924 3718
rect 42604 3232 42612 3296
rect 42676 3232 42692 3296
rect 42756 3232 42772 3296
rect 42836 3232 42852 3296
rect 42916 3232 42924 3296
rect 42604 2208 42924 3232
rect 42604 2144 42612 2208
rect 42676 2144 42692 2208
rect 42756 2144 42772 2208
rect 42836 2144 42852 2208
rect 42916 2144 42924 2208
rect 42604 2128 42924 2144
rect 46944 57152 47264 57712
rect 46944 57088 46952 57152
rect 47016 57088 47032 57152
rect 47096 57088 47112 57152
rect 47176 57088 47192 57152
rect 47256 57088 47264 57152
rect 46944 56064 47264 57088
rect 46944 56000 46952 56064
rect 47016 56000 47032 56064
rect 47096 56000 47112 56064
rect 47176 56000 47192 56064
rect 47256 56000 47264 56064
rect 46944 54976 47264 56000
rect 46944 54912 46952 54976
rect 47016 54912 47032 54976
rect 47096 54912 47112 54976
rect 47176 54912 47192 54976
rect 47256 54912 47264 54976
rect 46944 53888 47264 54912
rect 46944 53824 46952 53888
rect 47016 53824 47032 53888
rect 47096 53824 47112 53888
rect 47176 53824 47192 53888
rect 47256 53824 47264 53888
rect 46944 53294 47264 53824
rect 46944 53058 46986 53294
rect 47222 53058 47264 53294
rect 46944 52800 47264 53058
rect 46944 52736 46952 52800
rect 47016 52736 47032 52800
rect 47096 52736 47112 52800
rect 47176 52736 47192 52800
rect 47256 52736 47264 52800
rect 46944 51712 47264 52736
rect 46944 51648 46952 51712
rect 47016 51648 47032 51712
rect 47096 51648 47112 51712
rect 47176 51648 47192 51712
rect 47256 51648 47264 51712
rect 46944 50624 47264 51648
rect 46944 50560 46952 50624
rect 47016 50560 47032 50624
rect 47096 50560 47112 50624
rect 47176 50560 47192 50624
rect 47256 50560 47264 50624
rect 46944 49536 47264 50560
rect 46944 49472 46952 49536
rect 47016 49472 47032 49536
rect 47096 49472 47112 49536
rect 47176 49472 47192 49536
rect 47256 49472 47264 49536
rect 46944 48448 47264 49472
rect 46944 48384 46952 48448
rect 47016 48384 47032 48448
rect 47096 48384 47112 48448
rect 47176 48384 47192 48448
rect 47256 48384 47264 48448
rect 46944 48294 47264 48384
rect 46944 48058 46986 48294
rect 47222 48058 47264 48294
rect 46944 47360 47264 48058
rect 46944 47296 46952 47360
rect 47016 47296 47032 47360
rect 47096 47296 47112 47360
rect 47176 47296 47192 47360
rect 47256 47296 47264 47360
rect 46944 46272 47264 47296
rect 46944 46208 46952 46272
rect 47016 46208 47032 46272
rect 47096 46208 47112 46272
rect 47176 46208 47192 46272
rect 47256 46208 47264 46272
rect 46944 45184 47264 46208
rect 46944 45120 46952 45184
rect 47016 45120 47032 45184
rect 47096 45120 47112 45184
rect 47176 45120 47192 45184
rect 47256 45120 47264 45184
rect 46944 44096 47264 45120
rect 46944 44032 46952 44096
rect 47016 44032 47032 44096
rect 47096 44032 47112 44096
rect 47176 44032 47192 44096
rect 47256 44032 47264 44096
rect 46944 43294 47264 44032
rect 46944 43058 46986 43294
rect 47222 43058 47264 43294
rect 46944 43008 47264 43058
rect 46944 42944 46952 43008
rect 47016 42944 47032 43008
rect 47096 42944 47112 43008
rect 47176 42944 47192 43008
rect 47256 42944 47264 43008
rect 46944 41920 47264 42944
rect 46944 41856 46952 41920
rect 47016 41856 47032 41920
rect 47096 41856 47112 41920
rect 47176 41856 47192 41920
rect 47256 41856 47264 41920
rect 46944 40832 47264 41856
rect 46944 40768 46952 40832
rect 47016 40768 47032 40832
rect 47096 40768 47112 40832
rect 47176 40768 47192 40832
rect 47256 40768 47264 40832
rect 46944 39744 47264 40768
rect 46944 39680 46952 39744
rect 47016 39680 47032 39744
rect 47096 39680 47112 39744
rect 47176 39680 47192 39744
rect 47256 39680 47264 39744
rect 46944 38656 47264 39680
rect 46944 38592 46952 38656
rect 47016 38592 47032 38656
rect 47096 38592 47112 38656
rect 47176 38592 47192 38656
rect 47256 38592 47264 38656
rect 46944 38294 47264 38592
rect 46944 38058 46986 38294
rect 47222 38058 47264 38294
rect 46944 37568 47264 38058
rect 46944 37504 46952 37568
rect 47016 37504 47032 37568
rect 47096 37504 47112 37568
rect 47176 37504 47192 37568
rect 47256 37504 47264 37568
rect 46944 36480 47264 37504
rect 46944 36416 46952 36480
rect 47016 36416 47032 36480
rect 47096 36416 47112 36480
rect 47176 36416 47192 36480
rect 47256 36416 47264 36480
rect 46944 35392 47264 36416
rect 46944 35328 46952 35392
rect 47016 35328 47032 35392
rect 47096 35328 47112 35392
rect 47176 35328 47192 35392
rect 47256 35328 47264 35392
rect 46944 34304 47264 35328
rect 46944 34240 46952 34304
rect 47016 34240 47032 34304
rect 47096 34240 47112 34304
rect 47176 34240 47192 34304
rect 47256 34240 47264 34304
rect 46944 33294 47264 34240
rect 46944 33216 46986 33294
rect 47222 33216 47264 33294
rect 46944 33152 46952 33216
rect 47256 33152 47264 33216
rect 46944 33058 46986 33152
rect 47222 33058 47264 33152
rect 46944 32128 47264 33058
rect 46944 32064 46952 32128
rect 47016 32064 47032 32128
rect 47096 32064 47112 32128
rect 47176 32064 47192 32128
rect 47256 32064 47264 32128
rect 46944 31040 47264 32064
rect 46944 30976 46952 31040
rect 47016 30976 47032 31040
rect 47096 30976 47112 31040
rect 47176 30976 47192 31040
rect 47256 30976 47264 31040
rect 46944 29952 47264 30976
rect 46944 29888 46952 29952
rect 47016 29888 47032 29952
rect 47096 29888 47112 29952
rect 47176 29888 47192 29952
rect 47256 29888 47264 29952
rect 46944 28864 47264 29888
rect 46944 28800 46952 28864
rect 47016 28800 47032 28864
rect 47096 28800 47112 28864
rect 47176 28800 47192 28864
rect 47256 28800 47264 28864
rect 46944 28294 47264 28800
rect 46944 28058 46986 28294
rect 47222 28058 47264 28294
rect 46944 27776 47264 28058
rect 46944 27712 46952 27776
rect 47016 27712 47032 27776
rect 47096 27712 47112 27776
rect 47176 27712 47192 27776
rect 47256 27712 47264 27776
rect 46944 26688 47264 27712
rect 46944 26624 46952 26688
rect 47016 26624 47032 26688
rect 47096 26624 47112 26688
rect 47176 26624 47192 26688
rect 47256 26624 47264 26688
rect 46944 25600 47264 26624
rect 46944 25536 46952 25600
rect 47016 25536 47032 25600
rect 47096 25536 47112 25600
rect 47176 25536 47192 25600
rect 47256 25536 47264 25600
rect 46944 24512 47264 25536
rect 46944 24448 46952 24512
rect 47016 24448 47032 24512
rect 47096 24448 47112 24512
rect 47176 24448 47192 24512
rect 47256 24448 47264 24512
rect 46944 23424 47264 24448
rect 46944 23360 46952 23424
rect 47016 23360 47032 23424
rect 47096 23360 47112 23424
rect 47176 23360 47192 23424
rect 47256 23360 47264 23424
rect 46944 23294 47264 23360
rect 46944 23058 46986 23294
rect 47222 23058 47264 23294
rect 46944 22336 47264 23058
rect 46944 22272 46952 22336
rect 47016 22272 47032 22336
rect 47096 22272 47112 22336
rect 47176 22272 47192 22336
rect 47256 22272 47264 22336
rect 46944 21248 47264 22272
rect 46944 21184 46952 21248
rect 47016 21184 47032 21248
rect 47096 21184 47112 21248
rect 47176 21184 47192 21248
rect 47256 21184 47264 21248
rect 46944 20160 47264 21184
rect 46944 20096 46952 20160
rect 47016 20096 47032 20160
rect 47096 20096 47112 20160
rect 47176 20096 47192 20160
rect 47256 20096 47264 20160
rect 46944 19072 47264 20096
rect 46944 19008 46952 19072
rect 47016 19008 47032 19072
rect 47096 19008 47112 19072
rect 47176 19008 47192 19072
rect 47256 19008 47264 19072
rect 46944 18294 47264 19008
rect 46944 18058 46986 18294
rect 47222 18058 47264 18294
rect 46944 17984 47264 18058
rect 46944 17920 46952 17984
rect 47016 17920 47032 17984
rect 47096 17920 47112 17984
rect 47176 17920 47192 17984
rect 47256 17920 47264 17984
rect 46944 16896 47264 17920
rect 46944 16832 46952 16896
rect 47016 16832 47032 16896
rect 47096 16832 47112 16896
rect 47176 16832 47192 16896
rect 47256 16832 47264 16896
rect 46944 15808 47264 16832
rect 46944 15744 46952 15808
rect 47016 15744 47032 15808
rect 47096 15744 47112 15808
rect 47176 15744 47192 15808
rect 47256 15744 47264 15808
rect 46944 14720 47264 15744
rect 46944 14656 46952 14720
rect 47016 14656 47032 14720
rect 47096 14656 47112 14720
rect 47176 14656 47192 14720
rect 47256 14656 47264 14720
rect 46944 13632 47264 14656
rect 46944 13568 46952 13632
rect 47016 13568 47032 13632
rect 47096 13568 47112 13632
rect 47176 13568 47192 13632
rect 47256 13568 47264 13632
rect 46944 13294 47264 13568
rect 46944 13058 46986 13294
rect 47222 13058 47264 13294
rect 46944 12544 47264 13058
rect 46944 12480 46952 12544
rect 47016 12480 47032 12544
rect 47096 12480 47112 12544
rect 47176 12480 47192 12544
rect 47256 12480 47264 12544
rect 46944 11456 47264 12480
rect 46944 11392 46952 11456
rect 47016 11392 47032 11456
rect 47096 11392 47112 11456
rect 47176 11392 47192 11456
rect 47256 11392 47264 11456
rect 46944 10368 47264 11392
rect 46944 10304 46952 10368
rect 47016 10304 47032 10368
rect 47096 10304 47112 10368
rect 47176 10304 47192 10368
rect 47256 10304 47264 10368
rect 46944 9280 47264 10304
rect 46944 9216 46952 9280
rect 47016 9216 47032 9280
rect 47096 9216 47112 9280
rect 47176 9216 47192 9280
rect 47256 9216 47264 9280
rect 46944 8294 47264 9216
rect 46944 8192 46986 8294
rect 47222 8192 47264 8294
rect 46944 8128 46952 8192
rect 47256 8128 47264 8192
rect 46944 8058 46986 8128
rect 47222 8058 47264 8128
rect 46944 7104 47264 8058
rect 46944 7040 46952 7104
rect 47016 7040 47032 7104
rect 47096 7040 47112 7104
rect 47176 7040 47192 7104
rect 47256 7040 47264 7104
rect 46944 6016 47264 7040
rect 46944 5952 46952 6016
rect 47016 5952 47032 6016
rect 47096 5952 47112 6016
rect 47176 5952 47192 6016
rect 47256 5952 47264 6016
rect 46944 4928 47264 5952
rect 46944 4864 46952 4928
rect 47016 4864 47032 4928
rect 47096 4864 47112 4928
rect 47176 4864 47192 4928
rect 47256 4864 47264 4928
rect 46944 3840 47264 4864
rect 46944 3776 46952 3840
rect 47016 3776 47032 3840
rect 47096 3776 47112 3840
rect 47176 3776 47192 3840
rect 47256 3776 47264 3840
rect 46944 3294 47264 3776
rect 46944 3058 46986 3294
rect 47222 3058 47264 3294
rect 46944 2752 47264 3058
rect 46944 2688 46952 2752
rect 47016 2688 47032 2752
rect 47096 2688 47112 2752
rect 47176 2688 47192 2752
rect 47256 2688 47264 2752
rect 46944 2128 47264 2688
rect 47604 57696 47924 57712
rect 47604 57632 47612 57696
rect 47676 57632 47692 57696
rect 47756 57632 47772 57696
rect 47836 57632 47852 57696
rect 47916 57632 47924 57696
rect 47604 56608 47924 57632
rect 47604 56544 47612 56608
rect 47676 56544 47692 56608
rect 47756 56544 47772 56608
rect 47836 56544 47852 56608
rect 47916 56544 47924 56608
rect 47604 55520 47924 56544
rect 47604 55456 47612 55520
rect 47676 55456 47692 55520
rect 47756 55456 47772 55520
rect 47836 55456 47852 55520
rect 47916 55456 47924 55520
rect 47604 54432 47924 55456
rect 47604 54368 47612 54432
rect 47676 54368 47692 54432
rect 47756 54368 47772 54432
rect 47836 54368 47852 54432
rect 47916 54368 47924 54432
rect 47604 53954 47924 54368
rect 47604 53718 47646 53954
rect 47882 53718 47924 53954
rect 47604 53344 47924 53718
rect 47604 53280 47612 53344
rect 47676 53280 47692 53344
rect 47756 53280 47772 53344
rect 47836 53280 47852 53344
rect 47916 53280 47924 53344
rect 47604 52256 47924 53280
rect 47604 52192 47612 52256
rect 47676 52192 47692 52256
rect 47756 52192 47772 52256
rect 47836 52192 47852 52256
rect 47916 52192 47924 52256
rect 47604 51168 47924 52192
rect 47604 51104 47612 51168
rect 47676 51104 47692 51168
rect 47756 51104 47772 51168
rect 47836 51104 47852 51168
rect 47916 51104 47924 51168
rect 47604 50080 47924 51104
rect 47604 50016 47612 50080
rect 47676 50016 47692 50080
rect 47756 50016 47772 50080
rect 47836 50016 47852 50080
rect 47916 50016 47924 50080
rect 47604 48992 47924 50016
rect 47604 48928 47612 48992
rect 47676 48954 47692 48992
rect 47756 48954 47772 48992
rect 47836 48954 47852 48992
rect 47916 48928 47924 48992
rect 47604 48718 47646 48928
rect 47882 48718 47924 48928
rect 47604 47904 47924 48718
rect 47604 47840 47612 47904
rect 47676 47840 47692 47904
rect 47756 47840 47772 47904
rect 47836 47840 47852 47904
rect 47916 47840 47924 47904
rect 47604 46816 47924 47840
rect 47604 46752 47612 46816
rect 47676 46752 47692 46816
rect 47756 46752 47772 46816
rect 47836 46752 47852 46816
rect 47916 46752 47924 46816
rect 47604 45728 47924 46752
rect 47604 45664 47612 45728
rect 47676 45664 47692 45728
rect 47756 45664 47772 45728
rect 47836 45664 47852 45728
rect 47916 45664 47924 45728
rect 47604 44640 47924 45664
rect 47604 44576 47612 44640
rect 47676 44576 47692 44640
rect 47756 44576 47772 44640
rect 47836 44576 47852 44640
rect 47916 44576 47924 44640
rect 47604 43954 47924 44576
rect 47604 43718 47646 43954
rect 47882 43718 47924 43954
rect 47604 43552 47924 43718
rect 47604 43488 47612 43552
rect 47676 43488 47692 43552
rect 47756 43488 47772 43552
rect 47836 43488 47852 43552
rect 47916 43488 47924 43552
rect 47604 42464 47924 43488
rect 47604 42400 47612 42464
rect 47676 42400 47692 42464
rect 47756 42400 47772 42464
rect 47836 42400 47852 42464
rect 47916 42400 47924 42464
rect 47604 41376 47924 42400
rect 47604 41312 47612 41376
rect 47676 41312 47692 41376
rect 47756 41312 47772 41376
rect 47836 41312 47852 41376
rect 47916 41312 47924 41376
rect 47604 40288 47924 41312
rect 47604 40224 47612 40288
rect 47676 40224 47692 40288
rect 47756 40224 47772 40288
rect 47836 40224 47852 40288
rect 47916 40224 47924 40288
rect 47604 39200 47924 40224
rect 47604 39136 47612 39200
rect 47676 39136 47692 39200
rect 47756 39136 47772 39200
rect 47836 39136 47852 39200
rect 47916 39136 47924 39200
rect 47604 38954 47924 39136
rect 47604 38718 47646 38954
rect 47882 38718 47924 38954
rect 47604 38112 47924 38718
rect 47604 38048 47612 38112
rect 47676 38048 47692 38112
rect 47756 38048 47772 38112
rect 47836 38048 47852 38112
rect 47916 38048 47924 38112
rect 47604 37024 47924 38048
rect 47604 36960 47612 37024
rect 47676 36960 47692 37024
rect 47756 36960 47772 37024
rect 47836 36960 47852 37024
rect 47916 36960 47924 37024
rect 47604 35936 47924 36960
rect 47604 35872 47612 35936
rect 47676 35872 47692 35936
rect 47756 35872 47772 35936
rect 47836 35872 47852 35936
rect 47916 35872 47924 35936
rect 47604 34848 47924 35872
rect 47604 34784 47612 34848
rect 47676 34784 47692 34848
rect 47756 34784 47772 34848
rect 47836 34784 47852 34848
rect 47916 34784 47924 34848
rect 47604 33954 47924 34784
rect 47604 33760 47646 33954
rect 47882 33760 47924 33954
rect 47604 33696 47612 33760
rect 47676 33696 47692 33718
rect 47756 33696 47772 33718
rect 47836 33696 47852 33718
rect 47916 33696 47924 33760
rect 47604 32672 47924 33696
rect 47604 32608 47612 32672
rect 47676 32608 47692 32672
rect 47756 32608 47772 32672
rect 47836 32608 47852 32672
rect 47916 32608 47924 32672
rect 47604 31584 47924 32608
rect 47604 31520 47612 31584
rect 47676 31520 47692 31584
rect 47756 31520 47772 31584
rect 47836 31520 47852 31584
rect 47916 31520 47924 31584
rect 47604 30496 47924 31520
rect 47604 30432 47612 30496
rect 47676 30432 47692 30496
rect 47756 30432 47772 30496
rect 47836 30432 47852 30496
rect 47916 30432 47924 30496
rect 47604 29408 47924 30432
rect 47604 29344 47612 29408
rect 47676 29344 47692 29408
rect 47756 29344 47772 29408
rect 47836 29344 47852 29408
rect 47916 29344 47924 29408
rect 47604 28954 47924 29344
rect 47604 28718 47646 28954
rect 47882 28718 47924 28954
rect 47604 28320 47924 28718
rect 47604 28256 47612 28320
rect 47676 28256 47692 28320
rect 47756 28256 47772 28320
rect 47836 28256 47852 28320
rect 47916 28256 47924 28320
rect 47604 27232 47924 28256
rect 47604 27168 47612 27232
rect 47676 27168 47692 27232
rect 47756 27168 47772 27232
rect 47836 27168 47852 27232
rect 47916 27168 47924 27232
rect 47604 26144 47924 27168
rect 47604 26080 47612 26144
rect 47676 26080 47692 26144
rect 47756 26080 47772 26144
rect 47836 26080 47852 26144
rect 47916 26080 47924 26144
rect 47604 25056 47924 26080
rect 47604 24992 47612 25056
rect 47676 24992 47692 25056
rect 47756 24992 47772 25056
rect 47836 24992 47852 25056
rect 47916 24992 47924 25056
rect 47604 23968 47924 24992
rect 47604 23904 47612 23968
rect 47676 23954 47692 23968
rect 47756 23954 47772 23968
rect 47836 23954 47852 23968
rect 47916 23904 47924 23968
rect 47604 23718 47646 23904
rect 47882 23718 47924 23904
rect 47604 22880 47924 23718
rect 47604 22816 47612 22880
rect 47676 22816 47692 22880
rect 47756 22816 47772 22880
rect 47836 22816 47852 22880
rect 47916 22816 47924 22880
rect 47604 21792 47924 22816
rect 47604 21728 47612 21792
rect 47676 21728 47692 21792
rect 47756 21728 47772 21792
rect 47836 21728 47852 21792
rect 47916 21728 47924 21792
rect 47604 20704 47924 21728
rect 47604 20640 47612 20704
rect 47676 20640 47692 20704
rect 47756 20640 47772 20704
rect 47836 20640 47852 20704
rect 47916 20640 47924 20704
rect 47604 19616 47924 20640
rect 47604 19552 47612 19616
rect 47676 19552 47692 19616
rect 47756 19552 47772 19616
rect 47836 19552 47852 19616
rect 47916 19552 47924 19616
rect 47604 18954 47924 19552
rect 47604 18718 47646 18954
rect 47882 18718 47924 18954
rect 47604 18528 47924 18718
rect 47604 18464 47612 18528
rect 47676 18464 47692 18528
rect 47756 18464 47772 18528
rect 47836 18464 47852 18528
rect 47916 18464 47924 18528
rect 47604 17440 47924 18464
rect 47604 17376 47612 17440
rect 47676 17376 47692 17440
rect 47756 17376 47772 17440
rect 47836 17376 47852 17440
rect 47916 17376 47924 17440
rect 47604 16352 47924 17376
rect 47604 16288 47612 16352
rect 47676 16288 47692 16352
rect 47756 16288 47772 16352
rect 47836 16288 47852 16352
rect 47916 16288 47924 16352
rect 47604 15264 47924 16288
rect 47604 15200 47612 15264
rect 47676 15200 47692 15264
rect 47756 15200 47772 15264
rect 47836 15200 47852 15264
rect 47916 15200 47924 15264
rect 47604 14176 47924 15200
rect 47604 14112 47612 14176
rect 47676 14112 47692 14176
rect 47756 14112 47772 14176
rect 47836 14112 47852 14176
rect 47916 14112 47924 14176
rect 47604 13954 47924 14112
rect 47604 13718 47646 13954
rect 47882 13718 47924 13954
rect 47604 13088 47924 13718
rect 47604 13024 47612 13088
rect 47676 13024 47692 13088
rect 47756 13024 47772 13088
rect 47836 13024 47852 13088
rect 47916 13024 47924 13088
rect 47604 12000 47924 13024
rect 47604 11936 47612 12000
rect 47676 11936 47692 12000
rect 47756 11936 47772 12000
rect 47836 11936 47852 12000
rect 47916 11936 47924 12000
rect 47604 10912 47924 11936
rect 47604 10848 47612 10912
rect 47676 10848 47692 10912
rect 47756 10848 47772 10912
rect 47836 10848 47852 10912
rect 47916 10848 47924 10912
rect 47604 9824 47924 10848
rect 47604 9760 47612 9824
rect 47676 9760 47692 9824
rect 47756 9760 47772 9824
rect 47836 9760 47852 9824
rect 47916 9760 47924 9824
rect 47604 8954 47924 9760
rect 47604 8736 47646 8954
rect 47882 8736 47924 8954
rect 47604 8672 47612 8736
rect 47676 8672 47692 8718
rect 47756 8672 47772 8718
rect 47836 8672 47852 8718
rect 47916 8672 47924 8736
rect 47604 7648 47924 8672
rect 47604 7584 47612 7648
rect 47676 7584 47692 7648
rect 47756 7584 47772 7648
rect 47836 7584 47852 7648
rect 47916 7584 47924 7648
rect 47604 6560 47924 7584
rect 47604 6496 47612 6560
rect 47676 6496 47692 6560
rect 47756 6496 47772 6560
rect 47836 6496 47852 6560
rect 47916 6496 47924 6560
rect 47604 5472 47924 6496
rect 47604 5408 47612 5472
rect 47676 5408 47692 5472
rect 47756 5408 47772 5472
rect 47836 5408 47852 5472
rect 47916 5408 47924 5472
rect 47604 4384 47924 5408
rect 47604 4320 47612 4384
rect 47676 4320 47692 4384
rect 47756 4320 47772 4384
rect 47836 4320 47852 4384
rect 47916 4320 47924 4384
rect 47604 3954 47924 4320
rect 47604 3718 47646 3954
rect 47882 3718 47924 3954
rect 47604 3296 47924 3718
rect 47604 3232 47612 3296
rect 47676 3232 47692 3296
rect 47756 3232 47772 3296
rect 47836 3232 47852 3296
rect 47916 3232 47924 3296
rect 47604 2208 47924 3232
rect 47604 2144 47612 2208
rect 47676 2144 47692 2208
rect 47756 2144 47772 2208
rect 47836 2144 47852 2208
rect 47916 2144 47924 2208
rect 47604 2128 47924 2144
rect 51944 57152 52264 57712
rect 51944 57088 51952 57152
rect 52016 57088 52032 57152
rect 52096 57088 52112 57152
rect 52176 57088 52192 57152
rect 52256 57088 52264 57152
rect 51944 56064 52264 57088
rect 51944 56000 51952 56064
rect 52016 56000 52032 56064
rect 52096 56000 52112 56064
rect 52176 56000 52192 56064
rect 52256 56000 52264 56064
rect 51944 54976 52264 56000
rect 51944 54912 51952 54976
rect 52016 54912 52032 54976
rect 52096 54912 52112 54976
rect 52176 54912 52192 54976
rect 52256 54912 52264 54976
rect 51944 53888 52264 54912
rect 51944 53824 51952 53888
rect 52016 53824 52032 53888
rect 52096 53824 52112 53888
rect 52176 53824 52192 53888
rect 52256 53824 52264 53888
rect 51944 53294 52264 53824
rect 51944 53058 51986 53294
rect 52222 53058 52264 53294
rect 51944 52800 52264 53058
rect 51944 52736 51952 52800
rect 52016 52736 52032 52800
rect 52096 52736 52112 52800
rect 52176 52736 52192 52800
rect 52256 52736 52264 52800
rect 51944 51712 52264 52736
rect 51944 51648 51952 51712
rect 52016 51648 52032 51712
rect 52096 51648 52112 51712
rect 52176 51648 52192 51712
rect 52256 51648 52264 51712
rect 51944 50624 52264 51648
rect 51944 50560 51952 50624
rect 52016 50560 52032 50624
rect 52096 50560 52112 50624
rect 52176 50560 52192 50624
rect 52256 50560 52264 50624
rect 51944 49536 52264 50560
rect 51944 49472 51952 49536
rect 52016 49472 52032 49536
rect 52096 49472 52112 49536
rect 52176 49472 52192 49536
rect 52256 49472 52264 49536
rect 51944 48448 52264 49472
rect 51944 48384 51952 48448
rect 52016 48384 52032 48448
rect 52096 48384 52112 48448
rect 52176 48384 52192 48448
rect 52256 48384 52264 48448
rect 51944 48294 52264 48384
rect 51944 48058 51986 48294
rect 52222 48058 52264 48294
rect 51944 47360 52264 48058
rect 51944 47296 51952 47360
rect 52016 47296 52032 47360
rect 52096 47296 52112 47360
rect 52176 47296 52192 47360
rect 52256 47296 52264 47360
rect 51944 46272 52264 47296
rect 51944 46208 51952 46272
rect 52016 46208 52032 46272
rect 52096 46208 52112 46272
rect 52176 46208 52192 46272
rect 52256 46208 52264 46272
rect 51944 45184 52264 46208
rect 51944 45120 51952 45184
rect 52016 45120 52032 45184
rect 52096 45120 52112 45184
rect 52176 45120 52192 45184
rect 52256 45120 52264 45184
rect 51944 44096 52264 45120
rect 51944 44032 51952 44096
rect 52016 44032 52032 44096
rect 52096 44032 52112 44096
rect 52176 44032 52192 44096
rect 52256 44032 52264 44096
rect 51944 43294 52264 44032
rect 51944 43058 51986 43294
rect 52222 43058 52264 43294
rect 51944 43008 52264 43058
rect 51944 42944 51952 43008
rect 52016 42944 52032 43008
rect 52096 42944 52112 43008
rect 52176 42944 52192 43008
rect 52256 42944 52264 43008
rect 51944 41920 52264 42944
rect 51944 41856 51952 41920
rect 52016 41856 52032 41920
rect 52096 41856 52112 41920
rect 52176 41856 52192 41920
rect 52256 41856 52264 41920
rect 51944 40832 52264 41856
rect 51944 40768 51952 40832
rect 52016 40768 52032 40832
rect 52096 40768 52112 40832
rect 52176 40768 52192 40832
rect 52256 40768 52264 40832
rect 51944 39744 52264 40768
rect 51944 39680 51952 39744
rect 52016 39680 52032 39744
rect 52096 39680 52112 39744
rect 52176 39680 52192 39744
rect 52256 39680 52264 39744
rect 51944 38656 52264 39680
rect 51944 38592 51952 38656
rect 52016 38592 52032 38656
rect 52096 38592 52112 38656
rect 52176 38592 52192 38656
rect 52256 38592 52264 38656
rect 51944 38294 52264 38592
rect 51944 38058 51986 38294
rect 52222 38058 52264 38294
rect 51944 37568 52264 38058
rect 51944 37504 51952 37568
rect 52016 37504 52032 37568
rect 52096 37504 52112 37568
rect 52176 37504 52192 37568
rect 52256 37504 52264 37568
rect 51944 36480 52264 37504
rect 51944 36416 51952 36480
rect 52016 36416 52032 36480
rect 52096 36416 52112 36480
rect 52176 36416 52192 36480
rect 52256 36416 52264 36480
rect 51944 35392 52264 36416
rect 51944 35328 51952 35392
rect 52016 35328 52032 35392
rect 52096 35328 52112 35392
rect 52176 35328 52192 35392
rect 52256 35328 52264 35392
rect 51944 34304 52264 35328
rect 51944 34240 51952 34304
rect 52016 34240 52032 34304
rect 52096 34240 52112 34304
rect 52176 34240 52192 34304
rect 52256 34240 52264 34304
rect 51944 33294 52264 34240
rect 51944 33216 51986 33294
rect 52222 33216 52264 33294
rect 51944 33152 51952 33216
rect 52256 33152 52264 33216
rect 51944 33058 51986 33152
rect 52222 33058 52264 33152
rect 51944 32128 52264 33058
rect 51944 32064 51952 32128
rect 52016 32064 52032 32128
rect 52096 32064 52112 32128
rect 52176 32064 52192 32128
rect 52256 32064 52264 32128
rect 51944 31040 52264 32064
rect 51944 30976 51952 31040
rect 52016 30976 52032 31040
rect 52096 30976 52112 31040
rect 52176 30976 52192 31040
rect 52256 30976 52264 31040
rect 51944 29952 52264 30976
rect 51944 29888 51952 29952
rect 52016 29888 52032 29952
rect 52096 29888 52112 29952
rect 52176 29888 52192 29952
rect 52256 29888 52264 29952
rect 51944 28864 52264 29888
rect 51944 28800 51952 28864
rect 52016 28800 52032 28864
rect 52096 28800 52112 28864
rect 52176 28800 52192 28864
rect 52256 28800 52264 28864
rect 51944 28294 52264 28800
rect 51944 28058 51986 28294
rect 52222 28058 52264 28294
rect 51944 27776 52264 28058
rect 51944 27712 51952 27776
rect 52016 27712 52032 27776
rect 52096 27712 52112 27776
rect 52176 27712 52192 27776
rect 52256 27712 52264 27776
rect 51944 26688 52264 27712
rect 51944 26624 51952 26688
rect 52016 26624 52032 26688
rect 52096 26624 52112 26688
rect 52176 26624 52192 26688
rect 52256 26624 52264 26688
rect 51944 25600 52264 26624
rect 51944 25536 51952 25600
rect 52016 25536 52032 25600
rect 52096 25536 52112 25600
rect 52176 25536 52192 25600
rect 52256 25536 52264 25600
rect 51944 24512 52264 25536
rect 51944 24448 51952 24512
rect 52016 24448 52032 24512
rect 52096 24448 52112 24512
rect 52176 24448 52192 24512
rect 52256 24448 52264 24512
rect 51944 23424 52264 24448
rect 51944 23360 51952 23424
rect 52016 23360 52032 23424
rect 52096 23360 52112 23424
rect 52176 23360 52192 23424
rect 52256 23360 52264 23424
rect 51944 23294 52264 23360
rect 51944 23058 51986 23294
rect 52222 23058 52264 23294
rect 51944 22336 52264 23058
rect 51944 22272 51952 22336
rect 52016 22272 52032 22336
rect 52096 22272 52112 22336
rect 52176 22272 52192 22336
rect 52256 22272 52264 22336
rect 51944 21248 52264 22272
rect 51944 21184 51952 21248
rect 52016 21184 52032 21248
rect 52096 21184 52112 21248
rect 52176 21184 52192 21248
rect 52256 21184 52264 21248
rect 51944 20160 52264 21184
rect 51944 20096 51952 20160
rect 52016 20096 52032 20160
rect 52096 20096 52112 20160
rect 52176 20096 52192 20160
rect 52256 20096 52264 20160
rect 51944 19072 52264 20096
rect 51944 19008 51952 19072
rect 52016 19008 52032 19072
rect 52096 19008 52112 19072
rect 52176 19008 52192 19072
rect 52256 19008 52264 19072
rect 51944 18294 52264 19008
rect 51944 18058 51986 18294
rect 52222 18058 52264 18294
rect 51944 17984 52264 18058
rect 51944 17920 51952 17984
rect 52016 17920 52032 17984
rect 52096 17920 52112 17984
rect 52176 17920 52192 17984
rect 52256 17920 52264 17984
rect 51944 16896 52264 17920
rect 51944 16832 51952 16896
rect 52016 16832 52032 16896
rect 52096 16832 52112 16896
rect 52176 16832 52192 16896
rect 52256 16832 52264 16896
rect 51944 15808 52264 16832
rect 51944 15744 51952 15808
rect 52016 15744 52032 15808
rect 52096 15744 52112 15808
rect 52176 15744 52192 15808
rect 52256 15744 52264 15808
rect 51944 14720 52264 15744
rect 51944 14656 51952 14720
rect 52016 14656 52032 14720
rect 52096 14656 52112 14720
rect 52176 14656 52192 14720
rect 52256 14656 52264 14720
rect 51944 13632 52264 14656
rect 51944 13568 51952 13632
rect 52016 13568 52032 13632
rect 52096 13568 52112 13632
rect 52176 13568 52192 13632
rect 52256 13568 52264 13632
rect 51944 13294 52264 13568
rect 51944 13058 51986 13294
rect 52222 13058 52264 13294
rect 51944 12544 52264 13058
rect 51944 12480 51952 12544
rect 52016 12480 52032 12544
rect 52096 12480 52112 12544
rect 52176 12480 52192 12544
rect 52256 12480 52264 12544
rect 51944 11456 52264 12480
rect 51944 11392 51952 11456
rect 52016 11392 52032 11456
rect 52096 11392 52112 11456
rect 52176 11392 52192 11456
rect 52256 11392 52264 11456
rect 51944 10368 52264 11392
rect 51944 10304 51952 10368
rect 52016 10304 52032 10368
rect 52096 10304 52112 10368
rect 52176 10304 52192 10368
rect 52256 10304 52264 10368
rect 51944 9280 52264 10304
rect 51944 9216 51952 9280
rect 52016 9216 52032 9280
rect 52096 9216 52112 9280
rect 52176 9216 52192 9280
rect 52256 9216 52264 9280
rect 51944 8294 52264 9216
rect 51944 8192 51986 8294
rect 52222 8192 52264 8294
rect 51944 8128 51952 8192
rect 52256 8128 52264 8192
rect 51944 8058 51986 8128
rect 52222 8058 52264 8128
rect 51944 7104 52264 8058
rect 51944 7040 51952 7104
rect 52016 7040 52032 7104
rect 52096 7040 52112 7104
rect 52176 7040 52192 7104
rect 52256 7040 52264 7104
rect 51944 6016 52264 7040
rect 51944 5952 51952 6016
rect 52016 5952 52032 6016
rect 52096 5952 52112 6016
rect 52176 5952 52192 6016
rect 52256 5952 52264 6016
rect 51944 4928 52264 5952
rect 51944 4864 51952 4928
rect 52016 4864 52032 4928
rect 52096 4864 52112 4928
rect 52176 4864 52192 4928
rect 52256 4864 52264 4928
rect 51944 3840 52264 4864
rect 51944 3776 51952 3840
rect 52016 3776 52032 3840
rect 52096 3776 52112 3840
rect 52176 3776 52192 3840
rect 52256 3776 52264 3840
rect 51944 3294 52264 3776
rect 51944 3058 51986 3294
rect 52222 3058 52264 3294
rect 51944 2752 52264 3058
rect 51944 2688 51952 2752
rect 52016 2688 52032 2752
rect 52096 2688 52112 2752
rect 52176 2688 52192 2752
rect 52256 2688 52264 2752
rect 51944 2128 52264 2688
rect 52604 57696 52924 57712
rect 52604 57632 52612 57696
rect 52676 57632 52692 57696
rect 52756 57632 52772 57696
rect 52836 57632 52852 57696
rect 52916 57632 52924 57696
rect 52604 56608 52924 57632
rect 52604 56544 52612 56608
rect 52676 56544 52692 56608
rect 52756 56544 52772 56608
rect 52836 56544 52852 56608
rect 52916 56544 52924 56608
rect 52604 55520 52924 56544
rect 52604 55456 52612 55520
rect 52676 55456 52692 55520
rect 52756 55456 52772 55520
rect 52836 55456 52852 55520
rect 52916 55456 52924 55520
rect 52604 54432 52924 55456
rect 52604 54368 52612 54432
rect 52676 54368 52692 54432
rect 52756 54368 52772 54432
rect 52836 54368 52852 54432
rect 52916 54368 52924 54432
rect 52604 53954 52924 54368
rect 52604 53718 52646 53954
rect 52882 53718 52924 53954
rect 52604 53344 52924 53718
rect 52604 53280 52612 53344
rect 52676 53280 52692 53344
rect 52756 53280 52772 53344
rect 52836 53280 52852 53344
rect 52916 53280 52924 53344
rect 52604 52256 52924 53280
rect 52604 52192 52612 52256
rect 52676 52192 52692 52256
rect 52756 52192 52772 52256
rect 52836 52192 52852 52256
rect 52916 52192 52924 52256
rect 52604 51168 52924 52192
rect 52604 51104 52612 51168
rect 52676 51104 52692 51168
rect 52756 51104 52772 51168
rect 52836 51104 52852 51168
rect 52916 51104 52924 51168
rect 52604 50080 52924 51104
rect 52604 50016 52612 50080
rect 52676 50016 52692 50080
rect 52756 50016 52772 50080
rect 52836 50016 52852 50080
rect 52916 50016 52924 50080
rect 52604 48992 52924 50016
rect 52604 48928 52612 48992
rect 52676 48954 52692 48992
rect 52756 48954 52772 48992
rect 52836 48954 52852 48992
rect 52916 48928 52924 48992
rect 52604 48718 52646 48928
rect 52882 48718 52924 48928
rect 52604 47904 52924 48718
rect 52604 47840 52612 47904
rect 52676 47840 52692 47904
rect 52756 47840 52772 47904
rect 52836 47840 52852 47904
rect 52916 47840 52924 47904
rect 52604 46816 52924 47840
rect 52604 46752 52612 46816
rect 52676 46752 52692 46816
rect 52756 46752 52772 46816
rect 52836 46752 52852 46816
rect 52916 46752 52924 46816
rect 52604 45728 52924 46752
rect 52604 45664 52612 45728
rect 52676 45664 52692 45728
rect 52756 45664 52772 45728
rect 52836 45664 52852 45728
rect 52916 45664 52924 45728
rect 52604 44640 52924 45664
rect 52604 44576 52612 44640
rect 52676 44576 52692 44640
rect 52756 44576 52772 44640
rect 52836 44576 52852 44640
rect 52916 44576 52924 44640
rect 52604 43954 52924 44576
rect 52604 43718 52646 43954
rect 52882 43718 52924 43954
rect 52604 43552 52924 43718
rect 52604 43488 52612 43552
rect 52676 43488 52692 43552
rect 52756 43488 52772 43552
rect 52836 43488 52852 43552
rect 52916 43488 52924 43552
rect 52604 42464 52924 43488
rect 52604 42400 52612 42464
rect 52676 42400 52692 42464
rect 52756 42400 52772 42464
rect 52836 42400 52852 42464
rect 52916 42400 52924 42464
rect 52604 41376 52924 42400
rect 52604 41312 52612 41376
rect 52676 41312 52692 41376
rect 52756 41312 52772 41376
rect 52836 41312 52852 41376
rect 52916 41312 52924 41376
rect 52604 40288 52924 41312
rect 52604 40224 52612 40288
rect 52676 40224 52692 40288
rect 52756 40224 52772 40288
rect 52836 40224 52852 40288
rect 52916 40224 52924 40288
rect 52604 39200 52924 40224
rect 52604 39136 52612 39200
rect 52676 39136 52692 39200
rect 52756 39136 52772 39200
rect 52836 39136 52852 39200
rect 52916 39136 52924 39200
rect 52604 38954 52924 39136
rect 52604 38718 52646 38954
rect 52882 38718 52924 38954
rect 52604 38112 52924 38718
rect 52604 38048 52612 38112
rect 52676 38048 52692 38112
rect 52756 38048 52772 38112
rect 52836 38048 52852 38112
rect 52916 38048 52924 38112
rect 52604 37024 52924 38048
rect 52604 36960 52612 37024
rect 52676 36960 52692 37024
rect 52756 36960 52772 37024
rect 52836 36960 52852 37024
rect 52916 36960 52924 37024
rect 52604 35936 52924 36960
rect 52604 35872 52612 35936
rect 52676 35872 52692 35936
rect 52756 35872 52772 35936
rect 52836 35872 52852 35936
rect 52916 35872 52924 35936
rect 52604 34848 52924 35872
rect 52604 34784 52612 34848
rect 52676 34784 52692 34848
rect 52756 34784 52772 34848
rect 52836 34784 52852 34848
rect 52916 34784 52924 34848
rect 52604 33954 52924 34784
rect 52604 33760 52646 33954
rect 52882 33760 52924 33954
rect 52604 33696 52612 33760
rect 52676 33696 52692 33718
rect 52756 33696 52772 33718
rect 52836 33696 52852 33718
rect 52916 33696 52924 33760
rect 52604 32672 52924 33696
rect 52604 32608 52612 32672
rect 52676 32608 52692 32672
rect 52756 32608 52772 32672
rect 52836 32608 52852 32672
rect 52916 32608 52924 32672
rect 52604 31584 52924 32608
rect 52604 31520 52612 31584
rect 52676 31520 52692 31584
rect 52756 31520 52772 31584
rect 52836 31520 52852 31584
rect 52916 31520 52924 31584
rect 52604 30496 52924 31520
rect 52604 30432 52612 30496
rect 52676 30432 52692 30496
rect 52756 30432 52772 30496
rect 52836 30432 52852 30496
rect 52916 30432 52924 30496
rect 52604 29408 52924 30432
rect 52604 29344 52612 29408
rect 52676 29344 52692 29408
rect 52756 29344 52772 29408
rect 52836 29344 52852 29408
rect 52916 29344 52924 29408
rect 52604 28954 52924 29344
rect 52604 28718 52646 28954
rect 52882 28718 52924 28954
rect 52604 28320 52924 28718
rect 52604 28256 52612 28320
rect 52676 28256 52692 28320
rect 52756 28256 52772 28320
rect 52836 28256 52852 28320
rect 52916 28256 52924 28320
rect 52604 27232 52924 28256
rect 52604 27168 52612 27232
rect 52676 27168 52692 27232
rect 52756 27168 52772 27232
rect 52836 27168 52852 27232
rect 52916 27168 52924 27232
rect 52604 26144 52924 27168
rect 52604 26080 52612 26144
rect 52676 26080 52692 26144
rect 52756 26080 52772 26144
rect 52836 26080 52852 26144
rect 52916 26080 52924 26144
rect 52604 25056 52924 26080
rect 52604 24992 52612 25056
rect 52676 24992 52692 25056
rect 52756 24992 52772 25056
rect 52836 24992 52852 25056
rect 52916 24992 52924 25056
rect 52604 23968 52924 24992
rect 52604 23904 52612 23968
rect 52676 23954 52692 23968
rect 52756 23954 52772 23968
rect 52836 23954 52852 23968
rect 52916 23904 52924 23968
rect 52604 23718 52646 23904
rect 52882 23718 52924 23904
rect 52604 22880 52924 23718
rect 52604 22816 52612 22880
rect 52676 22816 52692 22880
rect 52756 22816 52772 22880
rect 52836 22816 52852 22880
rect 52916 22816 52924 22880
rect 52604 21792 52924 22816
rect 52604 21728 52612 21792
rect 52676 21728 52692 21792
rect 52756 21728 52772 21792
rect 52836 21728 52852 21792
rect 52916 21728 52924 21792
rect 52604 20704 52924 21728
rect 52604 20640 52612 20704
rect 52676 20640 52692 20704
rect 52756 20640 52772 20704
rect 52836 20640 52852 20704
rect 52916 20640 52924 20704
rect 52604 19616 52924 20640
rect 52604 19552 52612 19616
rect 52676 19552 52692 19616
rect 52756 19552 52772 19616
rect 52836 19552 52852 19616
rect 52916 19552 52924 19616
rect 52604 18954 52924 19552
rect 52604 18718 52646 18954
rect 52882 18718 52924 18954
rect 52604 18528 52924 18718
rect 52604 18464 52612 18528
rect 52676 18464 52692 18528
rect 52756 18464 52772 18528
rect 52836 18464 52852 18528
rect 52916 18464 52924 18528
rect 52604 17440 52924 18464
rect 52604 17376 52612 17440
rect 52676 17376 52692 17440
rect 52756 17376 52772 17440
rect 52836 17376 52852 17440
rect 52916 17376 52924 17440
rect 52604 16352 52924 17376
rect 52604 16288 52612 16352
rect 52676 16288 52692 16352
rect 52756 16288 52772 16352
rect 52836 16288 52852 16352
rect 52916 16288 52924 16352
rect 52604 15264 52924 16288
rect 52604 15200 52612 15264
rect 52676 15200 52692 15264
rect 52756 15200 52772 15264
rect 52836 15200 52852 15264
rect 52916 15200 52924 15264
rect 52604 14176 52924 15200
rect 52604 14112 52612 14176
rect 52676 14112 52692 14176
rect 52756 14112 52772 14176
rect 52836 14112 52852 14176
rect 52916 14112 52924 14176
rect 52604 13954 52924 14112
rect 52604 13718 52646 13954
rect 52882 13718 52924 13954
rect 52604 13088 52924 13718
rect 52604 13024 52612 13088
rect 52676 13024 52692 13088
rect 52756 13024 52772 13088
rect 52836 13024 52852 13088
rect 52916 13024 52924 13088
rect 52604 12000 52924 13024
rect 52604 11936 52612 12000
rect 52676 11936 52692 12000
rect 52756 11936 52772 12000
rect 52836 11936 52852 12000
rect 52916 11936 52924 12000
rect 52604 10912 52924 11936
rect 52604 10848 52612 10912
rect 52676 10848 52692 10912
rect 52756 10848 52772 10912
rect 52836 10848 52852 10912
rect 52916 10848 52924 10912
rect 52604 9824 52924 10848
rect 52604 9760 52612 9824
rect 52676 9760 52692 9824
rect 52756 9760 52772 9824
rect 52836 9760 52852 9824
rect 52916 9760 52924 9824
rect 52604 8954 52924 9760
rect 52604 8736 52646 8954
rect 52882 8736 52924 8954
rect 52604 8672 52612 8736
rect 52676 8672 52692 8718
rect 52756 8672 52772 8718
rect 52836 8672 52852 8718
rect 52916 8672 52924 8736
rect 52604 7648 52924 8672
rect 52604 7584 52612 7648
rect 52676 7584 52692 7648
rect 52756 7584 52772 7648
rect 52836 7584 52852 7648
rect 52916 7584 52924 7648
rect 52604 6560 52924 7584
rect 52604 6496 52612 6560
rect 52676 6496 52692 6560
rect 52756 6496 52772 6560
rect 52836 6496 52852 6560
rect 52916 6496 52924 6560
rect 52604 5472 52924 6496
rect 52604 5408 52612 5472
rect 52676 5408 52692 5472
rect 52756 5408 52772 5472
rect 52836 5408 52852 5472
rect 52916 5408 52924 5472
rect 52604 4384 52924 5408
rect 52604 4320 52612 4384
rect 52676 4320 52692 4384
rect 52756 4320 52772 4384
rect 52836 4320 52852 4384
rect 52916 4320 52924 4384
rect 52604 3954 52924 4320
rect 52604 3718 52646 3954
rect 52882 3718 52924 3954
rect 52604 3296 52924 3718
rect 52604 3232 52612 3296
rect 52676 3232 52692 3296
rect 52756 3232 52772 3296
rect 52836 3232 52852 3296
rect 52916 3232 52924 3296
rect 52604 2208 52924 3232
rect 52604 2144 52612 2208
rect 52676 2144 52692 2208
rect 52756 2144 52772 2208
rect 52836 2144 52852 2208
rect 52916 2144 52924 2208
rect 52604 2128 52924 2144
rect 56944 57152 57264 57712
rect 56944 57088 56952 57152
rect 57016 57088 57032 57152
rect 57096 57088 57112 57152
rect 57176 57088 57192 57152
rect 57256 57088 57264 57152
rect 56944 56064 57264 57088
rect 56944 56000 56952 56064
rect 57016 56000 57032 56064
rect 57096 56000 57112 56064
rect 57176 56000 57192 56064
rect 57256 56000 57264 56064
rect 56944 54976 57264 56000
rect 56944 54912 56952 54976
rect 57016 54912 57032 54976
rect 57096 54912 57112 54976
rect 57176 54912 57192 54976
rect 57256 54912 57264 54976
rect 56944 53888 57264 54912
rect 56944 53824 56952 53888
rect 57016 53824 57032 53888
rect 57096 53824 57112 53888
rect 57176 53824 57192 53888
rect 57256 53824 57264 53888
rect 56944 53294 57264 53824
rect 56944 53058 56986 53294
rect 57222 53058 57264 53294
rect 56944 52800 57264 53058
rect 56944 52736 56952 52800
rect 57016 52736 57032 52800
rect 57096 52736 57112 52800
rect 57176 52736 57192 52800
rect 57256 52736 57264 52800
rect 56944 51712 57264 52736
rect 56944 51648 56952 51712
rect 57016 51648 57032 51712
rect 57096 51648 57112 51712
rect 57176 51648 57192 51712
rect 57256 51648 57264 51712
rect 56944 50624 57264 51648
rect 56944 50560 56952 50624
rect 57016 50560 57032 50624
rect 57096 50560 57112 50624
rect 57176 50560 57192 50624
rect 57256 50560 57264 50624
rect 56944 49536 57264 50560
rect 56944 49472 56952 49536
rect 57016 49472 57032 49536
rect 57096 49472 57112 49536
rect 57176 49472 57192 49536
rect 57256 49472 57264 49536
rect 56944 48448 57264 49472
rect 56944 48384 56952 48448
rect 57016 48384 57032 48448
rect 57096 48384 57112 48448
rect 57176 48384 57192 48448
rect 57256 48384 57264 48448
rect 56944 48294 57264 48384
rect 56944 48058 56986 48294
rect 57222 48058 57264 48294
rect 56944 47360 57264 48058
rect 56944 47296 56952 47360
rect 57016 47296 57032 47360
rect 57096 47296 57112 47360
rect 57176 47296 57192 47360
rect 57256 47296 57264 47360
rect 56944 46272 57264 47296
rect 56944 46208 56952 46272
rect 57016 46208 57032 46272
rect 57096 46208 57112 46272
rect 57176 46208 57192 46272
rect 57256 46208 57264 46272
rect 56944 45184 57264 46208
rect 56944 45120 56952 45184
rect 57016 45120 57032 45184
rect 57096 45120 57112 45184
rect 57176 45120 57192 45184
rect 57256 45120 57264 45184
rect 56944 44096 57264 45120
rect 56944 44032 56952 44096
rect 57016 44032 57032 44096
rect 57096 44032 57112 44096
rect 57176 44032 57192 44096
rect 57256 44032 57264 44096
rect 56944 43294 57264 44032
rect 56944 43058 56986 43294
rect 57222 43058 57264 43294
rect 56944 43008 57264 43058
rect 56944 42944 56952 43008
rect 57016 42944 57032 43008
rect 57096 42944 57112 43008
rect 57176 42944 57192 43008
rect 57256 42944 57264 43008
rect 56944 41920 57264 42944
rect 56944 41856 56952 41920
rect 57016 41856 57032 41920
rect 57096 41856 57112 41920
rect 57176 41856 57192 41920
rect 57256 41856 57264 41920
rect 56944 40832 57264 41856
rect 56944 40768 56952 40832
rect 57016 40768 57032 40832
rect 57096 40768 57112 40832
rect 57176 40768 57192 40832
rect 57256 40768 57264 40832
rect 56944 39744 57264 40768
rect 56944 39680 56952 39744
rect 57016 39680 57032 39744
rect 57096 39680 57112 39744
rect 57176 39680 57192 39744
rect 57256 39680 57264 39744
rect 56944 38656 57264 39680
rect 56944 38592 56952 38656
rect 57016 38592 57032 38656
rect 57096 38592 57112 38656
rect 57176 38592 57192 38656
rect 57256 38592 57264 38656
rect 56944 38294 57264 38592
rect 56944 38058 56986 38294
rect 57222 38058 57264 38294
rect 56944 37568 57264 38058
rect 56944 37504 56952 37568
rect 57016 37504 57032 37568
rect 57096 37504 57112 37568
rect 57176 37504 57192 37568
rect 57256 37504 57264 37568
rect 56944 36480 57264 37504
rect 56944 36416 56952 36480
rect 57016 36416 57032 36480
rect 57096 36416 57112 36480
rect 57176 36416 57192 36480
rect 57256 36416 57264 36480
rect 56944 35392 57264 36416
rect 56944 35328 56952 35392
rect 57016 35328 57032 35392
rect 57096 35328 57112 35392
rect 57176 35328 57192 35392
rect 57256 35328 57264 35392
rect 56944 34304 57264 35328
rect 56944 34240 56952 34304
rect 57016 34240 57032 34304
rect 57096 34240 57112 34304
rect 57176 34240 57192 34304
rect 57256 34240 57264 34304
rect 56944 33294 57264 34240
rect 56944 33216 56986 33294
rect 57222 33216 57264 33294
rect 56944 33152 56952 33216
rect 57256 33152 57264 33216
rect 56944 33058 56986 33152
rect 57222 33058 57264 33152
rect 56944 32128 57264 33058
rect 56944 32064 56952 32128
rect 57016 32064 57032 32128
rect 57096 32064 57112 32128
rect 57176 32064 57192 32128
rect 57256 32064 57264 32128
rect 56944 31040 57264 32064
rect 56944 30976 56952 31040
rect 57016 30976 57032 31040
rect 57096 30976 57112 31040
rect 57176 30976 57192 31040
rect 57256 30976 57264 31040
rect 56944 29952 57264 30976
rect 56944 29888 56952 29952
rect 57016 29888 57032 29952
rect 57096 29888 57112 29952
rect 57176 29888 57192 29952
rect 57256 29888 57264 29952
rect 56944 28864 57264 29888
rect 56944 28800 56952 28864
rect 57016 28800 57032 28864
rect 57096 28800 57112 28864
rect 57176 28800 57192 28864
rect 57256 28800 57264 28864
rect 56944 28294 57264 28800
rect 56944 28058 56986 28294
rect 57222 28058 57264 28294
rect 56944 27776 57264 28058
rect 56944 27712 56952 27776
rect 57016 27712 57032 27776
rect 57096 27712 57112 27776
rect 57176 27712 57192 27776
rect 57256 27712 57264 27776
rect 56944 26688 57264 27712
rect 56944 26624 56952 26688
rect 57016 26624 57032 26688
rect 57096 26624 57112 26688
rect 57176 26624 57192 26688
rect 57256 26624 57264 26688
rect 56944 25600 57264 26624
rect 56944 25536 56952 25600
rect 57016 25536 57032 25600
rect 57096 25536 57112 25600
rect 57176 25536 57192 25600
rect 57256 25536 57264 25600
rect 56944 24512 57264 25536
rect 56944 24448 56952 24512
rect 57016 24448 57032 24512
rect 57096 24448 57112 24512
rect 57176 24448 57192 24512
rect 57256 24448 57264 24512
rect 56944 23424 57264 24448
rect 56944 23360 56952 23424
rect 57016 23360 57032 23424
rect 57096 23360 57112 23424
rect 57176 23360 57192 23424
rect 57256 23360 57264 23424
rect 56944 23294 57264 23360
rect 56944 23058 56986 23294
rect 57222 23058 57264 23294
rect 56944 22336 57264 23058
rect 56944 22272 56952 22336
rect 57016 22272 57032 22336
rect 57096 22272 57112 22336
rect 57176 22272 57192 22336
rect 57256 22272 57264 22336
rect 56944 21248 57264 22272
rect 56944 21184 56952 21248
rect 57016 21184 57032 21248
rect 57096 21184 57112 21248
rect 57176 21184 57192 21248
rect 57256 21184 57264 21248
rect 56944 20160 57264 21184
rect 56944 20096 56952 20160
rect 57016 20096 57032 20160
rect 57096 20096 57112 20160
rect 57176 20096 57192 20160
rect 57256 20096 57264 20160
rect 56944 19072 57264 20096
rect 56944 19008 56952 19072
rect 57016 19008 57032 19072
rect 57096 19008 57112 19072
rect 57176 19008 57192 19072
rect 57256 19008 57264 19072
rect 56944 18294 57264 19008
rect 56944 18058 56986 18294
rect 57222 18058 57264 18294
rect 56944 17984 57264 18058
rect 56944 17920 56952 17984
rect 57016 17920 57032 17984
rect 57096 17920 57112 17984
rect 57176 17920 57192 17984
rect 57256 17920 57264 17984
rect 56944 16896 57264 17920
rect 56944 16832 56952 16896
rect 57016 16832 57032 16896
rect 57096 16832 57112 16896
rect 57176 16832 57192 16896
rect 57256 16832 57264 16896
rect 56944 15808 57264 16832
rect 56944 15744 56952 15808
rect 57016 15744 57032 15808
rect 57096 15744 57112 15808
rect 57176 15744 57192 15808
rect 57256 15744 57264 15808
rect 56944 14720 57264 15744
rect 56944 14656 56952 14720
rect 57016 14656 57032 14720
rect 57096 14656 57112 14720
rect 57176 14656 57192 14720
rect 57256 14656 57264 14720
rect 56944 13632 57264 14656
rect 56944 13568 56952 13632
rect 57016 13568 57032 13632
rect 57096 13568 57112 13632
rect 57176 13568 57192 13632
rect 57256 13568 57264 13632
rect 56944 13294 57264 13568
rect 56944 13058 56986 13294
rect 57222 13058 57264 13294
rect 56944 12544 57264 13058
rect 56944 12480 56952 12544
rect 57016 12480 57032 12544
rect 57096 12480 57112 12544
rect 57176 12480 57192 12544
rect 57256 12480 57264 12544
rect 56944 11456 57264 12480
rect 56944 11392 56952 11456
rect 57016 11392 57032 11456
rect 57096 11392 57112 11456
rect 57176 11392 57192 11456
rect 57256 11392 57264 11456
rect 56944 10368 57264 11392
rect 56944 10304 56952 10368
rect 57016 10304 57032 10368
rect 57096 10304 57112 10368
rect 57176 10304 57192 10368
rect 57256 10304 57264 10368
rect 56944 9280 57264 10304
rect 56944 9216 56952 9280
rect 57016 9216 57032 9280
rect 57096 9216 57112 9280
rect 57176 9216 57192 9280
rect 57256 9216 57264 9280
rect 56944 8294 57264 9216
rect 56944 8192 56986 8294
rect 57222 8192 57264 8294
rect 56944 8128 56952 8192
rect 57256 8128 57264 8192
rect 56944 8058 56986 8128
rect 57222 8058 57264 8128
rect 56944 7104 57264 8058
rect 56944 7040 56952 7104
rect 57016 7040 57032 7104
rect 57096 7040 57112 7104
rect 57176 7040 57192 7104
rect 57256 7040 57264 7104
rect 56944 6016 57264 7040
rect 56944 5952 56952 6016
rect 57016 5952 57032 6016
rect 57096 5952 57112 6016
rect 57176 5952 57192 6016
rect 57256 5952 57264 6016
rect 56944 4928 57264 5952
rect 56944 4864 56952 4928
rect 57016 4864 57032 4928
rect 57096 4864 57112 4928
rect 57176 4864 57192 4928
rect 57256 4864 57264 4928
rect 56944 3840 57264 4864
rect 56944 3776 56952 3840
rect 57016 3776 57032 3840
rect 57096 3776 57112 3840
rect 57176 3776 57192 3840
rect 57256 3776 57264 3840
rect 56944 3294 57264 3776
rect 56944 3058 56986 3294
rect 57222 3058 57264 3294
rect 56944 2752 57264 3058
rect 56944 2688 56952 2752
rect 57016 2688 57032 2752
rect 57096 2688 57112 2752
rect 57176 2688 57192 2752
rect 57256 2688 57264 2752
rect 56944 2128 57264 2688
rect 57604 57696 57924 57712
rect 57604 57632 57612 57696
rect 57676 57632 57692 57696
rect 57756 57632 57772 57696
rect 57836 57632 57852 57696
rect 57916 57632 57924 57696
rect 57604 56608 57924 57632
rect 57604 56544 57612 56608
rect 57676 56544 57692 56608
rect 57756 56544 57772 56608
rect 57836 56544 57852 56608
rect 57916 56544 57924 56608
rect 57604 55520 57924 56544
rect 57604 55456 57612 55520
rect 57676 55456 57692 55520
rect 57756 55456 57772 55520
rect 57836 55456 57852 55520
rect 57916 55456 57924 55520
rect 57604 54432 57924 55456
rect 57604 54368 57612 54432
rect 57676 54368 57692 54432
rect 57756 54368 57772 54432
rect 57836 54368 57852 54432
rect 57916 54368 57924 54432
rect 57604 53954 57924 54368
rect 57604 53718 57646 53954
rect 57882 53718 57924 53954
rect 57604 53344 57924 53718
rect 57604 53280 57612 53344
rect 57676 53280 57692 53344
rect 57756 53280 57772 53344
rect 57836 53280 57852 53344
rect 57916 53280 57924 53344
rect 57604 52256 57924 53280
rect 57604 52192 57612 52256
rect 57676 52192 57692 52256
rect 57756 52192 57772 52256
rect 57836 52192 57852 52256
rect 57916 52192 57924 52256
rect 57604 51168 57924 52192
rect 57604 51104 57612 51168
rect 57676 51104 57692 51168
rect 57756 51104 57772 51168
rect 57836 51104 57852 51168
rect 57916 51104 57924 51168
rect 57604 50080 57924 51104
rect 57604 50016 57612 50080
rect 57676 50016 57692 50080
rect 57756 50016 57772 50080
rect 57836 50016 57852 50080
rect 57916 50016 57924 50080
rect 57604 48992 57924 50016
rect 57604 48928 57612 48992
rect 57676 48954 57692 48992
rect 57756 48954 57772 48992
rect 57836 48954 57852 48992
rect 57916 48928 57924 48992
rect 57604 48718 57646 48928
rect 57882 48718 57924 48928
rect 57604 47904 57924 48718
rect 57604 47840 57612 47904
rect 57676 47840 57692 47904
rect 57756 47840 57772 47904
rect 57836 47840 57852 47904
rect 57916 47840 57924 47904
rect 57604 46816 57924 47840
rect 57604 46752 57612 46816
rect 57676 46752 57692 46816
rect 57756 46752 57772 46816
rect 57836 46752 57852 46816
rect 57916 46752 57924 46816
rect 57604 45728 57924 46752
rect 57604 45664 57612 45728
rect 57676 45664 57692 45728
rect 57756 45664 57772 45728
rect 57836 45664 57852 45728
rect 57916 45664 57924 45728
rect 57604 44640 57924 45664
rect 57604 44576 57612 44640
rect 57676 44576 57692 44640
rect 57756 44576 57772 44640
rect 57836 44576 57852 44640
rect 57916 44576 57924 44640
rect 57604 43954 57924 44576
rect 57604 43718 57646 43954
rect 57882 43718 57924 43954
rect 57604 43552 57924 43718
rect 57604 43488 57612 43552
rect 57676 43488 57692 43552
rect 57756 43488 57772 43552
rect 57836 43488 57852 43552
rect 57916 43488 57924 43552
rect 57604 42464 57924 43488
rect 57604 42400 57612 42464
rect 57676 42400 57692 42464
rect 57756 42400 57772 42464
rect 57836 42400 57852 42464
rect 57916 42400 57924 42464
rect 57604 41376 57924 42400
rect 57604 41312 57612 41376
rect 57676 41312 57692 41376
rect 57756 41312 57772 41376
rect 57836 41312 57852 41376
rect 57916 41312 57924 41376
rect 57604 40288 57924 41312
rect 57604 40224 57612 40288
rect 57676 40224 57692 40288
rect 57756 40224 57772 40288
rect 57836 40224 57852 40288
rect 57916 40224 57924 40288
rect 57604 39200 57924 40224
rect 57604 39136 57612 39200
rect 57676 39136 57692 39200
rect 57756 39136 57772 39200
rect 57836 39136 57852 39200
rect 57916 39136 57924 39200
rect 57604 38954 57924 39136
rect 57604 38718 57646 38954
rect 57882 38718 57924 38954
rect 57604 38112 57924 38718
rect 57604 38048 57612 38112
rect 57676 38048 57692 38112
rect 57756 38048 57772 38112
rect 57836 38048 57852 38112
rect 57916 38048 57924 38112
rect 57604 37024 57924 38048
rect 57604 36960 57612 37024
rect 57676 36960 57692 37024
rect 57756 36960 57772 37024
rect 57836 36960 57852 37024
rect 57916 36960 57924 37024
rect 57604 35936 57924 36960
rect 57604 35872 57612 35936
rect 57676 35872 57692 35936
rect 57756 35872 57772 35936
rect 57836 35872 57852 35936
rect 57916 35872 57924 35936
rect 57604 34848 57924 35872
rect 57604 34784 57612 34848
rect 57676 34784 57692 34848
rect 57756 34784 57772 34848
rect 57836 34784 57852 34848
rect 57916 34784 57924 34848
rect 57604 33954 57924 34784
rect 57604 33760 57646 33954
rect 57882 33760 57924 33954
rect 57604 33696 57612 33760
rect 57676 33696 57692 33718
rect 57756 33696 57772 33718
rect 57836 33696 57852 33718
rect 57916 33696 57924 33760
rect 57604 32672 57924 33696
rect 57604 32608 57612 32672
rect 57676 32608 57692 32672
rect 57756 32608 57772 32672
rect 57836 32608 57852 32672
rect 57916 32608 57924 32672
rect 57604 31584 57924 32608
rect 57604 31520 57612 31584
rect 57676 31520 57692 31584
rect 57756 31520 57772 31584
rect 57836 31520 57852 31584
rect 57916 31520 57924 31584
rect 57604 30496 57924 31520
rect 57604 30432 57612 30496
rect 57676 30432 57692 30496
rect 57756 30432 57772 30496
rect 57836 30432 57852 30496
rect 57916 30432 57924 30496
rect 57604 29408 57924 30432
rect 57604 29344 57612 29408
rect 57676 29344 57692 29408
rect 57756 29344 57772 29408
rect 57836 29344 57852 29408
rect 57916 29344 57924 29408
rect 57604 28954 57924 29344
rect 57604 28718 57646 28954
rect 57882 28718 57924 28954
rect 57604 28320 57924 28718
rect 57604 28256 57612 28320
rect 57676 28256 57692 28320
rect 57756 28256 57772 28320
rect 57836 28256 57852 28320
rect 57916 28256 57924 28320
rect 57604 27232 57924 28256
rect 57604 27168 57612 27232
rect 57676 27168 57692 27232
rect 57756 27168 57772 27232
rect 57836 27168 57852 27232
rect 57916 27168 57924 27232
rect 57604 26144 57924 27168
rect 57604 26080 57612 26144
rect 57676 26080 57692 26144
rect 57756 26080 57772 26144
rect 57836 26080 57852 26144
rect 57916 26080 57924 26144
rect 57604 25056 57924 26080
rect 57604 24992 57612 25056
rect 57676 24992 57692 25056
rect 57756 24992 57772 25056
rect 57836 24992 57852 25056
rect 57916 24992 57924 25056
rect 57604 23968 57924 24992
rect 57604 23904 57612 23968
rect 57676 23954 57692 23968
rect 57756 23954 57772 23968
rect 57836 23954 57852 23968
rect 57916 23904 57924 23968
rect 57604 23718 57646 23904
rect 57882 23718 57924 23904
rect 57604 22880 57924 23718
rect 57604 22816 57612 22880
rect 57676 22816 57692 22880
rect 57756 22816 57772 22880
rect 57836 22816 57852 22880
rect 57916 22816 57924 22880
rect 57604 21792 57924 22816
rect 57604 21728 57612 21792
rect 57676 21728 57692 21792
rect 57756 21728 57772 21792
rect 57836 21728 57852 21792
rect 57916 21728 57924 21792
rect 57604 20704 57924 21728
rect 57604 20640 57612 20704
rect 57676 20640 57692 20704
rect 57756 20640 57772 20704
rect 57836 20640 57852 20704
rect 57916 20640 57924 20704
rect 57604 19616 57924 20640
rect 57604 19552 57612 19616
rect 57676 19552 57692 19616
rect 57756 19552 57772 19616
rect 57836 19552 57852 19616
rect 57916 19552 57924 19616
rect 57604 18954 57924 19552
rect 57604 18718 57646 18954
rect 57882 18718 57924 18954
rect 57604 18528 57924 18718
rect 57604 18464 57612 18528
rect 57676 18464 57692 18528
rect 57756 18464 57772 18528
rect 57836 18464 57852 18528
rect 57916 18464 57924 18528
rect 57604 17440 57924 18464
rect 57604 17376 57612 17440
rect 57676 17376 57692 17440
rect 57756 17376 57772 17440
rect 57836 17376 57852 17440
rect 57916 17376 57924 17440
rect 57604 16352 57924 17376
rect 57604 16288 57612 16352
rect 57676 16288 57692 16352
rect 57756 16288 57772 16352
rect 57836 16288 57852 16352
rect 57916 16288 57924 16352
rect 57604 15264 57924 16288
rect 57604 15200 57612 15264
rect 57676 15200 57692 15264
rect 57756 15200 57772 15264
rect 57836 15200 57852 15264
rect 57916 15200 57924 15264
rect 57604 14176 57924 15200
rect 57604 14112 57612 14176
rect 57676 14112 57692 14176
rect 57756 14112 57772 14176
rect 57836 14112 57852 14176
rect 57916 14112 57924 14176
rect 57604 13954 57924 14112
rect 57604 13718 57646 13954
rect 57882 13718 57924 13954
rect 57604 13088 57924 13718
rect 57604 13024 57612 13088
rect 57676 13024 57692 13088
rect 57756 13024 57772 13088
rect 57836 13024 57852 13088
rect 57916 13024 57924 13088
rect 57604 12000 57924 13024
rect 57604 11936 57612 12000
rect 57676 11936 57692 12000
rect 57756 11936 57772 12000
rect 57836 11936 57852 12000
rect 57916 11936 57924 12000
rect 57604 10912 57924 11936
rect 57604 10848 57612 10912
rect 57676 10848 57692 10912
rect 57756 10848 57772 10912
rect 57836 10848 57852 10912
rect 57916 10848 57924 10912
rect 57604 9824 57924 10848
rect 57604 9760 57612 9824
rect 57676 9760 57692 9824
rect 57756 9760 57772 9824
rect 57836 9760 57852 9824
rect 57916 9760 57924 9824
rect 57604 8954 57924 9760
rect 57604 8736 57646 8954
rect 57882 8736 57924 8954
rect 57604 8672 57612 8736
rect 57676 8672 57692 8718
rect 57756 8672 57772 8718
rect 57836 8672 57852 8718
rect 57916 8672 57924 8736
rect 57604 7648 57924 8672
rect 57604 7584 57612 7648
rect 57676 7584 57692 7648
rect 57756 7584 57772 7648
rect 57836 7584 57852 7648
rect 57916 7584 57924 7648
rect 57604 6560 57924 7584
rect 57604 6496 57612 6560
rect 57676 6496 57692 6560
rect 57756 6496 57772 6560
rect 57836 6496 57852 6560
rect 57916 6496 57924 6560
rect 57604 5472 57924 6496
rect 57604 5408 57612 5472
rect 57676 5408 57692 5472
rect 57756 5408 57772 5472
rect 57836 5408 57852 5472
rect 57916 5408 57924 5472
rect 57604 4384 57924 5408
rect 57604 4320 57612 4384
rect 57676 4320 57692 4384
rect 57756 4320 57772 4384
rect 57836 4320 57852 4384
rect 57916 4320 57924 4384
rect 57604 3954 57924 4320
rect 57604 3718 57646 3954
rect 57882 3718 57924 3954
rect 57604 3296 57924 3718
rect 57604 3232 57612 3296
rect 57676 3232 57692 3296
rect 57756 3232 57772 3296
rect 57836 3232 57852 3296
rect 57916 3232 57924 3296
rect 57604 2208 57924 3232
rect 57604 2144 57612 2208
rect 57676 2144 57692 2208
rect 57756 2144 57772 2208
rect 57836 2144 57852 2208
rect 57916 2144 57924 2208
rect 57604 2128 57924 2144
<< via4 >>
rect 1986 53058 2222 53294
rect 1986 48058 2222 48294
rect 1986 43058 2222 43294
rect 1986 38058 2222 38294
rect 1986 33216 2222 33294
rect 1986 33152 2016 33216
rect 2016 33152 2032 33216
rect 2032 33152 2096 33216
rect 2096 33152 2112 33216
rect 2112 33152 2176 33216
rect 2176 33152 2192 33216
rect 2192 33152 2222 33216
rect 1986 33058 2222 33152
rect 1986 28058 2222 28294
rect 1986 23058 2222 23294
rect 1986 18058 2222 18294
rect 1986 13058 2222 13294
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1986 3058 2222 3294
rect 2646 53718 2882 53954
rect 2646 48928 2676 48954
rect 2676 48928 2692 48954
rect 2692 48928 2756 48954
rect 2756 48928 2772 48954
rect 2772 48928 2836 48954
rect 2836 48928 2852 48954
rect 2852 48928 2882 48954
rect 2646 48718 2882 48928
rect 2646 43718 2882 43954
rect 2646 38718 2882 38954
rect 2646 33760 2882 33954
rect 2646 33718 2676 33760
rect 2676 33718 2692 33760
rect 2692 33718 2756 33760
rect 2756 33718 2772 33760
rect 2772 33718 2836 33760
rect 2836 33718 2852 33760
rect 2852 33718 2882 33760
rect 2646 28718 2882 28954
rect 2646 23904 2676 23954
rect 2676 23904 2692 23954
rect 2692 23904 2756 23954
rect 2756 23904 2772 23954
rect 2772 23904 2836 23954
rect 2836 23904 2852 23954
rect 2852 23904 2882 23954
rect 2646 23718 2882 23904
rect 2646 18718 2882 18954
rect 2646 13718 2882 13954
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 2646 3718 2882 3954
rect 6986 53058 7222 53294
rect 6986 48058 7222 48294
rect 6986 43058 7222 43294
rect 6986 38058 7222 38294
rect 6986 33216 7222 33294
rect 6986 33152 7016 33216
rect 7016 33152 7032 33216
rect 7032 33152 7096 33216
rect 7096 33152 7112 33216
rect 7112 33152 7176 33216
rect 7176 33152 7192 33216
rect 7192 33152 7222 33216
rect 6986 33058 7222 33152
rect 6986 28058 7222 28294
rect 6986 23058 7222 23294
rect 6986 18058 7222 18294
rect 6986 13058 7222 13294
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 6986 3058 7222 3294
rect 7646 53718 7882 53954
rect 7646 48928 7676 48954
rect 7676 48928 7692 48954
rect 7692 48928 7756 48954
rect 7756 48928 7772 48954
rect 7772 48928 7836 48954
rect 7836 48928 7852 48954
rect 7852 48928 7882 48954
rect 7646 48718 7882 48928
rect 7646 43718 7882 43954
rect 7646 38718 7882 38954
rect 7646 33760 7882 33954
rect 7646 33718 7676 33760
rect 7676 33718 7692 33760
rect 7692 33718 7756 33760
rect 7756 33718 7772 33760
rect 7772 33718 7836 33760
rect 7836 33718 7852 33760
rect 7852 33718 7882 33760
rect 7646 28718 7882 28954
rect 7646 23904 7676 23954
rect 7676 23904 7692 23954
rect 7692 23904 7756 23954
rect 7756 23904 7772 23954
rect 7772 23904 7836 23954
rect 7836 23904 7852 23954
rect 7852 23904 7882 23954
rect 7646 23718 7882 23904
rect 7646 18718 7882 18954
rect 7646 13718 7882 13954
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 7646 3718 7882 3954
rect 11986 53058 12222 53294
rect 11986 48058 12222 48294
rect 11986 43058 12222 43294
rect 11986 38058 12222 38294
rect 11986 33216 12222 33294
rect 11986 33152 12016 33216
rect 12016 33152 12032 33216
rect 12032 33152 12096 33216
rect 12096 33152 12112 33216
rect 12112 33152 12176 33216
rect 12176 33152 12192 33216
rect 12192 33152 12222 33216
rect 11986 33058 12222 33152
rect 11986 28058 12222 28294
rect 11986 23058 12222 23294
rect 11986 18058 12222 18294
rect 11986 13058 12222 13294
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 11986 3058 12222 3294
rect 12646 53718 12882 53954
rect 12646 48928 12676 48954
rect 12676 48928 12692 48954
rect 12692 48928 12756 48954
rect 12756 48928 12772 48954
rect 12772 48928 12836 48954
rect 12836 48928 12852 48954
rect 12852 48928 12882 48954
rect 12646 48718 12882 48928
rect 12646 43718 12882 43954
rect 12646 38718 12882 38954
rect 12646 33760 12882 33954
rect 12646 33718 12676 33760
rect 12676 33718 12692 33760
rect 12692 33718 12756 33760
rect 12756 33718 12772 33760
rect 12772 33718 12836 33760
rect 12836 33718 12852 33760
rect 12852 33718 12882 33760
rect 12646 28718 12882 28954
rect 12646 23904 12676 23954
rect 12676 23904 12692 23954
rect 12692 23904 12756 23954
rect 12756 23904 12772 23954
rect 12772 23904 12836 23954
rect 12836 23904 12852 23954
rect 12852 23904 12882 23954
rect 12646 23718 12882 23904
rect 12646 18718 12882 18954
rect 12646 13718 12882 13954
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 12646 3718 12882 3954
rect 16986 53058 17222 53294
rect 16986 48058 17222 48294
rect 16986 43058 17222 43294
rect 16986 38058 17222 38294
rect 16986 33216 17222 33294
rect 16986 33152 17016 33216
rect 17016 33152 17032 33216
rect 17032 33152 17096 33216
rect 17096 33152 17112 33216
rect 17112 33152 17176 33216
rect 17176 33152 17192 33216
rect 17192 33152 17222 33216
rect 16986 33058 17222 33152
rect 16986 28058 17222 28294
rect 16986 23058 17222 23294
rect 16986 18058 17222 18294
rect 16986 13058 17222 13294
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 16986 3058 17222 3294
rect 17646 53718 17882 53954
rect 17646 48928 17676 48954
rect 17676 48928 17692 48954
rect 17692 48928 17756 48954
rect 17756 48928 17772 48954
rect 17772 48928 17836 48954
rect 17836 48928 17852 48954
rect 17852 48928 17882 48954
rect 17646 48718 17882 48928
rect 17646 43718 17882 43954
rect 17646 38718 17882 38954
rect 17646 33760 17882 33954
rect 17646 33718 17676 33760
rect 17676 33718 17692 33760
rect 17692 33718 17756 33760
rect 17756 33718 17772 33760
rect 17772 33718 17836 33760
rect 17836 33718 17852 33760
rect 17852 33718 17882 33760
rect 17646 28718 17882 28954
rect 17646 23904 17676 23954
rect 17676 23904 17692 23954
rect 17692 23904 17756 23954
rect 17756 23904 17772 23954
rect 17772 23904 17836 23954
rect 17836 23904 17852 23954
rect 17852 23904 17882 23954
rect 17646 23718 17882 23904
rect 17646 18718 17882 18954
rect 17646 13718 17882 13954
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 17646 3718 17882 3954
rect 21986 53058 22222 53294
rect 21986 48058 22222 48294
rect 21986 43058 22222 43294
rect 21986 38058 22222 38294
rect 21986 33216 22222 33294
rect 21986 33152 22016 33216
rect 22016 33152 22032 33216
rect 22032 33152 22096 33216
rect 22096 33152 22112 33216
rect 22112 33152 22176 33216
rect 22176 33152 22192 33216
rect 22192 33152 22222 33216
rect 21986 33058 22222 33152
rect 21986 28058 22222 28294
rect 21986 23058 22222 23294
rect 21986 18058 22222 18294
rect 21986 13058 22222 13294
rect 21986 8192 22222 8294
rect 21986 8128 22016 8192
rect 22016 8128 22032 8192
rect 22032 8128 22096 8192
rect 22096 8128 22112 8192
rect 22112 8128 22176 8192
rect 22176 8128 22192 8192
rect 22192 8128 22222 8192
rect 21986 8058 22222 8128
rect 21986 3058 22222 3294
rect 22646 53718 22882 53954
rect 22646 48928 22676 48954
rect 22676 48928 22692 48954
rect 22692 48928 22756 48954
rect 22756 48928 22772 48954
rect 22772 48928 22836 48954
rect 22836 48928 22852 48954
rect 22852 48928 22882 48954
rect 22646 48718 22882 48928
rect 22646 43718 22882 43954
rect 22646 38718 22882 38954
rect 22646 33760 22882 33954
rect 22646 33718 22676 33760
rect 22676 33718 22692 33760
rect 22692 33718 22756 33760
rect 22756 33718 22772 33760
rect 22772 33718 22836 33760
rect 22836 33718 22852 33760
rect 22852 33718 22882 33760
rect 22646 28718 22882 28954
rect 22646 23904 22676 23954
rect 22676 23904 22692 23954
rect 22692 23904 22756 23954
rect 22756 23904 22772 23954
rect 22772 23904 22836 23954
rect 22836 23904 22852 23954
rect 22852 23904 22882 23954
rect 22646 23718 22882 23904
rect 22646 18718 22882 18954
rect 22646 13718 22882 13954
rect 22646 8736 22882 8954
rect 22646 8718 22676 8736
rect 22676 8718 22692 8736
rect 22692 8718 22756 8736
rect 22756 8718 22772 8736
rect 22772 8718 22836 8736
rect 22836 8718 22852 8736
rect 22852 8718 22882 8736
rect 22646 3718 22882 3954
rect 26986 53058 27222 53294
rect 26986 48058 27222 48294
rect 26986 43058 27222 43294
rect 26986 38058 27222 38294
rect 26986 33216 27222 33294
rect 26986 33152 27016 33216
rect 27016 33152 27032 33216
rect 27032 33152 27096 33216
rect 27096 33152 27112 33216
rect 27112 33152 27176 33216
rect 27176 33152 27192 33216
rect 27192 33152 27222 33216
rect 26986 33058 27222 33152
rect 26986 28058 27222 28294
rect 26986 23058 27222 23294
rect 26986 18058 27222 18294
rect 26986 13058 27222 13294
rect 26986 8192 27222 8294
rect 26986 8128 27016 8192
rect 27016 8128 27032 8192
rect 27032 8128 27096 8192
rect 27096 8128 27112 8192
rect 27112 8128 27176 8192
rect 27176 8128 27192 8192
rect 27192 8128 27222 8192
rect 26986 8058 27222 8128
rect 26986 3058 27222 3294
rect 27646 53718 27882 53954
rect 27646 48928 27676 48954
rect 27676 48928 27692 48954
rect 27692 48928 27756 48954
rect 27756 48928 27772 48954
rect 27772 48928 27836 48954
rect 27836 48928 27852 48954
rect 27852 48928 27882 48954
rect 27646 48718 27882 48928
rect 27646 43718 27882 43954
rect 27646 38718 27882 38954
rect 27646 33760 27882 33954
rect 27646 33718 27676 33760
rect 27676 33718 27692 33760
rect 27692 33718 27756 33760
rect 27756 33718 27772 33760
rect 27772 33718 27836 33760
rect 27836 33718 27852 33760
rect 27852 33718 27882 33760
rect 27646 28718 27882 28954
rect 27646 23904 27676 23954
rect 27676 23904 27692 23954
rect 27692 23904 27756 23954
rect 27756 23904 27772 23954
rect 27772 23904 27836 23954
rect 27836 23904 27852 23954
rect 27852 23904 27882 23954
rect 27646 23718 27882 23904
rect 27646 18718 27882 18954
rect 27646 13718 27882 13954
rect 27646 8736 27882 8954
rect 27646 8718 27676 8736
rect 27676 8718 27692 8736
rect 27692 8718 27756 8736
rect 27756 8718 27772 8736
rect 27772 8718 27836 8736
rect 27836 8718 27852 8736
rect 27852 8718 27882 8736
rect 27646 3718 27882 3954
rect 31986 53058 32222 53294
rect 31986 48058 32222 48294
rect 31986 43058 32222 43294
rect 31986 38058 32222 38294
rect 31986 33216 32222 33294
rect 31986 33152 32016 33216
rect 32016 33152 32032 33216
rect 32032 33152 32096 33216
rect 32096 33152 32112 33216
rect 32112 33152 32176 33216
rect 32176 33152 32192 33216
rect 32192 33152 32222 33216
rect 31986 33058 32222 33152
rect 31986 28058 32222 28294
rect 31986 23058 32222 23294
rect 31986 18058 32222 18294
rect 31986 13058 32222 13294
rect 31986 8192 32222 8294
rect 31986 8128 32016 8192
rect 32016 8128 32032 8192
rect 32032 8128 32096 8192
rect 32096 8128 32112 8192
rect 32112 8128 32176 8192
rect 32176 8128 32192 8192
rect 32192 8128 32222 8192
rect 31986 8058 32222 8128
rect 31986 3058 32222 3294
rect 32646 53718 32882 53954
rect 32646 48928 32676 48954
rect 32676 48928 32692 48954
rect 32692 48928 32756 48954
rect 32756 48928 32772 48954
rect 32772 48928 32836 48954
rect 32836 48928 32852 48954
rect 32852 48928 32882 48954
rect 32646 48718 32882 48928
rect 32646 43718 32882 43954
rect 32646 38718 32882 38954
rect 32646 33760 32882 33954
rect 32646 33718 32676 33760
rect 32676 33718 32692 33760
rect 32692 33718 32756 33760
rect 32756 33718 32772 33760
rect 32772 33718 32836 33760
rect 32836 33718 32852 33760
rect 32852 33718 32882 33760
rect 32646 28718 32882 28954
rect 32646 23904 32676 23954
rect 32676 23904 32692 23954
rect 32692 23904 32756 23954
rect 32756 23904 32772 23954
rect 32772 23904 32836 23954
rect 32836 23904 32852 23954
rect 32852 23904 32882 23954
rect 32646 23718 32882 23904
rect 32646 18718 32882 18954
rect 32646 13718 32882 13954
rect 32646 8736 32882 8954
rect 32646 8718 32676 8736
rect 32676 8718 32692 8736
rect 32692 8718 32756 8736
rect 32756 8718 32772 8736
rect 32772 8718 32836 8736
rect 32836 8718 32852 8736
rect 32852 8718 32882 8736
rect 32646 3718 32882 3954
rect 36986 53058 37222 53294
rect 36986 48058 37222 48294
rect 36986 43058 37222 43294
rect 36986 38058 37222 38294
rect 36986 33216 37222 33294
rect 36986 33152 37016 33216
rect 37016 33152 37032 33216
rect 37032 33152 37096 33216
rect 37096 33152 37112 33216
rect 37112 33152 37176 33216
rect 37176 33152 37192 33216
rect 37192 33152 37222 33216
rect 36986 33058 37222 33152
rect 36986 28058 37222 28294
rect 36986 23058 37222 23294
rect 36986 18058 37222 18294
rect 36986 13058 37222 13294
rect 36986 8192 37222 8294
rect 36986 8128 37016 8192
rect 37016 8128 37032 8192
rect 37032 8128 37096 8192
rect 37096 8128 37112 8192
rect 37112 8128 37176 8192
rect 37176 8128 37192 8192
rect 37192 8128 37222 8192
rect 36986 8058 37222 8128
rect 36986 3058 37222 3294
rect 37646 53718 37882 53954
rect 37646 48928 37676 48954
rect 37676 48928 37692 48954
rect 37692 48928 37756 48954
rect 37756 48928 37772 48954
rect 37772 48928 37836 48954
rect 37836 48928 37852 48954
rect 37852 48928 37882 48954
rect 37646 48718 37882 48928
rect 37646 43718 37882 43954
rect 37646 38718 37882 38954
rect 37646 33760 37882 33954
rect 37646 33718 37676 33760
rect 37676 33718 37692 33760
rect 37692 33718 37756 33760
rect 37756 33718 37772 33760
rect 37772 33718 37836 33760
rect 37836 33718 37852 33760
rect 37852 33718 37882 33760
rect 37646 28718 37882 28954
rect 37646 23904 37676 23954
rect 37676 23904 37692 23954
rect 37692 23904 37756 23954
rect 37756 23904 37772 23954
rect 37772 23904 37836 23954
rect 37836 23904 37852 23954
rect 37852 23904 37882 23954
rect 37646 23718 37882 23904
rect 37646 18718 37882 18954
rect 37646 13718 37882 13954
rect 37646 8736 37882 8954
rect 37646 8718 37676 8736
rect 37676 8718 37692 8736
rect 37692 8718 37756 8736
rect 37756 8718 37772 8736
rect 37772 8718 37836 8736
rect 37836 8718 37852 8736
rect 37852 8718 37882 8736
rect 37646 3718 37882 3954
rect 41986 53058 42222 53294
rect 41986 48058 42222 48294
rect 41986 43058 42222 43294
rect 41986 38058 42222 38294
rect 41986 33216 42222 33294
rect 41986 33152 42016 33216
rect 42016 33152 42032 33216
rect 42032 33152 42096 33216
rect 42096 33152 42112 33216
rect 42112 33152 42176 33216
rect 42176 33152 42192 33216
rect 42192 33152 42222 33216
rect 41986 33058 42222 33152
rect 41986 28058 42222 28294
rect 41986 23058 42222 23294
rect 41986 18058 42222 18294
rect 41986 13058 42222 13294
rect 41986 8192 42222 8294
rect 41986 8128 42016 8192
rect 42016 8128 42032 8192
rect 42032 8128 42096 8192
rect 42096 8128 42112 8192
rect 42112 8128 42176 8192
rect 42176 8128 42192 8192
rect 42192 8128 42222 8192
rect 41986 8058 42222 8128
rect 41986 3058 42222 3294
rect 42646 53718 42882 53954
rect 42646 48928 42676 48954
rect 42676 48928 42692 48954
rect 42692 48928 42756 48954
rect 42756 48928 42772 48954
rect 42772 48928 42836 48954
rect 42836 48928 42852 48954
rect 42852 48928 42882 48954
rect 42646 48718 42882 48928
rect 42646 43718 42882 43954
rect 42646 38718 42882 38954
rect 42646 33760 42882 33954
rect 42646 33718 42676 33760
rect 42676 33718 42692 33760
rect 42692 33718 42756 33760
rect 42756 33718 42772 33760
rect 42772 33718 42836 33760
rect 42836 33718 42852 33760
rect 42852 33718 42882 33760
rect 42646 28718 42882 28954
rect 42646 23904 42676 23954
rect 42676 23904 42692 23954
rect 42692 23904 42756 23954
rect 42756 23904 42772 23954
rect 42772 23904 42836 23954
rect 42836 23904 42852 23954
rect 42852 23904 42882 23954
rect 42646 23718 42882 23904
rect 42646 18718 42882 18954
rect 42646 13718 42882 13954
rect 42646 8736 42882 8954
rect 42646 8718 42676 8736
rect 42676 8718 42692 8736
rect 42692 8718 42756 8736
rect 42756 8718 42772 8736
rect 42772 8718 42836 8736
rect 42836 8718 42852 8736
rect 42852 8718 42882 8736
rect 42646 3718 42882 3954
rect 46986 53058 47222 53294
rect 46986 48058 47222 48294
rect 46986 43058 47222 43294
rect 46986 38058 47222 38294
rect 46986 33216 47222 33294
rect 46986 33152 47016 33216
rect 47016 33152 47032 33216
rect 47032 33152 47096 33216
rect 47096 33152 47112 33216
rect 47112 33152 47176 33216
rect 47176 33152 47192 33216
rect 47192 33152 47222 33216
rect 46986 33058 47222 33152
rect 46986 28058 47222 28294
rect 46986 23058 47222 23294
rect 46986 18058 47222 18294
rect 46986 13058 47222 13294
rect 46986 8192 47222 8294
rect 46986 8128 47016 8192
rect 47016 8128 47032 8192
rect 47032 8128 47096 8192
rect 47096 8128 47112 8192
rect 47112 8128 47176 8192
rect 47176 8128 47192 8192
rect 47192 8128 47222 8192
rect 46986 8058 47222 8128
rect 46986 3058 47222 3294
rect 47646 53718 47882 53954
rect 47646 48928 47676 48954
rect 47676 48928 47692 48954
rect 47692 48928 47756 48954
rect 47756 48928 47772 48954
rect 47772 48928 47836 48954
rect 47836 48928 47852 48954
rect 47852 48928 47882 48954
rect 47646 48718 47882 48928
rect 47646 43718 47882 43954
rect 47646 38718 47882 38954
rect 47646 33760 47882 33954
rect 47646 33718 47676 33760
rect 47676 33718 47692 33760
rect 47692 33718 47756 33760
rect 47756 33718 47772 33760
rect 47772 33718 47836 33760
rect 47836 33718 47852 33760
rect 47852 33718 47882 33760
rect 47646 28718 47882 28954
rect 47646 23904 47676 23954
rect 47676 23904 47692 23954
rect 47692 23904 47756 23954
rect 47756 23904 47772 23954
rect 47772 23904 47836 23954
rect 47836 23904 47852 23954
rect 47852 23904 47882 23954
rect 47646 23718 47882 23904
rect 47646 18718 47882 18954
rect 47646 13718 47882 13954
rect 47646 8736 47882 8954
rect 47646 8718 47676 8736
rect 47676 8718 47692 8736
rect 47692 8718 47756 8736
rect 47756 8718 47772 8736
rect 47772 8718 47836 8736
rect 47836 8718 47852 8736
rect 47852 8718 47882 8736
rect 47646 3718 47882 3954
rect 51986 53058 52222 53294
rect 51986 48058 52222 48294
rect 51986 43058 52222 43294
rect 51986 38058 52222 38294
rect 51986 33216 52222 33294
rect 51986 33152 52016 33216
rect 52016 33152 52032 33216
rect 52032 33152 52096 33216
rect 52096 33152 52112 33216
rect 52112 33152 52176 33216
rect 52176 33152 52192 33216
rect 52192 33152 52222 33216
rect 51986 33058 52222 33152
rect 51986 28058 52222 28294
rect 51986 23058 52222 23294
rect 51986 18058 52222 18294
rect 51986 13058 52222 13294
rect 51986 8192 52222 8294
rect 51986 8128 52016 8192
rect 52016 8128 52032 8192
rect 52032 8128 52096 8192
rect 52096 8128 52112 8192
rect 52112 8128 52176 8192
rect 52176 8128 52192 8192
rect 52192 8128 52222 8192
rect 51986 8058 52222 8128
rect 51986 3058 52222 3294
rect 52646 53718 52882 53954
rect 52646 48928 52676 48954
rect 52676 48928 52692 48954
rect 52692 48928 52756 48954
rect 52756 48928 52772 48954
rect 52772 48928 52836 48954
rect 52836 48928 52852 48954
rect 52852 48928 52882 48954
rect 52646 48718 52882 48928
rect 52646 43718 52882 43954
rect 52646 38718 52882 38954
rect 52646 33760 52882 33954
rect 52646 33718 52676 33760
rect 52676 33718 52692 33760
rect 52692 33718 52756 33760
rect 52756 33718 52772 33760
rect 52772 33718 52836 33760
rect 52836 33718 52852 33760
rect 52852 33718 52882 33760
rect 52646 28718 52882 28954
rect 52646 23904 52676 23954
rect 52676 23904 52692 23954
rect 52692 23904 52756 23954
rect 52756 23904 52772 23954
rect 52772 23904 52836 23954
rect 52836 23904 52852 23954
rect 52852 23904 52882 23954
rect 52646 23718 52882 23904
rect 52646 18718 52882 18954
rect 52646 13718 52882 13954
rect 52646 8736 52882 8954
rect 52646 8718 52676 8736
rect 52676 8718 52692 8736
rect 52692 8718 52756 8736
rect 52756 8718 52772 8736
rect 52772 8718 52836 8736
rect 52836 8718 52852 8736
rect 52852 8718 52882 8736
rect 52646 3718 52882 3954
rect 56986 53058 57222 53294
rect 56986 48058 57222 48294
rect 56986 43058 57222 43294
rect 56986 38058 57222 38294
rect 56986 33216 57222 33294
rect 56986 33152 57016 33216
rect 57016 33152 57032 33216
rect 57032 33152 57096 33216
rect 57096 33152 57112 33216
rect 57112 33152 57176 33216
rect 57176 33152 57192 33216
rect 57192 33152 57222 33216
rect 56986 33058 57222 33152
rect 56986 28058 57222 28294
rect 56986 23058 57222 23294
rect 56986 18058 57222 18294
rect 56986 13058 57222 13294
rect 56986 8192 57222 8294
rect 56986 8128 57016 8192
rect 57016 8128 57032 8192
rect 57032 8128 57096 8192
rect 57096 8128 57112 8192
rect 57112 8128 57176 8192
rect 57176 8128 57192 8192
rect 57192 8128 57222 8192
rect 56986 8058 57222 8128
rect 56986 3058 57222 3294
rect 57646 53718 57882 53954
rect 57646 48928 57676 48954
rect 57676 48928 57692 48954
rect 57692 48928 57756 48954
rect 57756 48928 57772 48954
rect 57772 48928 57836 48954
rect 57836 48928 57852 48954
rect 57852 48928 57882 48954
rect 57646 48718 57882 48928
rect 57646 43718 57882 43954
rect 57646 38718 57882 38954
rect 57646 33760 57882 33954
rect 57646 33718 57676 33760
rect 57676 33718 57692 33760
rect 57692 33718 57756 33760
rect 57756 33718 57772 33760
rect 57772 33718 57836 33760
rect 57836 33718 57852 33760
rect 57852 33718 57882 33760
rect 57646 28718 57882 28954
rect 57646 23904 57676 23954
rect 57676 23904 57692 23954
rect 57692 23904 57756 23954
rect 57756 23904 57772 23954
rect 57772 23904 57836 23954
rect 57836 23904 57852 23954
rect 57852 23904 57882 23954
rect 57646 23718 57882 23904
rect 57646 18718 57882 18954
rect 57646 13718 57882 13954
rect 57646 8736 57882 8954
rect 57646 8718 57676 8736
rect 57676 8718 57692 8736
rect 57692 8718 57756 8736
rect 57756 8718 57772 8736
rect 57772 8718 57836 8736
rect 57836 8718 57852 8736
rect 57852 8718 57882 8736
rect 57646 3718 57882 3954
<< metal5 >>
rect 1056 53954 58928 53996
rect 1056 53718 2646 53954
rect 2882 53718 7646 53954
rect 7882 53718 12646 53954
rect 12882 53718 17646 53954
rect 17882 53718 22646 53954
rect 22882 53718 27646 53954
rect 27882 53718 32646 53954
rect 32882 53718 37646 53954
rect 37882 53718 42646 53954
rect 42882 53718 47646 53954
rect 47882 53718 52646 53954
rect 52882 53718 57646 53954
rect 57882 53718 58928 53954
rect 1056 53676 58928 53718
rect 1056 53294 58928 53336
rect 1056 53058 1986 53294
rect 2222 53058 6986 53294
rect 7222 53058 11986 53294
rect 12222 53058 16986 53294
rect 17222 53058 21986 53294
rect 22222 53058 26986 53294
rect 27222 53058 31986 53294
rect 32222 53058 36986 53294
rect 37222 53058 41986 53294
rect 42222 53058 46986 53294
rect 47222 53058 51986 53294
rect 52222 53058 56986 53294
rect 57222 53058 58928 53294
rect 1056 53016 58928 53058
rect 1056 48954 58928 48996
rect 1056 48718 2646 48954
rect 2882 48718 7646 48954
rect 7882 48718 12646 48954
rect 12882 48718 17646 48954
rect 17882 48718 22646 48954
rect 22882 48718 27646 48954
rect 27882 48718 32646 48954
rect 32882 48718 37646 48954
rect 37882 48718 42646 48954
rect 42882 48718 47646 48954
rect 47882 48718 52646 48954
rect 52882 48718 57646 48954
rect 57882 48718 58928 48954
rect 1056 48676 58928 48718
rect 1056 48294 58928 48336
rect 1056 48058 1986 48294
rect 2222 48058 6986 48294
rect 7222 48058 11986 48294
rect 12222 48058 16986 48294
rect 17222 48058 21986 48294
rect 22222 48058 26986 48294
rect 27222 48058 31986 48294
rect 32222 48058 36986 48294
rect 37222 48058 41986 48294
rect 42222 48058 46986 48294
rect 47222 48058 51986 48294
rect 52222 48058 56986 48294
rect 57222 48058 58928 48294
rect 1056 48016 58928 48058
rect 1056 43954 58928 43996
rect 1056 43718 2646 43954
rect 2882 43718 7646 43954
rect 7882 43718 12646 43954
rect 12882 43718 17646 43954
rect 17882 43718 22646 43954
rect 22882 43718 27646 43954
rect 27882 43718 32646 43954
rect 32882 43718 37646 43954
rect 37882 43718 42646 43954
rect 42882 43718 47646 43954
rect 47882 43718 52646 43954
rect 52882 43718 57646 43954
rect 57882 43718 58928 43954
rect 1056 43676 58928 43718
rect 1056 43294 58928 43336
rect 1056 43058 1986 43294
rect 2222 43058 6986 43294
rect 7222 43058 11986 43294
rect 12222 43058 16986 43294
rect 17222 43058 21986 43294
rect 22222 43058 26986 43294
rect 27222 43058 31986 43294
rect 32222 43058 36986 43294
rect 37222 43058 41986 43294
rect 42222 43058 46986 43294
rect 47222 43058 51986 43294
rect 52222 43058 56986 43294
rect 57222 43058 58928 43294
rect 1056 43016 58928 43058
rect 1056 38954 58928 38996
rect 1056 38718 2646 38954
rect 2882 38718 7646 38954
rect 7882 38718 12646 38954
rect 12882 38718 17646 38954
rect 17882 38718 22646 38954
rect 22882 38718 27646 38954
rect 27882 38718 32646 38954
rect 32882 38718 37646 38954
rect 37882 38718 42646 38954
rect 42882 38718 47646 38954
rect 47882 38718 52646 38954
rect 52882 38718 57646 38954
rect 57882 38718 58928 38954
rect 1056 38676 58928 38718
rect 1056 38294 58928 38336
rect 1056 38058 1986 38294
rect 2222 38058 6986 38294
rect 7222 38058 11986 38294
rect 12222 38058 16986 38294
rect 17222 38058 21986 38294
rect 22222 38058 26986 38294
rect 27222 38058 31986 38294
rect 32222 38058 36986 38294
rect 37222 38058 41986 38294
rect 42222 38058 46986 38294
rect 47222 38058 51986 38294
rect 52222 38058 56986 38294
rect 57222 38058 58928 38294
rect 1056 38016 58928 38058
rect 1056 33954 58928 33996
rect 1056 33718 2646 33954
rect 2882 33718 7646 33954
rect 7882 33718 12646 33954
rect 12882 33718 17646 33954
rect 17882 33718 22646 33954
rect 22882 33718 27646 33954
rect 27882 33718 32646 33954
rect 32882 33718 37646 33954
rect 37882 33718 42646 33954
rect 42882 33718 47646 33954
rect 47882 33718 52646 33954
rect 52882 33718 57646 33954
rect 57882 33718 58928 33954
rect 1056 33676 58928 33718
rect 1056 33294 58928 33336
rect 1056 33058 1986 33294
rect 2222 33058 6986 33294
rect 7222 33058 11986 33294
rect 12222 33058 16986 33294
rect 17222 33058 21986 33294
rect 22222 33058 26986 33294
rect 27222 33058 31986 33294
rect 32222 33058 36986 33294
rect 37222 33058 41986 33294
rect 42222 33058 46986 33294
rect 47222 33058 51986 33294
rect 52222 33058 56986 33294
rect 57222 33058 58928 33294
rect 1056 33016 58928 33058
rect 1056 28954 58928 28996
rect 1056 28718 2646 28954
rect 2882 28718 7646 28954
rect 7882 28718 12646 28954
rect 12882 28718 17646 28954
rect 17882 28718 22646 28954
rect 22882 28718 27646 28954
rect 27882 28718 32646 28954
rect 32882 28718 37646 28954
rect 37882 28718 42646 28954
rect 42882 28718 47646 28954
rect 47882 28718 52646 28954
rect 52882 28718 57646 28954
rect 57882 28718 58928 28954
rect 1056 28676 58928 28718
rect 1056 28294 58928 28336
rect 1056 28058 1986 28294
rect 2222 28058 6986 28294
rect 7222 28058 11986 28294
rect 12222 28058 16986 28294
rect 17222 28058 21986 28294
rect 22222 28058 26986 28294
rect 27222 28058 31986 28294
rect 32222 28058 36986 28294
rect 37222 28058 41986 28294
rect 42222 28058 46986 28294
rect 47222 28058 51986 28294
rect 52222 28058 56986 28294
rect 57222 28058 58928 28294
rect 1056 28016 58928 28058
rect 1056 23954 58928 23996
rect 1056 23718 2646 23954
rect 2882 23718 7646 23954
rect 7882 23718 12646 23954
rect 12882 23718 17646 23954
rect 17882 23718 22646 23954
rect 22882 23718 27646 23954
rect 27882 23718 32646 23954
rect 32882 23718 37646 23954
rect 37882 23718 42646 23954
rect 42882 23718 47646 23954
rect 47882 23718 52646 23954
rect 52882 23718 57646 23954
rect 57882 23718 58928 23954
rect 1056 23676 58928 23718
rect 1056 23294 58928 23336
rect 1056 23058 1986 23294
rect 2222 23058 6986 23294
rect 7222 23058 11986 23294
rect 12222 23058 16986 23294
rect 17222 23058 21986 23294
rect 22222 23058 26986 23294
rect 27222 23058 31986 23294
rect 32222 23058 36986 23294
rect 37222 23058 41986 23294
rect 42222 23058 46986 23294
rect 47222 23058 51986 23294
rect 52222 23058 56986 23294
rect 57222 23058 58928 23294
rect 1056 23016 58928 23058
rect 1056 18954 58928 18996
rect 1056 18718 2646 18954
rect 2882 18718 7646 18954
rect 7882 18718 12646 18954
rect 12882 18718 17646 18954
rect 17882 18718 22646 18954
rect 22882 18718 27646 18954
rect 27882 18718 32646 18954
rect 32882 18718 37646 18954
rect 37882 18718 42646 18954
rect 42882 18718 47646 18954
rect 47882 18718 52646 18954
rect 52882 18718 57646 18954
rect 57882 18718 58928 18954
rect 1056 18676 58928 18718
rect 1056 18294 58928 18336
rect 1056 18058 1986 18294
rect 2222 18058 6986 18294
rect 7222 18058 11986 18294
rect 12222 18058 16986 18294
rect 17222 18058 21986 18294
rect 22222 18058 26986 18294
rect 27222 18058 31986 18294
rect 32222 18058 36986 18294
rect 37222 18058 41986 18294
rect 42222 18058 46986 18294
rect 47222 18058 51986 18294
rect 52222 18058 56986 18294
rect 57222 18058 58928 18294
rect 1056 18016 58928 18058
rect 1056 13954 58928 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 22646 13954
rect 22882 13718 27646 13954
rect 27882 13718 32646 13954
rect 32882 13718 37646 13954
rect 37882 13718 42646 13954
rect 42882 13718 47646 13954
rect 47882 13718 52646 13954
rect 52882 13718 57646 13954
rect 57882 13718 58928 13954
rect 1056 13676 58928 13718
rect 1056 13294 58928 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 21986 13294
rect 22222 13058 26986 13294
rect 27222 13058 31986 13294
rect 32222 13058 36986 13294
rect 37222 13058 41986 13294
rect 42222 13058 46986 13294
rect 47222 13058 51986 13294
rect 52222 13058 56986 13294
rect 57222 13058 58928 13294
rect 1056 13016 58928 13058
rect 1056 8954 58928 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 22646 8954
rect 22882 8718 27646 8954
rect 27882 8718 32646 8954
rect 32882 8718 37646 8954
rect 37882 8718 42646 8954
rect 42882 8718 47646 8954
rect 47882 8718 52646 8954
rect 52882 8718 57646 8954
rect 57882 8718 58928 8954
rect 1056 8676 58928 8718
rect 1056 8294 58928 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 21986 8294
rect 22222 8058 26986 8294
rect 27222 8058 31986 8294
rect 32222 8058 36986 8294
rect 37222 8058 41986 8294
rect 42222 8058 46986 8294
rect 47222 8058 51986 8294
rect 52222 8058 56986 8294
rect 57222 8058 58928 8294
rect 1056 8016 58928 8058
rect 1056 3954 58928 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 22646 3954
rect 22882 3718 27646 3954
rect 27882 3718 32646 3954
rect 32882 3718 37646 3954
rect 37882 3718 42646 3954
rect 42882 3718 47646 3954
rect 47882 3718 52646 3954
rect 52882 3718 57646 3954
rect 57882 3718 58928 3954
rect 1056 3676 58928 3718
rect 1056 3294 58928 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 21986 3294
rect 22222 3058 26986 3294
rect 27222 3058 31986 3294
rect 32222 3058 36986 3294
rect 37222 3058 41986 3294
rect 42222 3058 46986 3294
rect 47222 3058 51986 3294
rect 52222 3058 56986 3294
rect 57222 3058 58928 3294
rect 1056 3016 58928 3058
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 0
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 0
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 0
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 0
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 0
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 0
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 0
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 0
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 0
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 0
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 0
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 0
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 0
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 0
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 0
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 0
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 0
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 0
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 0
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 0
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_461
timestamp 0
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 0
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_477
timestamp 0
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_489
timestamp 0
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 0
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_505
timestamp 0
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_517
timestamp 0
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 0
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_533
timestamp 0
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_545
timestamp 0
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 0
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_561
timestamp 0
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_573
timestamp 0
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 0
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_589
timestamp 0
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_601
timestamp 0
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 0
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_617
timestamp 0
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 0
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 0
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 0
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 0
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 0
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 0
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 0
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 0
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 0
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 0
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 0
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 0
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 0
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 0
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 0
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 0
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 0
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 0
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 0
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 0
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 0
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 0
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 0
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 0
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 0
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 0
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 0
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_473
timestamp 0
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_485
timestamp 0
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_497
timestamp 0
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 0
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_505
timestamp 0
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_517
timestamp 0
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_529
timestamp 0
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_541
timestamp 0
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_553
timestamp 0
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 0
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_561
timestamp 0
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_573
timestamp 0
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_585
timestamp 0
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_597
timestamp 0
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_609
timestamp 0
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_615
timestamp 0
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_617
timestamp 0
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 0
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 0
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 0
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 0
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 0
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 0
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 0
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 0
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 0
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 0
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 0
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 0
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 0
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 0
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 0
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 0
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 0
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 0
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 0
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 0
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 0
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 0
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 0
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 0
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 0
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 0
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_469
timestamp 0
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 0
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 0
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 0
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 0
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 0
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 0
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 0
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 0
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 0
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 0
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_569
timestamp 0
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_581
timestamp 0
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 0
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_589
timestamp 0
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_601
timestamp 0
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_613
timestamp 0
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 0
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 0
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 0
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 0
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 0
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 0
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 0
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 0
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 0
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 0
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 0
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 0
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 0
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 0
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 0
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 0
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 0
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 0
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 0
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 0
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 0
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 0
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 0
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 0
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 0
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 0
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 0
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 0
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 0
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_505
timestamp 0
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_517
timestamp 0
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 0
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 0
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 0
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 0
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 0
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 0
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 0
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_597
timestamp 0
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_609
timestamp 0
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 0
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_617
timestamp 0
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 0
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 0
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 0
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 0
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 0
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 0
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 0
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 0
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 0
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 0
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 0
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 0
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 0
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 0
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 0
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 0
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 0
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 0
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 0
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 0
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 0
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 0
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 0
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 0
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 0
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 0
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 0
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 0
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 0
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 0
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 0
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 0
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 0
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_501
timestamp 0
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_513
timestamp 0
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_525
timestamp 0
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 0
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 0
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 0
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 0
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 0
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 0
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 0
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 0
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 0
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_613
timestamp 0
transform 1 0 57500 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_621
timestamp 0
transform 1 0 58236 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 0
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 0
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 0
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 0
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 0
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 0
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 0
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 0
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 0
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 0
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 0
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 0
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 0
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 0
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 0
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 0
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 0
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 0
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 0
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 0
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 0
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 0
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 0
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 0
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 0
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 0
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 0
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 0
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 0
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 0
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 0
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 0
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 0
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 0
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_517
timestamp 0
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_529
timestamp 0
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_541
timestamp 0
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 0
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 0
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 0
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 0
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 0
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 0
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 0
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 0
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_617
timestamp 0
transform 1 0 57868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_621
timestamp 0
transform 1 0 58236 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 0
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 0
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 0
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 0
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 0
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 0
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 0
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 0
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 0
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 0
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 0
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 0
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 0
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 0
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 0
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 0
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 0
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 0
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 0
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 0
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 0
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 0
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 0
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 0
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 0
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 0
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 0
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 0
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 0
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 0
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 0
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 0
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 0
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 0
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 0
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_489
timestamp 0
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_501
timestamp 0
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_513
timestamp 0
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_525
timestamp 0
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 0
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 0
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 0
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 0
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 0
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 0
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 0
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 0
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 0
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 0
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 0
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 0
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 0
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 0
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 0
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 0
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 0
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 0
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 0
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 0
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 0
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 0
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 0
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 0
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 0
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 0
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 0
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 0
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 0
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 0
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 0
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 0
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 0
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 0
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 0
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 0
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 0
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 0
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_473
timestamp 0
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_485
timestamp 0
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_497
timestamp 0
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_503
timestamp 0
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_505
timestamp 0
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_517
timestamp 0
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_529
timestamp 0
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_541
timestamp 0
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_553
timestamp 0
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 0
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_561
timestamp 0
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_573
timestamp 0
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_585
timestamp 0
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_597
timestamp 0
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 0
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 0
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_617
timestamp 0
transform 1 0 57868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_621
timestamp 0
transform 1 0 58236 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 0
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 0
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 0
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 0
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 0
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 0
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 0
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 0
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 0
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 0
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 0
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 0
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 0
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 0
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 0
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 0
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 0
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 0
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 0
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 0
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 0
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 0
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 0
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 0
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 0
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 0
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 0
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 0
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 0
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 0
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 0
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 0
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 0
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_489
timestamp 0
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_501
timestamp 0
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_513
timestamp 0
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_525
timestamp 0
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 0
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_533
timestamp 0
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_545
timestamp 0
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_557
timestamp 0
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 0
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 0
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 0
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 0
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 0
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_613
timestamp 0
transform 1 0 57500 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_621
timestamp 0
transform 1 0 58236 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 0
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 0
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 0
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 0
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 0
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 0
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 0
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 0
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 0
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 0
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 0
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 0
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 0
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 0
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 0
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 0
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 0
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 0
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 0
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 0
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 0
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 0
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 0
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 0
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 0
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 0
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 0
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 0
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 0
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 0
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 0
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_485
timestamp 0
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_497
timestamp 0
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 0
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 0
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_517
timestamp 0
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_529
timestamp 0
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_541
timestamp 0
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_553
timestamp 0
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_559
timestamp 0
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_561
timestamp 0
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 0
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 0
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 0
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 0
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 0
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_617
timestamp 0
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 0
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 0
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 0
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 0
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 0
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 0
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 0
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 0
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 0
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 0
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 0
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 0
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 0
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 0
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 0
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 0
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 0
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 0
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 0
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 0
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 0
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 0
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 0
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 0
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 0
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 0
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 0
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 0
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 0
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 0
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 0
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 0
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 0
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 0
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_489
timestamp 0
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_501
timestamp 0
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_513
timestamp 0
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_525
timestamp 0
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_531
timestamp 0
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 0
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 0
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 0
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 0
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 0
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 0
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 0
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 0
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_613
timestamp 0
transform 1 0 57500 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_621
timestamp 0
transform 1 0 58236 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 0
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 0
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 0
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 0
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 0
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 0
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 0
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 0
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 0
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 0
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 0
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 0
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 0
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 0
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 0
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 0
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 0
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 0
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 0
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 0
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 0
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 0
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 0
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 0
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 0
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 0
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 0
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 0
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 0
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 0
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 0
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 0
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_473
timestamp 0
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_485
timestamp 0
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_497
timestamp 0
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 0
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_505
timestamp 0
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 0
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_529
timestamp 0
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_541
timestamp 0
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_553
timestamp 0
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 0
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 0
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 0
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 0
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 0
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 0
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 0
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_617
timestamp 0
transform 1 0 57868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_621
timestamp 0
transform 1 0 58236 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 0
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 0
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 0
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 0
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 0
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 0
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 0
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 0
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 0
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 0
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 0
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 0
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 0
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 0
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 0
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 0
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 0
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 0
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 0
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 0
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 0
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 0
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 0
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 0
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 0
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 0
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 0
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 0
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 0
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 0
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 0
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 0
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 0
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_489
timestamp 0
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_501
timestamp 0
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_513
timestamp 0
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_525
timestamp 0
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 0
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 0
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 0
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 0
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 0
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 0
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 0
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 0
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 0
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 0
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 0
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 0
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 0
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 0
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 0
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 0
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 0
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 0
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 0
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 0
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 0
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 0
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 0
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 0
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 0
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 0
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 0
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 0
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 0
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 0
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 0
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 0
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 0
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 0
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 0
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 0
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 0
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 0
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 0
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 0
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 0
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_473
timestamp 0
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_485
timestamp 0
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_497
timestamp 0
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 0
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 0
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_517
timestamp 0
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_529
timestamp 0
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_541
timestamp 0
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 0
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 0
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_561
timestamp 0
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_573
timestamp 0
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_585
timestamp 0
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_597
timestamp 0
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_609
timestamp 0
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 0
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_617
timestamp 0
transform 1 0 57868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_621
timestamp 0
transform 1 0 58236 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 0
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 0
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 0
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 0
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 0
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 0
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 0
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 0
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 0
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 0
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 0
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 0
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 0
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 0
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 0
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 0
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 0
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 0
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 0
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 0
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 0
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 0
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 0
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_401
timestamp 0
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_413
timestamp 0
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 0
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 0
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_433
timestamp 0
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 0
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_457
timestamp 0
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_469
timestamp 0
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 0
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_477
timestamp 0
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_489
timestamp 0
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_501
timestamp 0
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_513
timestamp 0
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_525
timestamp 0
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 0
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_533
timestamp 0
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_545
timestamp 0
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_557
timestamp 0
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_569
timestamp 0
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_581
timestamp 0
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_587
timestamp 0
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_589
timestamp 0
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_601
timestamp 0
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_613
timestamp 0
transform 1 0 57500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_621
timestamp 0
transform 1 0 58236 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 0
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 0
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 0
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 0
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 0
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 0
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 0
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 0
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 0
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 0
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 0
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 0
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 0
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 0
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 0
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 0
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 0
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 0
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 0
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 0
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 0
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 0
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 0
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 0
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_429
timestamp 0
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_441
timestamp 0
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_447
timestamp 0
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 0
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_461
timestamp 0
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_473
timestamp 0
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_485
timestamp 0
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_497
timestamp 0
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_503
timestamp 0
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_505
timestamp 0
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_517
timestamp 0
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_529
timestamp 0
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_541
timestamp 0
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_553
timestamp 0
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_559
timestamp 0
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_561
timestamp 0
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_573
timestamp 0
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_585
timestamp 0
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_597
timestamp 0
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_609
timestamp 0
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_615
timestamp 0
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_617
timestamp 0
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 0
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 0
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 0
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 0
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 0
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 0
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 0
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 0
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 0
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 0
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 0
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 0
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 0
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 0
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 0
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 0
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 0
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 0
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 0
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 0
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 0
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_401
timestamp 0
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_413
timestamp 0
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 0
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 0
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 0
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_445
timestamp 0
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_457
timestamp 0
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_469
timestamp 0
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_475
timestamp 0
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_477
timestamp 0
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_489
timestamp 0
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_501
timestamp 0
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_513
timestamp 0
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_525
timestamp 0
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_531
timestamp 0
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_533
timestamp 0
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_545
timestamp 0
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_557
timestamp 0
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_569
timestamp 0
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_581
timestamp 0
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_587
timestamp 0
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_589
timestamp 0
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_601
timestamp 0
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_613
timestamp 0
transform 1 0 57500 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_621
timestamp 0
transform 1 0 58236 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 0
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 0
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 0
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 0
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 0
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 0
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 0
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 0
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 0
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 0
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 0
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 0
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 0
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 0
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 0
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 0
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 0
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 0
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 0
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 0
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 0
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 0
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 0
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 0
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 0
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_429
timestamp 0
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_441
timestamp 0
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 0
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 0
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_461
timestamp 0
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_473
timestamp 0
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_485
timestamp 0
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_497
timestamp 0
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_503
timestamp 0
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_505
timestamp 0
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_517
timestamp 0
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_529
timestamp 0
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_541
timestamp 0
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_553
timestamp 0
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_559
timestamp 0
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_561
timestamp 0
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_573
timestamp 0
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_585
timestamp 0
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_597
timestamp 0
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_609
timestamp 0
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 0
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_617
timestamp 0
transform 1 0 57868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_621
timestamp 0
transform 1 0 58236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 0
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 0
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 0
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 0
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 0
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 0
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 0
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 0
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 0
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 0
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 0
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 0
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 0
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 0
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 0
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 0
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 0
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 0
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 0
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 0
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 0
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 0
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 0
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 0
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 0
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 0
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 0
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 0
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_457
timestamp 0
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_469
timestamp 0
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 0
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_477
timestamp 0
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_489
timestamp 0
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_501
timestamp 0
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_513
timestamp 0
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_525
timestamp 0
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_531
timestamp 0
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_533
timestamp 0
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_545
timestamp 0
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_557
timestamp 0
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_569
timestamp 0
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_581
timestamp 0
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_587
timestamp 0
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_589
timestamp 0
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_601
timestamp 0
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_613
timestamp 0
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 0
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 0
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 0
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 0
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 0
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 0
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 0
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 0
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 0
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 0
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 0
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 0
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 0
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 0
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 0
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 0
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 0
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 0
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 0
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 0
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 0
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 0
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 0
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 0
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 0
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 0
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_405
timestamp 0
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_417
timestamp 0
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_429
timestamp 0
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_441
timestamp 0
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 0
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_449
timestamp 0
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_461
timestamp 0
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_473
timestamp 0
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_485
timestamp 0
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_497
timestamp 0
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_503
timestamp 0
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_505
timestamp 0
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_517
timestamp 0
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_529
timestamp 0
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_541
timestamp 0
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_553
timestamp 0
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_559
timestamp 0
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_561
timestamp 0
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_573
timestamp 0
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_585
timestamp 0
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_597
timestamp 0
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_609
timestamp 0
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_615
timestamp 0
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_617
timestamp 0
transform 1 0 57868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_621
timestamp 0
transform 1 0 58236 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 0
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 0
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 0
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 0
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 0
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 0
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 0
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 0
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 0
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 0
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 0
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 0
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 0
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 0
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 0
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 0
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 0
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 0
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 0
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 0
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 0
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 0
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 0
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 0
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 0
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_401
timestamp 0
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_413
timestamp 0
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_419
timestamp 0
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_421
timestamp 0
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_433
timestamp 0
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_445
timestamp 0
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_457
timestamp 0
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_469
timestamp 0
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_475
timestamp 0
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_477
timestamp 0
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_489
timestamp 0
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_501
timestamp 0
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_513
timestamp 0
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_525
timestamp 0
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_531
timestamp 0
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_533
timestamp 0
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_545
timestamp 0
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_557
timestamp 0
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_569
timestamp 0
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_581
timestamp 0
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_587
timestamp 0
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_589
timestamp 0
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_601
timestamp 0
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_613
timestamp 0
transform 1 0 57500 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_621
timestamp 0
transform 1 0 58236 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 0
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 0
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 0
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 0
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 0
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 0
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 0
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 0
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 0
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 0
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 0
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 0
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 0
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 0
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 0
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 0
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 0
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 0
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 0
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 0
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 0
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 0
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 0
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 0
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_417
timestamp 0
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_429
timestamp 0
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_441
timestamp 0
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_447
timestamp 0
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 0
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_461
timestamp 0
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_473
timestamp 0
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_485
timestamp 0
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_497
timestamp 0
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_503
timestamp 0
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_505
timestamp 0
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_517
timestamp 0
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_529
timestamp 0
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_541
timestamp 0
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_553
timestamp 0
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_559
timestamp 0
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_561
timestamp 0
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_573
timestamp 0
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_585
timestamp 0
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_597
timestamp 0
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_609
timestamp 0
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_615
timestamp 0
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_617
timestamp 0
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 0
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 0
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 0
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 0
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 0
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 0
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 0
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 0
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 0
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 0
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 0
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 0
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 0
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 0
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 0
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 0
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 0
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 0
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 0
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 0
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 0
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 0
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_401
timestamp 0
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 0
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 0
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 0
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_433
timestamp 0
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_445
timestamp 0
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_457
timestamp 0
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_469
timestamp 0
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_475
timestamp 0
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_477
timestamp 0
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_489
timestamp 0
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_501
timestamp 0
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_513
timestamp 0
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_525
timestamp 0
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_531
timestamp 0
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_533
timestamp 0
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_545
timestamp 0
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_557
timestamp 0
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_569
timestamp 0
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_581
timestamp 0
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_587
timestamp 0
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_589
timestamp 0
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_601
timestamp 0
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_613
timestamp 0
transform 1 0 57500 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_621
timestamp 0
transform 1 0 58236 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 0
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 0
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 0
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 0
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 0
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 0
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 0
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 0
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 0
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 0
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 0
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 0
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 0
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 0
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 0
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 0
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 0
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 0
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 0
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 0
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 0
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 0
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_405
timestamp 0
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_417
timestamp 0
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_429
timestamp 0
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_441
timestamp 0
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 0
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_449
timestamp 0
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_461
timestamp 0
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_473
timestamp 0
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_485
timestamp 0
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_497
timestamp 0
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_503
timestamp 0
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_505
timestamp 0
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_517
timestamp 0
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_529
timestamp 0
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_541
timestamp 0
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_553
timestamp 0
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_559
timestamp 0
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_561
timestamp 0
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_573
timestamp 0
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_585
timestamp 0
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_597
timestamp 0
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_609
timestamp 0
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_615
timestamp 0
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_617
timestamp 0
transform 1 0 57868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_621
timestamp 0
transform 1 0 58236 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 0
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 0
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 0
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 0
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 0
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 0
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 0
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 0
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 0
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 0
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 0
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 0
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 0
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 0
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 0
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 0
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 0
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 0
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 0
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 0
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 0
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 0
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 0
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 0
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_421
timestamp 0
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_433
timestamp 0
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_445
timestamp 0
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_457
timestamp 0
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_469
timestamp 0
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_475
timestamp 0
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_477
timestamp 0
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_489
timestamp 0
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_501
timestamp 0
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_513
timestamp 0
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_525
timestamp 0
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_531
timestamp 0
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_533
timestamp 0
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_545
timestamp 0
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_557
timestamp 0
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_569
timestamp 0
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_581
timestamp 0
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_587
timestamp 0
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_589
timestamp 0
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_601
timestamp 0
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_613
timestamp 0
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 0
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 0
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 0
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 0
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 0
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 0
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 0
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 0
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 0
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 0
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 0
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 0
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 0
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 0
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 0
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 0
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 0
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 0
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 0
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 0
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 0
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 0
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 0
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 0
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 0
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 0
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 0
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_429
timestamp 0
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_441
timestamp 0
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 0
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_449
timestamp 0
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_461
timestamp 0
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_473
timestamp 0
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_485
timestamp 0
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_497
timestamp 0
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_503
timestamp 0
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_505
timestamp 0
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_517
timestamp 0
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_529
timestamp 0
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_541
timestamp 0
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_553
timestamp 0
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_559
timestamp 0
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_561
timestamp 0
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_573
timestamp 0
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_585
timestamp 0
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_597
timestamp 0
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_609
timestamp 0
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_615
timestamp 0
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_617
timestamp 0
transform 1 0 57868 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_621
timestamp 0
transform 1 0 58236 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 0
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 0
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 0
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 0
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 0
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 0
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 0
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 0
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 0
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 0
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 0
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 0
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 0
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 0
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 0
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 0
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 0
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 0
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 0
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 0
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_401
timestamp 0
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_413
timestamp 0
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 0
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 0
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_433
timestamp 0
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_445
timestamp 0
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_457
timestamp 0
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_469
timestamp 0
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_475
timestamp 0
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_477
timestamp 0
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_489
timestamp 0
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_501
timestamp 0
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_513
timestamp 0
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_525
timestamp 0
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_531
timestamp 0
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_533
timestamp 0
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_545
timestamp 0
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_557
timestamp 0
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_569
timestamp 0
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_581
timestamp 0
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_587
timestamp 0
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_589
timestamp 0
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_601
timestamp 0
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_613
timestamp 0
transform 1 0 57500 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_621
timestamp 0
transform 1 0 58236 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 0
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 0
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 0
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 0
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 0
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 0
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 0
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 0
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 0
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 0
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 0
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 0
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 0
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 0
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 0
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 0
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 0
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 0
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 0
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 0
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 0
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 0
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 0
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 0
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 0
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 0
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 0
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 0
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 0
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_417
timestamp 0
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_429
timestamp 0
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_441
timestamp 0
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_447
timestamp 0
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_449
timestamp 0
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_461
timestamp 0
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_473
timestamp 0
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_485
timestamp 0
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_497
timestamp 0
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_503
timestamp 0
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_505
timestamp 0
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_517
timestamp 0
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_529
timestamp 0
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_541
timestamp 0
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_553
timestamp 0
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_559
timestamp 0
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_561
timestamp 0
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_573
timestamp 0
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_585
timestamp 0
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_597
timestamp 0
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_609
timestamp 0
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_615
timestamp 0
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_617
timestamp 0
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 0
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 0
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 0
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 0
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 0
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 0
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 0
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 0
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 0
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 0
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 0
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 0
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 0
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 0
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 0
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 0
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 0
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 0
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 0
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 0
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 0
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 0
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 0
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 0
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 0
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 0
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 0
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_401
timestamp 0
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_413
timestamp 0
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 0
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 0
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 0
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_445
timestamp 0
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_457
timestamp 0
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_469
timestamp 0
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_475
timestamp 0
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_477
timestamp 0
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_489
timestamp 0
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_501
timestamp 0
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_513
timestamp 0
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_525
timestamp 0
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_531
timestamp 0
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_533
timestamp 0
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_545
timestamp 0
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_557
timestamp 0
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_569
timestamp 0
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_581
timestamp 0
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_587
timestamp 0
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_589
timestamp 0
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_601
timestamp 0
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_613
timestamp 0
transform 1 0 57500 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_621
timestamp 0
transform 1 0 58236 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 0
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 0
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 0
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 0
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 0
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 0
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 0
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 0
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 0
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 0
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 0
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 0
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 0
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 0
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 0
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 0
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 0
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 0
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 0
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 0
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 0
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 0
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 0
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 0
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 0
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 0
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_405
timestamp 0
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_417
timestamp 0
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_429
timestamp 0
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_441
timestamp 0
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 0
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 0
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_461
timestamp 0
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_473
timestamp 0
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_485
timestamp 0
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_497
timestamp 0
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_503
timestamp 0
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_505
timestamp 0
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_517
timestamp 0
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_529
timestamp 0
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_541
timestamp 0
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_553
timestamp 0
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_559
timestamp 0
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_561
timestamp 0
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_573
timestamp 0
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_585
timestamp 0
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_597
timestamp 0
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_609
timestamp 0
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_615
timestamp 0
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_617
timestamp 0
transform 1 0 57868 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_621
timestamp 0
transform 1 0 58236 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 0
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 0
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 0
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 0
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 0
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 0
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 0
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 0
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 0
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 0
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 0
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 0
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 0
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 0
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 0
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 0
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 0
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 0
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 0
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 0
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 0
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 0
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 0
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 0
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 0
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 0
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 0
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_401
timestamp 0
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_413
timestamp 0
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 0
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_421
timestamp 0
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_433
timestamp 0
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_445
timestamp 0
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_457
timestamp 0
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_469
timestamp 0
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 0
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_477
timestamp 0
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_489
timestamp 0
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_501
timestamp 0
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_513
timestamp 0
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_525
timestamp 0
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_531
timestamp 0
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_533
timestamp 0
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_545
timestamp 0
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_557
timestamp 0
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_569
timestamp 0
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_581
timestamp 0
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_587
timestamp 0
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 0
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_601
timestamp 0
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_613
timestamp 0
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 0
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 0
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 0
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 0
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 0
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 0
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 0
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 0
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 0
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 0
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 0
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 0
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 0
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 0
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 0
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 0
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 0
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 0
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 0
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 0
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 0
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 0
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 0
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 0
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 0
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 0
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 0
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 0
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 0
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 0
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 0
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 0
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 0
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 0
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_429
timestamp 0
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_441
timestamp 0
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 0
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_449
timestamp 0
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_461
timestamp 0
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_473
timestamp 0
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_485
timestamp 0
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_497
timestamp 0
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_503
timestamp 0
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_505
timestamp 0
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_517
timestamp 0
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_529
timestamp 0
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_541
timestamp 0
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_553
timestamp 0
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_559
timestamp 0
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_561
timestamp 0
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_573
timestamp 0
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_585
timestamp 0
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_597
timestamp 0
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_609
timestamp 0
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_615
timestamp 0
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_617
timestamp 0
transform 1 0 57868 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_621
timestamp 0
transform 1 0 58236 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 0
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 0
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 0
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 0
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 0
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 0
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 0
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 0
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 0
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 0
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 0
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 0
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 0
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 0
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 0
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 0
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 0
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 0
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 0
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 0
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 0
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 0
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 0
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 0
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 0
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 0
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_401
timestamp 0
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_413
timestamp 0
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 0
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 0
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_433
timestamp 0
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_445
timestamp 0
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_457
timestamp 0
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_469
timestamp 0
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_475
timestamp 0
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_477
timestamp 0
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_489
timestamp 0
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_501
timestamp 0
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_513
timestamp 0
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_525
timestamp 0
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_531
timestamp 0
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_533
timestamp 0
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_545
timestamp 0
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_557
timestamp 0
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_569
timestamp 0
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_581
timestamp 0
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_587
timestamp 0
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_589
timestamp 0
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_601
timestamp 0
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_613
timestamp 0
transform 1 0 57500 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_621
timestamp 0
transform 1 0 58236 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 0
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 0
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 0
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 0
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 0
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 0
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 0
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 0
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 0
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 0
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 0
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 0
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 0
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 0
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 0
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 0
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 0
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 0
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 0
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 0
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 0
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 0
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 0
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 0
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 0
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 0
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 0
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 0
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 0
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 0
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 0
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 0
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_405
timestamp 0
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_417
timestamp 0
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_429
timestamp 0
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_441
timestamp 0
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 0
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 0
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_461
timestamp 0
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_473
timestamp 0
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_485
timestamp 0
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_497
timestamp 0
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_503
timestamp 0
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_505
timestamp 0
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_517
timestamp 0
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_529
timestamp 0
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_541
timestamp 0
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_553
timestamp 0
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_559
timestamp 0
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_561
timestamp 0
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_573
timestamp 0
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_585
timestamp 0
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_597
timestamp 0
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_609
timestamp 0
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_615
timestamp 0
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_617
timestamp 0
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 0
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 0
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 0
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 0
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 0
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 0
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 0
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 0
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 0
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 0
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 0
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 0
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 0
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 0
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 0
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 0
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 0
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 0
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 0
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 0
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 0
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 0
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 0
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 0
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 0
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 0
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 0
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 0
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 0
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 0
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 0
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_401
timestamp 0
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_413
timestamp 0
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 0
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 0
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_433
timestamp 0
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_445
timestamp 0
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_457
timestamp 0
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_469
timestamp 0
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 0
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_477
timestamp 0
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_489
timestamp 0
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_501
timestamp 0
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_513
timestamp 0
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_525
timestamp 0
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_531
timestamp 0
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_533
timestamp 0
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_545
timestamp 0
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_557
timestamp 0
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_569
timestamp 0
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_581
timestamp 0
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_587
timestamp 0
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_589
timestamp 0
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_601
timestamp 0
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_613
timestamp 0
transform 1 0 57500 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_621
timestamp 0
transform 1 0 58236 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 0
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 0
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 0
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 0
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 0
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 0
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 0
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 0
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 0
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 0
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 0
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 0
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 0
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 0
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 0
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 0
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 0
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 0
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 0
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 0
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 0
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 0
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 0
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 0
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 0
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 0
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 0
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 0
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 0
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 0
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 0
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 0
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 0
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 0
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_429
timestamp 0
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_441
timestamp 0
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_447
timestamp 0
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_449
timestamp 0
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_461
timestamp 0
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_473
timestamp 0
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_485
timestamp 0
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_497
timestamp 0
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_503
timestamp 0
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_505
timestamp 0
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_517
timestamp 0
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_529
timestamp 0
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_541
timestamp 0
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_553
timestamp 0
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_559
timestamp 0
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_561
timestamp 0
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_573
timestamp 0
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_585
timestamp 0
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_597
timestamp 0
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_609
timestamp 0
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_615
timestamp 0
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_617
timestamp 0
transform 1 0 57868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_621
timestamp 0
transform 1 0 58236 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 0
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 0
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 0
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 0
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 0
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 0
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 0
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 0
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 0
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 0
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 0
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 0
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 0
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 0
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 0
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 0
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 0
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 0
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 0
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 0
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 0
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 0
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 0
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 0
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 0
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 0
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 0
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_401
timestamp 0
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_413
timestamp 0
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 0
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 0
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_433
timestamp 0
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_445
timestamp 0
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_457
timestamp 0
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_469
timestamp 0
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_475
timestamp 0
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_477
timestamp 0
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_489
timestamp 0
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_501
timestamp 0
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_513
timestamp 0
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_525
timestamp 0
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_531
timestamp 0
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_533
timestamp 0
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_545
timestamp 0
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_557
timestamp 0
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_569
timestamp 0
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_581
timestamp 0
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_587
timestamp 0
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_589
timestamp 0
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_601
timestamp 0
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_613
timestamp 0
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 0
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 0
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 0
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 0
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 0
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 0
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 0
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 0
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 0
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 0
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 0
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 0
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 0
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 0
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 0
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 0
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 0
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 0
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 0
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 0
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 0
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 0
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 0
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 0
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 0
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 0
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 0
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 0
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 0
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 0
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 0
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 0
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 0
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 0
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_405
timestamp 0
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_417
timestamp 0
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_429
timestamp 0
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_441
timestamp 0
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_447
timestamp 0
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 0
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_461
timestamp 0
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_473
timestamp 0
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_485
timestamp 0
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_497
timestamp 0
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_503
timestamp 0
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_505
timestamp 0
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_517
timestamp 0
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_529
timestamp 0
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_541
timestamp 0
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_553
timestamp 0
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_559
timestamp 0
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_561
timestamp 0
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_573
timestamp 0
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_585
timestamp 0
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_597
timestamp 0
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_609
timestamp 0
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_615
timestamp 0
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_617
timestamp 0
transform 1 0 57868 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_621
timestamp 0
transform 1 0 58236 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 0
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 0
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 0
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 0
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 0
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 0
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 0
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 0
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 0
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 0
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 0
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 0
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 0
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 0
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 0
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 0
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 0
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 0
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 0
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 0
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 0
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 0
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 0
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 0
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 0
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 0
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 0
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 0
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 0
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 0
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 0
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 0
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 0
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 0
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_401
timestamp 0
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_413
timestamp 0
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 0
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_421
timestamp 0
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_433
timestamp 0
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_445
timestamp 0
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_457
timestamp 0
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_469
timestamp 0
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_475
timestamp 0
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_477
timestamp 0
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_489
timestamp 0
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_501
timestamp 0
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_513
timestamp 0
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_525
timestamp 0
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_531
timestamp 0
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_533
timestamp 0
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_545
timestamp 0
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_557
timestamp 0
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_569
timestamp 0
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_581
timestamp 0
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_587
timestamp 0
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_589
timestamp 0
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_601
timestamp 0
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_613
timestamp 0
transform 1 0 57500 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_621
timestamp 0
transform 1 0 58236 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 0
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 0
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 0
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 0
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 0
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 0
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 0
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 0
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 0
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 0
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 0
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 0
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 0
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 0
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 0
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 0
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 0
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 0
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 0
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 0
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 0
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 0
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 0
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 0
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 0
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 0
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 0
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 0
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 0
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 0
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 0
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 0
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 0
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_429
timestamp 0
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_441
timestamp 0
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 0
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_449
timestamp 0
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_461
timestamp 0
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_473
timestamp 0
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_485
timestamp 0
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_497
timestamp 0
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_503
timestamp 0
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_505
timestamp 0
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_517
timestamp 0
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_529
timestamp 0
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_541
timestamp 0
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_553
timestamp 0
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_559
timestamp 0
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_561
timestamp 0
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_573
timestamp 0
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_585
timestamp 0
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_597
timestamp 0
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_609
timestamp 0
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 0
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_617
timestamp 0
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 0
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 0
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 0
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 0
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 0
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 0
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 0
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 0
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 0
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 0
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 0
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 0
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 0
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 0
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 0
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 0
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 0
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 0
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 0
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 0
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 0
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 0
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 0
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 0
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 0
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 0
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 0
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 0
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 0
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 0
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 0
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 0
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 0
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_401
timestamp 0
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_413
timestamp 0
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 0
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 0
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_433
timestamp 0
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_445
timestamp 0
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_457
timestamp 0
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_469
timestamp 0
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_475
timestamp 0
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_477
timestamp 0
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_489
timestamp 0
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_501
timestamp 0
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_513
timestamp 0
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_525
timestamp 0
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_531
timestamp 0
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_533
timestamp 0
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_545
timestamp 0
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_557
timestamp 0
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_569
timestamp 0
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_581
timestamp 0
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_587
timestamp 0
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_589
timestamp 0
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_601
timestamp 0
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_613
timestamp 0
transform 1 0 57500 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_621
timestamp 0
transform 1 0 58236 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 0
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 0
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 0
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 0
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 0
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 0
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 0
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 0
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 0
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 0
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 0
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 0
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 0
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 0
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 0
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 0
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 0
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 0
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 0
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 0
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 0
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 0
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 0
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 0
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 0
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 0
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 0
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 0
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 0
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 0
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 0
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 0
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 0
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 0
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 0
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 0
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 0
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 0
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 0
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_429
timestamp 0
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_441
timestamp 0
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_447
timestamp 0
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 0
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_461
timestamp 0
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_473
timestamp 0
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_485
timestamp 0
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_497
timestamp 0
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 0
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_505
timestamp 0
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_517
timestamp 0
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_529
timestamp 0
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_541
timestamp 0
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_553
timestamp 0
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_559
timestamp 0
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_561
timestamp 0
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_573
timestamp 0
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_585
timestamp 0
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_597
timestamp 0
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_609
timestamp 0
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_615
timestamp 0
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_617
timestamp 0
transform 1 0 57868 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_621
timestamp 0
transform 1 0 58236 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 0
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 0
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 0
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 0
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 0
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 0
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 0
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 0
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 0
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 0
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 0
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 0
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 0
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 0
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 0
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 0
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 0
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 0
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 0
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 0
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 0
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 0
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 0
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 0
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 0
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 0
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 0
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 0
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 0
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 0
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 0
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 0
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 0
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 0
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 0
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 0
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 0
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 0
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 0
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 0
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 0
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 0
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 0
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_457
timestamp 0
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_469
timestamp 0
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_475
timestamp 0
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_477
timestamp 0
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_489
timestamp 0
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_501
timestamp 0
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_513
timestamp 0
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 0
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 0
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 0
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_545
timestamp 0
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_557
timestamp 0
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_569
timestamp 0
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_581
timestamp 0
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_587
timestamp 0
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_589
timestamp 0
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_601
timestamp 0
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_613
timestamp 0
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 0
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 0
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 0
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 0
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 0
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 0
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 0
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 0
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 0
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 0
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 0
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 0
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 0
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 0
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 0
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 0
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 0
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 0
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 0
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 0
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 0
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 0
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 0
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 0
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 0
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 0
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 0
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 0
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 0
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 0
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 0
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 0
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 0
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 0
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 0
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 0
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 0
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 0
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 0
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 0
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 0
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 0
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_461
timestamp 0
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_473
timestamp 0
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_485
timestamp 0
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_497
timestamp 0
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 0
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_505
timestamp 0
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_517
timestamp 0
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_529
timestamp 0
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_541
timestamp 0
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_553
timestamp 0
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_559
timestamp 0
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_561
timestamp 0
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_573
timestamp 0
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_585
timestamp 0
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_597
timestamp 0
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_609
timestamp 0
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_615
timestamp 0
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_617
timestamp 0
transform 1 0 57868 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_621
timestamp 0
transform 1 0 58236 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 0
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 0
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 0
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 0
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 0
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 0
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 0
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 0
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 0
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 0
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 0
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 0
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 0
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 0
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 0
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 0
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 0
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 0
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 0
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 0
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 0
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 0
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 0
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 0
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 0
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 0
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 0
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 0
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 0
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 0
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 0
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 0
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 0
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 0
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 0
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 0
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 0
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 0
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 0
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 0
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 0
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 0
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 0
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_457
timestamp 0
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_469
timestamp 0
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_475
timestamp 0
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_477
timestamp 0
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_489
timestamp 0
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_501
timestamp 0
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_513
timestamp 0
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_525
timestamp 0
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_531
timestamp 0
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_533
timestamp 0
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_545
timestamp 0
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_557
timestamp 0
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_569
timestamp 0
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_581
timestamp 0
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_587
timestamp 0
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 0
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 0
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_613
timestamp 0
transform 1 0 57500 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_621
timestamp 0
transform 1 0 58236 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 0
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 0
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 0
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 0
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 0
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 0
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 0
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 0
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 0
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 0
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 0
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 0
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 0
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 0
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 0
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 0
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 0
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 0
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 0
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 0
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 0
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 0
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 0
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 0
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 0
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 0
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 0
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 0
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 0
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 0
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 0
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 0
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 0
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 0
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 0
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 0
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 0
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 0
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 0
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 0
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 0
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 0
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 0
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_461
timestamp 0
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_473
timestamp 0
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_485
timestamp 0
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_497
timestamp 0
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 0
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_505
timestamp 0
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_517
timestamp 0
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_529
timestamp 0
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_541
timestamp 0
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_553
timestamp 0
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 0
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_561
timestamp 0
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_573
timestamp 0
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_585
timestamp 0
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_597
timestamp 0
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_609
timestamp 0
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_615
timestamp 0
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_617
timestamp 0
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 0
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 0
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 0
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 0
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 0
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 0
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 0
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 0
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 0
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 0
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 0
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 0
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 0
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 0
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 0
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 0
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 0
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 0
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 0
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 0
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 0
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 0
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 0
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 0
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 0
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 0
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 0
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 0
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 0
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 0
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 0
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 0
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 0
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 0
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 0
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 0
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 0
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_401
timestamp 0
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_413
timestamp 0
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 0
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 0
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 0
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_445
timestamp 0
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_457
timestamp 0
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_469
timestamp 0
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_475
timestamp 0
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 0
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 0
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_501
timestamp 0
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_513
timestamp 0
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_525
timestamp 0
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_531
timestamp 0
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 0
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_545
timestamp 0
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_557
timestamp 0
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_569
timestamp 0
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_581
timestamp 0
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_587
timestamp 0
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 0
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 0
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_613
timestamp 0
transform 1 0 57500 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_621
timestamp 0
transform 1 0 58236 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 0
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 0
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 0
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 0
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 0
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 0
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 0
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 0
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 0
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 0
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 0
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 0
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 0
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 0
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 0
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 0
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 0
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 0
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 0
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 0
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 0
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 0
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 0
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 0
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 0
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 0
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 0
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 0
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 0
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 0
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 0
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 0
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 0
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 0
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 0
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 0
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 0
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 0
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 0
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 0
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 0
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 0
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 0
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 0
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 0
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_429
timestamp 0
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_441
timestamp 0
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_447
timestamp 0
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_449
timestamp 0
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_461
timestamp 0
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_473
timestamp 0
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_485
timestamp 0
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_497
timestamp 0
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_503
timestamp 0
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_505
timestamp 0
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_517
timestamp 0
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_529
timestamp 0
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_541
timestamp 0
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_553
timestamp 0
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_559
timestamp 0
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_561
timestamp 0
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_573
timestamp 0
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_585
timestamp 0
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_597
timestamp 0
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_609
timestamp 0
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_615
timestamp 0
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_617
timestamp 0
transform 1 0 57868 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_621
timestamp 0
transform 1 0 58236 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 0
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 0
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 0
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 0
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 0
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 0
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 0
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 0
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 0
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 0
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 0
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 0
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 0
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 0
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 0
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 0
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 0
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 0
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 0
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 0
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 0
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 0
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 0
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 0
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 0
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 0
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 0
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 0
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 0
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 0
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 0
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 0
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 0
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 0
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 0
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 0
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 0
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 0
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 0
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 0
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 0
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 0
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_401
timestamp 0
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_413
timestamp 0
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 0
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 0
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_433
timestamp 0
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_445
timestamp 0
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_457
timestamp 0
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_469
timestamp 0
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_475
timestamp 0
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_477
timestamp 0
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_489
timestamp 0
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_501
timestamp 0
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_513
timestamp 0
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_525
timestamp 0
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_531
timestamp 0
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_533
timestamp 0
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_545
timestamp 0
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_557
timestamp 0
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_569
timestamp 0
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_581
timestamp 0
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_587
timestamp 0
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_589
timestamp 0
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_601
timestamp 0
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_613
timestamp 0
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 0
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 0
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 0
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 0
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 0
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 0
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 0
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 0
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 0
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 0
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 0
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 0
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 0
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 0
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 0
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 0
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 0
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 0
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 0
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 0
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 0
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 0
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 0
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 0
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 0
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 0
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 0
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 0
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 0
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 0
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 0
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 0
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 0
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 0
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 0
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 0
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 0
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 0
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 0
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 0
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 0
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 0
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 0
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_405
timestamp 0
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_417
timestamp 0
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_429
timestamp 0
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_441
timestamp 0
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_447
timestamp 0
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_449
timestamp 0
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_461
timestamp 0
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_473
timestamp 0
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_485
timestamp 0
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_497
timestamp 0
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_503
timestamp 0
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_505
timestamp 0
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_517
timestamp 0
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_529
timestamp 0
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_541
timestamp 0
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_553
timestamp 0
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_559
timestamp 0
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_561
timestamp 0
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_573
timestamp 0
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_585
timestamp 0
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_597
timestamp 0
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_609
timestamp 0
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_615
timestamp 0
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_617
timestamp 0
transform 1 0 57868 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_621
timestamp 0
transform 1 0 58236 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 0
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 0
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 0
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 0
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 0
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 0
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 0
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 0
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 0
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 0
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 0
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 0
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 0
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 0
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 0
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 0
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 0
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 0
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 0
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 0
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 0
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 0
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 0
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 0
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 0
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 0
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 0
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 0
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 0
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 0
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 0
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 0
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 0
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 0
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 0
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 0
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 0
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 0
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 0
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 0
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 0
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 0
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_401
timestamp 0
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_413
timestamp 0
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_419
timestamp 0
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 0
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 0
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_445
timestamp 0
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_457
timestamp 0
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_469
timestamp 0
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_475
timestamp 0
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_477
timestamp 0
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_489
timestamp 0
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_501
timestamp 0
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_513
timestamp 0
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_525
timestamp 0
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_531
timestamp 0
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_533
timestamp 0
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_545
timestamp 0
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_557
timestamp 0
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_569
timestamp 0
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_581
timestamp 0
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_587
timestamp 0
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_589
timestamp 0
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_601
timestamp 0
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_613
timestamp 0
transform 1 0 57500 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_621
timestamp 0
transform 1 0 58236 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 0
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 0
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 0
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 0
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 0
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 0
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 0
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 0
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 0
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 0
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 0
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 0
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 0
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 0
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 0
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 0
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 0
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 0
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 0
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 0
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 0
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 0
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 0
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 0
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 0
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 0
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 0
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 0
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 0
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 0
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 0
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 0
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 0
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 0
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 0
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 0
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 0
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 0
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 0
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 0
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 0
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 0
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 0
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 0
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 0
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_429
timestamp 0
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_441
timestamp 0
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_447
timestamp 0
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_449
timestamp 0
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_461
timestamp 0
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_473
timestamp 0
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_485
timestamp 0
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_497
timestamp 0
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_503
timestamp 0
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_505
timestamp 0
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_517
timestamp 0
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_529
timestamp 0
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_541
timestamp 0
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_553
timestamp 0
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_559
timestamp 0
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_561
timestamp 0
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_573
timestamp 0
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_585
timestamp 0
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_597
timestamp 0
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_609
timestamp 0
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_615
timestamp 0
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_617
timestamp 0
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 0
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 0
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 0
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 0
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 0
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 0
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 0
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 0
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 0
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 0
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 0
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 0
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 0
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 0
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 0
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 0
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 0
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 0
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 0
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 0
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 0
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 0
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 0
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 0
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 0
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 0
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 0
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 0
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 0
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 0
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 0
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 0
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 0
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 0
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 0
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 0
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 0
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 0
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 0
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 0
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 0
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 0
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_401
timestamp 0
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_413
timestamp 0
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 0
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 0
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_433
timestamp 0
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_445
timestamp 0
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_457
timestamp 0
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_469
timestamp 0
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_475
timestamp 0
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_477
timestamp 0
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_489
timestamp 0
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_501
timestamp 0
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_513
timestamp 0
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_525
timestamp 0
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_531
timestamp 0
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_533
timestamp 0
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_545
timestamp 0
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_557
timestamp 0
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_569
timestamp 0
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_581
timestamp 0
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_587
timestamp 0
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_589
timestamp 0
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_601
timestamp 0
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_613
timestamp 0
transform 1 0 57500 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_621
timestamp 0
transform 1 0 58236 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 0
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 0
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 0
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 0
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 0
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 0
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 0
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 0
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 0
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 0
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 0
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 0
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 0
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 0
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 0
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 0
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 0
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 0
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 0
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 0
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 0
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 0
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 0
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 0
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 0
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 0
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 0
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 0
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 0
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 0
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 0
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 0
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 0
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 0
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 0
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 0
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 0
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 0
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 0
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 0
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 0
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 0
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 0
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 0
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 0
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_429
timestamp 0
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_441
timestamp 0
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_447
timestamp 0
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 0
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_461
timestamp 0
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_473
timestamp 0
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_485
timestamp 0
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_497
timestamp 0
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_503
timestamp 0
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_505
timestamp 0
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_517
timestamp 0
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_529
timestamp 0
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_541
timestamp 0
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_553
timestamp 0
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_559
timestamp 0
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_561
timestamp 0
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_573
timestamp 0
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_585
timestamp 0
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_597
timestamp 0
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_609
timestamp 0
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_615
timestamp 0
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_617
timestamp 0
transform 1 0 57868 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_621
timestamp 0
transform 1 0 58236 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 0
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 0
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 0
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 0
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 0
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 0
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 0
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 0
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 0
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 0
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 0
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 0
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 0
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 0
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 0
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 0
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 0
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 0
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 0
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 0
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 0
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 0
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 0
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 0
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 0
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 0
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 0
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 0
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 0
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 0
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 0
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 0
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 0
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 0
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 0
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 0
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 0
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 0
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 0
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 0
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 0
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 0
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_401
timestamp 0
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_413
timestamp 0
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 0
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 0
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 0
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 0
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_457
timestamp 0
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_469
timestamp 0
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_475
timestamp 0
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_477
timestamp 0
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_489
timestamp 0
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_501
timestamp 0
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_513
timestamp 0
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_525
timestamp 0
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_531
timestamp 0
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_533
timestamp 0
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_545
timestamp 0
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_557
timestamp 0
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_569
timestamp 0
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_581
timestamp 0
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_587
timestamp 0
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_589
timestamp 0
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_601
timestamp 0
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_613
timestamp 0
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 0
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 0
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 0
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 0
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 0
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 0
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 0
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 0
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 0
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 0
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 0
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 0
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 0
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 0
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 0
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 0
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 0
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 0
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 0
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 0
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 0
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 0
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 0
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 0
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 0
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 0
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 0
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 0
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 0
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 0
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 0
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 0
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 0
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 0
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 0
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 0
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 0
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 0
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 0
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 0
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 0
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 0
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 0
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 0
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 0
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 0
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_441
timestamp 0
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_447
timestamp 0
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 0
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_461
timestamp 0
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_473
timestamp 0
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_485
timestamp 0
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_497
timestamp 0
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_503
timestamp 0
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_505
timestamp 0
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_517
timestamp 0
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_529
timestamp 0
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_541
timestamp 0
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_553
timestamp 0
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_559
timestamp 0
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_561
timestamp 0
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_573
timestamp 0
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_585
timestamp 0
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_597
timestamp 0
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_609
timestamp 0
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_615
timestamp 0
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_617
timestamp 0
transform 1 0 57868 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_621
timestamp 0
transform 1 0 58236 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 0
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 0
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 0
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 0
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 0
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 0
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 0
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 0
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 0
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 0
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 0
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 0
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 0
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 0
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 0
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 0
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 0
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 0
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 0
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 0
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 0
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 0
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 0
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 0
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 0
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 0
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 0
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 0
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 0
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 0
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 0
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 0
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 0
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 0
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 0
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 0
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 0
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 0
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 0
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 0
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 0
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 0
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 0
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 0
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 0
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_421
timestamp 0
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_433
timestamp 0
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_445
timestamp 0
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_457
timestamp 0
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_469
timestamp 0
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_475
timestamp 0
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_477
timestamp 0
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_489
timestamp 0
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_501
timestamp 0
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_513
timestamp 0
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_525
timestamp 0
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_531
timestamp 0
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_533
timestamp 0
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_545
timestamp 0
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_557
timestamp 0
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_569
timestamp 0
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_581
timestamp 0
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_587
timestamp 0
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_589
timestamp 0
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_601
timestamp 0
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_613
timestamp 0
transform 1 0 57500 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_621
timestamp 0
transform 1 0 58236 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 0
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 0
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 0
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 0
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 0
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 0
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 0
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 0
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 0
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 0
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 0
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 0
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 0
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 0
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 0
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 0
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 0
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 0
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 0
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 0
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 0
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 0
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 0
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 0
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 0
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 0
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 0
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 0
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 0
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 0
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 0
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 0
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 0
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 0
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 0
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 0
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 0
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 0
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 0
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 0
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 0
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 0
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 0
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 0
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 0
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_429
timestamp 0
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_441
timestamp 0
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 0
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_449
timestamp 0
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_461
timestamp 0
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_473
timestamp 0
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_485
timestamp 0
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_497
timestamp 0
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_503
timestamp 0
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_505
timestamp 0
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_517
timestamp 0
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_529
timestamp 0
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_541
timestamp 0
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_553
timestamp 0
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_559
timestamp 0
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_561
timestamp 0
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_573
timestamp 0
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_585
timestamp 0
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_597
timestamp 0
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_609
timestamp 0
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_615
timestamp 0
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_617
timestamp 0
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 0
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 0
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 0
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 0
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 0
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 0
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 0
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 0
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 0
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 0
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 0
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 0
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 0
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 0
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 0
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 0
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 0
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 0
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 0
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 0
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 0
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 0
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 0
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 0
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 0
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 0
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 0
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 0
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 0
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 0
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 0
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 0
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 0
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 0
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 0
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 0
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 0
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 0
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 0
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 0
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 0
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 0
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 0
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 0
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 0
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 0
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_433
timestamp 0
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_445
timestamp 0
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_457
timestamp 0
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_469
timestamp 0
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_475
timestamp 0
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_477
timestamp 0
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_489
timestamp 0
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_501
timestamp 0
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_513
timestamp 0
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_525
timestamp 0
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_531
timestamp 0
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_533
timestamp 0
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_545
timestamp 0
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_557
timestamp 0
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_569
timestamp 0
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_581
timestamp 0
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_587
timestamp 0
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_589
timestamp 0
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_601
timestamp 0
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_613
timestamp 0
transform 1 0 57500 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_621
timestamp 0
transform 1 0 58236 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 0
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 0
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 0
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 0
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 0
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 0
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 0
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 0
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 0
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 0
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 0
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 0
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 0
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 0
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 0
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 0
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 0
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 0
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 0
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 0
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 0
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 0
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 0
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 0
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 0
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 0
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 0
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 0
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 0
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 0
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 0
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 0
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 0
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 0
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 0
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 0
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 0
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 0
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 0
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 0
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 0
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 0
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 0
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 0
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 0
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 0
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 0
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 0
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 0
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_461
timestamp 0
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_473
timestamp 0
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_485
timestamp 0
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_497
timestamp 0
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_503
timestamp 0
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_505
timestamp 0
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_517
timestamp 0
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_529
timestamp 0
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_541
timestamp 0
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_553
timestamp 0
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_559
timestamp 0
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_561
timestamp 0
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_573
timestamp 0
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_585
timestamp 0
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_597
timestamp 0
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_609
timestamp 0
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_615
timestamp 0
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_617
timestamp 0
transform 1 0 57868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_621
timestamp 0
transform 1 0 58236 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 0
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 0
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 0
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 0
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 0
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 0
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 0
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 0
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 0
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 0
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 0
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 0
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 0
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 0
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 0
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 0
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 0
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 0
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 0
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 0
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 0
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 0
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 0
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 0
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 0
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 0
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 0
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 0
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 0
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 0
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 0
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 0
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 0
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 0
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 0
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 0
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 0
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 0
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 0
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 0
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 0
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 0
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 0
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 0
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 0
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 0
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 0
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 0
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_457
timestamp 0
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_469
timestamp 0
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_475
timestamp 0
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_477
timestamp 0
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_489
timestamp 0
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_501
timestamp 0
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_513
timestamp 0
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_525
timestamp 0
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_531
timestamp 0
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_533
timestamp 0
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_545
timestamp 0
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_557
timestamp 0
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_569
timestamp 0
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_581
timestamp 0
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_587
timestamp 0
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_589
timestamp 0
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_601
timestamp 0
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_613
timestamp 0
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 0
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 0
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 0
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 0
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 0
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 0
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 0
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 0
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 0
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 0
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 0
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 0
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 0
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 0
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 0
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 0
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 0
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 0
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 0
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 0
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 0
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 0
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 0
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 0
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 0
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 0
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 0
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 0
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 0
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 0
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 0
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 0
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 0
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 0
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 0
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 0
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 0
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 0
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 0
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 0
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 0
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 0
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 0
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 0
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 0
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 0
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 0
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 0
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 0
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 0
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_473
timestamp 0
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_485
timestamp 0
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_497
timestamp 0
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_503
timestamp 0
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_505
timestamp 0
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_517
timestamp 0
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_529
timestamp 0
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_541
timestamp 0
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_553
timestamp 0
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_559
timestamp 0
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_561
timestamp 0
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_573
timestamp 0
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_585
timestamp 0
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_597
timestamp 0
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_609
timestamp 0
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_615
timestamp 0
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_617
timestamp 0
transform 1 0 57868 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_621
timestamp 0
transform 1 0 58236 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 0
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 0
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 0
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 0
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 0
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 0
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 0
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 0
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 0
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 0
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 0
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 0
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 0
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 0
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 0
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 0
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 0
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 0
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 0
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 0
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 0
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 0
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 0
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 0
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 0
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 0
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 0
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 0
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 0
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 0
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 0
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 0
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 0
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 0
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 0
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 0
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 0
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 0
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 0
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 0
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 0
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 0
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 0
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 0
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 0
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 0
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 0
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_445
timestamp 0
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_457
timestamp 0
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_469
timestamp 0
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_475
timestamp 0
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_477
timestamp 0
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_489
timestamp 0
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_501
timestamp 0
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_513
timestamp 0
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_525
timestamp 0
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_531
timestamp 0
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_533
timestamp 0
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_545
timestamp 0
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_557
timestamp 0
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_569
timestamp 0
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_581
timestamp 0
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_587
timestamp 0
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_589
timestamp 0
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_601
timestamp 0
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_613
timestamp 0
transform 1 0 57500 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_621
timestamp 0
transform 1 0 58236 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 0
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 0
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 0
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 0
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 0
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 0
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 0
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 0
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 0
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 0
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 0
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 0
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 0
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 0
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 0
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 0
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 0
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 0
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 0
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 0
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 0
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 0
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 0
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 0
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 0
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 0
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 0
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 0
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 0
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 0
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 0
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 0
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 0
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 0
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 0
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 0
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 0
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 0
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 0
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 0
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 0
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 0
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 0
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 0
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 0
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_429
timestamp 0
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_441
timestamp 0
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_447
timestamp 0
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_449
timestamp 0
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_461
timestamp 0
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_473
timestamp 0
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_485
timestamp 0
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_497
timestamp 0
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_503
timestamp 0
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_505
timestamp 0
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_517
timestamp 0
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_529
timestamp 0
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_541
timestamp 0
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_553
timestamp 0
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_559
timestamp 0
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_561
timestamp 0
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_573
timestamp 0
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_585
timestamp 0
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_597
timestamp 0
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_609
timestamp 0
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_615
timestamp 0
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_617
timestamp 0
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 0
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 0
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 0
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 0
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 0
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 0
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 0
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 0
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 0
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 0
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 0
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 0
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 0
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 0
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 0
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 0
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 0
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 0
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_177
timestamp 0
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_189
timestamp 0
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_195
timestamp 0
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 0
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 0
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 0
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 0
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 0
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 0
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 0
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 0
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 0
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 0
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 0
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 0
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 0
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 0
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 0
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 0
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 0
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 0
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 0
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 0
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 0
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 0
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 0
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 0
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 0
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 0
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_445
timestamp 0
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_457
timestamp 0
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_469
timestamp 0
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_475
timestamp 0
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_477
timestamp 0
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_489
timestamp 0
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_501
timestamp 0
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_513
timestamp 0
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_525
timestamp 0
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_531
timestamp 0
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_533
timestamp 0
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_545
timestamp 0
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_557
timestamp 0
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_569
timestamp 0
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_581
timestamp 0
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_587
timestamp 0
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_589
timestamp 0
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_601
timestamp 0
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_613
timestamp 0
transform 1 0 57500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_621
timestamp 0
transform 1 0 58236 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 0
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 0
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 0
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 0
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 0
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 0
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 0
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 0
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 0
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 0
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 0
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 0
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 0
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 0
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 0
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 0
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 0
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 0
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 0
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 0
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 0
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 0
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 0
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 0
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 0
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 0
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 0
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_261
timestamp 0
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_273
timestamp 0
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 0
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 0
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 0
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 0
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 0
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 0
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 0
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 0
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 0
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 0
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 0
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 0
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 0
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 0
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 0
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 0
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_429
timestamp 0
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_441
timestamp 0
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_447
timestamp 0
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_449
timestamp 0
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_461
timestamp 0
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_473
timestamp 0
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_485
timestamp 0
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_497
timestamp 0
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_503
timestamp 0
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_505
timestamp 0
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_517
timestamp 0
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_529
timestamp 0
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_541
timestamp 0
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_553
timestamp 0
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_559
timestamp 0
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_561
timestamp 0
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_573
timestamp 0
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_585
timestamp 0
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_597
timestamp 0
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_609
timestamp 0
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_615
timestamp 0
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_617
timestamp 0
transform 1 0 57868 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_621
timestamp 0
transform 1 0 58236 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 0
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 0
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 0
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 0
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 0
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 0
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 0
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 0
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 0
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 0
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 0
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 0
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 0
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 0
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 0
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 0
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 0
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 0
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 0
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 0
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 0
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 0
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_209
timestamp 0
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_221
timestamp 0
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_233
timestamp 0
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 0
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 0
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 0
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 0
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 0
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 0
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 0
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 0
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 0
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 0
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 0
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 0
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 0
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 0
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 0
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 0
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 0
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 0
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 0
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 0
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 0
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_433
timestamp 0
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_445
timestamp 0
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_457
timestamp 0
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_469
timestamp 0
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_475
timestamp 0
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_477
timestamp 0
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_489
timestamp 0
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_501
timestamp 0
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_513
timestamp 0
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_525
timestamp 0
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_531
timestamp 0
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_533
timestamp 0
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_545
timestamp 0
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_557
timestamp 0
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_569
timestamp 0
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_581
timestamp 0
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_587
timestamp 0
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_589
timestamp 0
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_601
timestamp 0
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_613
timestamp 0
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 0
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 0
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 0
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 0
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 0
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 0
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 0
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 0
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 0
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 0
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 0
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 0
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 0
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 0
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 0
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 0
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 0
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 0
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 0
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 0
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 0
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 0
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 0
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 0
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 0
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_237
timestamp 0
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_249
timestamp 0
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 0
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 0
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 0
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 0
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 0
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 0
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 0
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 0
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 0
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 0
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 0
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 0
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 0
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 0
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 0
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 0
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 0
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 0
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_429
timestamp 0
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_441
timestamp 0
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_447
timestamp 0
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_449
timestamp 0
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_461
timestamp 0
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_473
timestamp 0
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_485
timestamp 0
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_497
timestamp 0
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_503
timestamp 0
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_505
timestamp 0
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_517
timestamp 0
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_529
timestamp 0
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_541
timestamp 0
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_553
timestamp 0
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_559
timestamp 0
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_561
timestamp 0
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_573
timestamp 0
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_585
timestamp 0
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_597
timestamp 0
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_609
timestamp 0
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_615
timestamp 0
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_617
timestamp 0
transform 1 0 57868 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_621
timestamp 0
transform 1 0 58236 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 0
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 0
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 0
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 0
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 0
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 0
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 0
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 0
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 0
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 0
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 0
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 0
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 0
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 0
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 0
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 0
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 0
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 0
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 0
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 0
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 0
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 0
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 0
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 0
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_233
timestamp 0
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_245
timestamp 0
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 0
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 0
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 0
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_277
timestamp 0
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 0
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 0
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 0
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 0
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 0
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_333
timestamp 0
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 0
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 0
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 0
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 0
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 0
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 0
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 0
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 0
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 0
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 0
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_433
timestamp 0
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_445
timestamp 0
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_457
timestamp 0
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_469
timestamp 0
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_475
timestamp 0
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_477
timestamp 0
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_489
timestamp 0
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_501
timestamp 0
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_513
timestamp 0
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_525
timestamp 0
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_531
timestamp 0
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_533
timestamp 0
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_545
timestamp 0
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_557
timestamp 0
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_569
timestamp 0
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_581
timestamp 0
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_587
timestamp 0
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_589
timestamp 0
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_601
timestamp 0
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_613
timestamp 0
transform 1 0 57500 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_621
timestamp 0
transform 1 0 58236 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 0
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 0
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 0
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 0
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 0
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 0
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 0
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 0
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 0
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 0
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 0
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 0
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 0
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 0
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 0
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 0
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 0
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 0
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 0
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 0
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 0
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_205
timestamp 0
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_217
timestamp 0
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 0
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 0
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 0
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 0
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 0
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 0
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 0
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 0
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 0
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 0
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 0
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 0
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 0
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 0
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 0
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 0
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 0
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 0
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 0
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 0
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 0
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 0
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_429
timestamp 0
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_441
timestamp 0
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_447
timestamp 0
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_449
timestamp 0
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_461
timestamp 0
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_473
timestamp 0
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_485
timestamp 0
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_497
timestamp 0
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_503
timestamp 0
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_505
timestamp 0
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_517
timestamp 0
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_529
timestamp 0
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_541
timestamp 0
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_553
timestamp 0
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_559
timestamp 0
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_561
timestamp 0
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_573
timestamp 0
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_585
timestamp 0
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_597
timestamp 0
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_609
timestamp 0
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_615
timestamp 0
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_617
timestamp 0
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 0
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 0
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 0
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 0
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 0
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 0
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 0
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 0
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 0
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 0
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 0
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 0
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 0
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 0
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 0
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 0
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 0
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 0
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 0
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 0
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 0
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 0
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 0
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 0
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 0
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 0
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 0
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 0
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 0
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 0
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 0
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 0
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 0
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 0
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 0
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 0
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 0
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 0
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 0
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 0
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 0
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 0
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 0
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 0
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 0
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 0
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_433
timestamp 0
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_445
timestamp 0
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_457
timestamp 0
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_469
timestamp 0
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_475
timestamp 0
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_477
timestamp 0
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_489
timestamp 0
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_501
timestamp 0
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_513
timestamp 0
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_525
timestamp 0
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_531
timestamp 0
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_533
timestamp 0
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_545
timestamp 0
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_557
timestamp 0
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_569
timestamp 0
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_581
timestamp 0
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_587
timestamp 0
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_589
timestamp 0
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_601
timestamp 0
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_613
timestamp 0
transform 1 0 57500 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_621
timestamp 0
transform 1 0 58236 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 0
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 0
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 0
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 0
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 0
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 0
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 0
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 0
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 0
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 0
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 0
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 0
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 0
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 0
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 0
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 0
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 0
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 0
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 0
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 0
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 0
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 0
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 0
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 0
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 0
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 0
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 0
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_261
timestamp 0
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 0
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 0
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 0
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 0
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 0
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 0
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 0
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 0
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 0
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 0
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 0
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 0
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 0
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 0
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 0
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 0
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 0
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 0
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_441
timestamp 0
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 0
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_449
timestamp 0
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_461
timestamp 0
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_473
timestamp 0
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_485
timestamp 0
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_497
timestamp 0
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_503
timestamp 0
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_505
timestamp 0
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_517
timestamp 0
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_529
timestamp 0
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_541
timestamp 0
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_553
timestamp 0
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_559
timestamp 0
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_561
timestamp 0
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_573
timestamp 0
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_585
timestamp 0
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_597
timestamp 0
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_609
timestamp 0
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_615
timestamp 0
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_617
timestamp 0
transform 1 0 57868 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_621
timestamp 0
transform 1 0 58236 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 0
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 0
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 0
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 0
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 0
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 0
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 0
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 0
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 0
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 0
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 0
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 0
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 0
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 0
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 0
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 0
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 0
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 0
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 0
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 0
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 0
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 0
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 0
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 0
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 0
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 0
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 0
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 0
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 0
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 0
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 0
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_301
timestamp 0
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 0
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 0
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 0
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 0
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 0
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 0
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 0
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 0
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 0
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 0
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 0
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 0
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 0
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 0
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_433
timestamp 0
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_445
timestamp 0
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_457
timestamp 0
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_469
timestamp 0
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_475
timestamp 0
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_477
timestamp 0
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_489
timestamp 0
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_501
timestamp 0
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_513
timestamp 0
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_525
timestamp 0
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_531
timestamp 0
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_533
timestamp 0
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_545
timestamp 0
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_557
timestamp 0
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_569
timestamp 0
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_581
timestamp 0
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_587
timestamp 0
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_589
timestamp 0
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_601
timestamp 0
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_613
timestamp 0
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 0
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 0
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 0
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 0
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 0
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 0
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 0
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 0
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 0
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 0
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 0
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 0
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 0
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 0
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 0
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 0
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 0
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 0
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 0
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 0
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_193
timestamp 0
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_205
timestamp 0
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_217
timestamp 0
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 0
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 0
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 0
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_249
timestamp 0
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_261
timestamp 0
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_273
timestamp 0
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_279
timestamp 0
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 0
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 0
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_305
timestamp 0
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_317
timestamp 0
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_329
timestamp 0
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 0
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_337
timestamp 0
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_349
timestamp 0
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_361
timestamp 0
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_373
timestamp 0
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_385
timestamp 0
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 0
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 0
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 0
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 0
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_429
timestamp 0
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_441
timestamp 0
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_447
timestamp 0
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_449
timestamp 0
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_461
timestamp 0
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_473
timestamp 0
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_485
timestamp 0
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_497
timestamp 0
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_503
timestamp 0
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_505
timestamp 0
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_517
timestamp 0
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_529
timestamp 0
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_541
timestamp 0
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_553
timestamp 0
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_559
timestamp 0
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_561
timestamp 0
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_573
timestamp 0
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_585
timestamp 0
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_597
timestamp 0
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_609
timestamp 0
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_615
timestamp 0
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_617
timestamp 0
transform 1 0 57868 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_621
timestamp 0
transform 1 0 58236 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 0
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 0
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 0
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 0
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 0
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 0
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 0
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 0
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 0
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 0
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 0
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 0
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 0
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 0
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 0
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 0
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 0
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 0
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 0
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 0
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 0
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_197
timestamp 0
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_209
timestamp 0
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_221
timestamp 0
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_233
timestamp 0
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_245
timestamp 0
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_251
timestamp 0
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_253
timestamp 0
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_265
timestamp 0
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_277
timestamp 0
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_289
timestamp 0
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_301
timestamp 0
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_307
timestamp 0
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 0
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 0
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 0
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 0
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 0
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 0
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_365
timestamp 0
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_377
timestamp 0
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_389
timestamp 0
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_401
timestamp 0
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_413
timestamp 0
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_419
timestamp 0
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_421
timestamp 0
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_433
timestamp 0
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_445
timestamp 0
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_457
timestamp 0
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_469
timestamp 0
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_475
timestamp 0
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_477
timestamp 0
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_489
timestamp 0
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_501
timestamp 0
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_513
timestamp 0
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_525
timestamp 0
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_531
timestamp 0
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_533
timestamp 0
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_545
timestamp 0
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_557
timestamp 0
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_569
timestamp 0
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_581
timestamp 0
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_587
timestamp 0
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_589
timestamp 0
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_601
timestamp 0
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_613
timestamp 0
transform 1 0 57500 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_621
timestamp 0
transform 1 0 58236 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 0
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 0
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 0
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 0
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 0
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 0
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 0
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 0
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 0
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 0
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 0
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 0
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 0
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 0
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 0
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 0
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 0
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 0
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 0
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_181
timestamp 0
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_193
timestamp 0
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_205
timestamp 0
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 0
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 0
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 0
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 0
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 0
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 0
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 0
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 0
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 0
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_293
timestamp 0
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_305
timestamp 0
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_317
timestamp 0
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 0
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 0
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 0
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_349
timestamp 0
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_361
timestamp 0
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_373
timestamp 0
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_385
timestamp 0
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_391
timestamp 0
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 0
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 0
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 0
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_429
timestamp 0
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_441
timestamp 0
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_447
timestamp 0
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_449
timestamp 0
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_461
timestamp 0
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_473
timestamp 0
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_485
timestamp 0
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_497
timestamp 0
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_503
timestamp 0
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_505
timestamp 0
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_517
timestamp 0
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_529
timestamp 0
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_541
timestamp 0
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_553
timestamp 0
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_559
timestamp 0
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_561
timestamp 0
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_573
timestamp 0
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_585
timestamp 0
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_597
timestamp 0
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_609
timestamp 0
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_615
timestamp 0
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_617
timestamp 0
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 0
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 0
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 0
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 0
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 0
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 0
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 0
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 0
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 0
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 0
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 0
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 0
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 0
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 0
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 0
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 0
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 0
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 0
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 0
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_189
timestamp 0
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 0
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_197
timestamp 0
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_209
timestamp 0
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_221
timestamp 0
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_233
timestamp 0
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_245
timestamp 0
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 0
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_253
timestamp 0
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_265
timestamp 0
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_277
timestamp 0
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_289
timestamp 0
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_301
timestamp 0
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_307
timestamp 0
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 0
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_321
timestamp 0
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_333
timestamp 0
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_345
timestamp 0
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 0
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 0
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 0
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 0
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 0
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 0
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 0
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 0
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_421
timestamp 0
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_433
timestamp 0
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_445
timestamp 0
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_457
timestamp 0
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_469
timestamp 0
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_475
timestamp 0
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_477
timestamp 0
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_489
timestamp 0
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_501
timestamp 0
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_513
timestamp 0
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_525
timestamp 0
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_531
timestamp 0
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_533
timestamp 0
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_545
timestamp 0
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_557
timestamp 0
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_569
timestamp 0
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_581
timestamp 0
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_587
timestamp 0
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_589
timestamp 0
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_601
timestamp 0
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_613
timestamp 0
transform 1 0 57500 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_621
timestamp 0
transform 1 0 58236 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 0
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 0
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 0
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 0
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 0
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 0
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 0
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 0
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 0
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 0
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 0
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 0
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 0
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 0
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 0
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 0
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 0
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 0
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 0
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_181
timestamp 0
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_193
timestamp 0
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_205
timestamp 0
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_217
timestamp 0
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 0
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 0
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 0
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 0
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 0
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 0
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 0
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 0
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 0
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 0
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 0
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 0
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 0
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 0
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 0
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 0
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 0
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 0
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 0
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 0
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 0
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 0
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_429
timestamp 0
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_441
timestamp 0
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_447
timestamp 0
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_449
timestamp 0
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_461
timestamp 0
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_473
timestamp 0
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_485
timestamp 0
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_497
timestamp 0
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_503
timestamp 0
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_505
timestamp 0
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_517
timestamp 0
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_529
timestamp 0
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_541
timestamp 0
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_553
timestamp 0
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_559
timestamp 0
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_561
timestamp 0
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_573
timestamp 0
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_585
timestamp 0
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_597
timestamp 0
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_609
timestamp 0
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_615
timestamp 0
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_617
timestamp 0
transform 1 0 57868 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_621
timestamp 0
transform 1 0 58236 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 0
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 0
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 0
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 0
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 0
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 0
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 0
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 0
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 0
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 0
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 0
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 0
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 0
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 0
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 0
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 0
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 0
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 0
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 0
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_189
timestamp 0
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 0
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_197
timestamp 0
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_209
timestamp 0
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_221
timestamp 0
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_233
timestamp 0
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_245
timestamp 0
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_251
timestamp 0
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 0
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 0
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 0
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 0
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 0
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 0
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 0
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 0
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_333
timestamp 0
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_345
timestamp 0
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_357
timestamp 0
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_363
timestamp 0
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 0
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 0
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 0
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 0
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 0
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 0
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_421
timestamp 0
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_433
timestamp 0
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_445
timestamp 0
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_457
timestamp 0
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_469
timestamp 0
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_475
timestamp 0
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_477
timestamp 0
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_489
timestamp 0
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_501
timestamp 0
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_513
timestamp 0
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_525
timestamp 0
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_531
timestamp 0
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_533
timestamp 0
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_545
timestamp 0
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_557
timestamp 0
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_569
timestamp 0
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_581
timestamp 0
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_587
timestamp 0
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_589
timestamp 0
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_601
timestamp 0
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_613
timestamp 0
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 0
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 0
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 0
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 0
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 0
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 0
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 0
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 0
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_81
timestamp 0
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_93
timestamp 0
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_105
timestamp 0
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_111
timestamp 0
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 0
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 0
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 0
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 0
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 0
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 0
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 0
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 0
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_193
timestamp 0
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_205
timestamp 0
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_217
timestamp 0
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_223
timestamp 0
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 0
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_237
timestamp 0
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_249
timestamp 0
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_261
timestamp 0
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_273
timestamp 0
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 0
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 0
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 0
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_305
timestamp 0
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_317
timestamp 0
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_329
timestamp 0
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_335
timestamp 0
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 0
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 0
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 0
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 0
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 0
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 0
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 0
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 0
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 0
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_429
timestamp 0
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_441
timestamp 0
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_447
timestamp 0
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_449
timestamp 0
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_461
timestamp 0
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_473
timestamp 0
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_485
timestamp 0
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_497
timestamp 0
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_503
timestamp 0
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_505
timestamp 0
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_517
timestamp 0
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_529
timestamp 0
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_541
timestamp 0
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_553
timestamp 0
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_559
timestamp 0
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_561
timestamp 0
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_573
timestamp 0
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_585
timestamp 0
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_597
timestamp 0
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_609
timestamp 0
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_615
timestamp 0
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_617
timestamp 0
transform 1 0 57868 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_621
timestamp 0
transform 1 0 58236 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_3
timestamp 0
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_15
timestamp 0
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 0
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 0
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 0
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 0
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 0
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 0
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 0
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 0
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 0
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 0
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 0
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 0
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 0
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_141
timestamp 0
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 0
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_165
timestamp 0
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_177
timestamp 0
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_189
timestamp 0
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_195
timestamp 0
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 0
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 0
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_221
timestamp 0
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_233
timestamp 0
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_245
timestamp 0
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 0
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 0
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_265
timestamp 0
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_277
timestamp 0
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_289
timestamp 0
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_301
timestamp 0
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 0
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 0
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 0
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_333
timestamp 0
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_345
timestamp 0
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_357
timestamp 0
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_363
timestamp 0
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 0
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 0
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_389
timestamp 0
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_401
timestamp 0
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_413
timestamp 0
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_419
timestamp 0
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_421
timestamp 0
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_433
timestamp 0
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_445
timestamp 0
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_457
timestamp 0
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_469
timestamp 0
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_475
timestamp 0
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_477
timestamp 0
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_489
timestamp 0
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_501
timestamp 0
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_513
timestamp 0
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_525
timestamp 0
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_531
timestamp 0
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_533
timestamp 0
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_545
timestamp 0
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_557
timestamp 0
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_569
timestamp 0
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_581
timestamp 0
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_587
timestamp 0
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_589
timestamp 0
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_601
timestamp 0
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_613
timestamp 0
transform 1 0 57500 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_621
timestamp 0
transform 1 0 58236 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_3
timestamp 0
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_15
timestamp 0
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_27
timestamp 0
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_39
timestamp 0
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_51
timestamp 0
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 0
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 0
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 0
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 0
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 0
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 0
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 0
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 0
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 0
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 0
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 0
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 0
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 0
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 0
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_181
timestamp 0
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_193
timestamp 0
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_205
timestamp 0
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_217
timestamp 0
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_223
timestamp 0
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_225
timestamp 0
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_237
timestamp 0
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_249
timestamp 0
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_261
timestamp 0
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_273
timestamp 0
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_279
timestamp 0
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_281
timestamp 0
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_293
timestamp 0
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_305
timestamp 0
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_317
timestamp 0
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_329
timestamp 0
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_335
timestamp 0
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_337
timestamp 0
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_349
timestamp 0
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_361
timestamp 0
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_373
timestamp 0
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_385
timestamp 0
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_391
timestamp 0
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_393
timestamp 0
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_405
timestamp 0
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_417
timestamp 0
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_429
timestamp 0
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_441
timestamp 0
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_447
timestamp 0
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_449
timestamp 0
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_461
timestamp 0
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_473
timestamp 0
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_485
timestamp 0
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_497
timestamp 0
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_503
timestamp 0
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_505
timestamp 0
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_517
timestamp 0
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_529
timestamp 0
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_541
timestamp 0
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_553
timestamp 0
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_559
timestamp 0
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_561
timestamp 0
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_573
timestamp 0
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_585
timestamp 0
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_597
timestamp 0
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_609
timestamp 0
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_615
timestamp 0
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_617
timestamp 0
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 0
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 0
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 0
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 0
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 0
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_53
timestamp 0
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_65
timestamp 0
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_77
timestamp 0
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 0
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_85
timestamp 0
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_97
timestamp 0
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_109
timestamp 0
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_121
timestamp 0
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_133
timestamp 0
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_139
timestamp 0
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 0
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 0
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_165
timestamp 0
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_177
timestamp 0
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_189
timestamp 0
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_195
timestamp 0
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_197
timestamp 0
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_209
timestamp 0
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_221
timestamp 0
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_233
timestamp 0
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_245
timestamp 0
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_251
timestamp 0
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_253
timestamp 0
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_265
timestamp 0
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_277
timestamp 0
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_289
timestamp 0
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_301
timestamp 0
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_307
timestamp 0
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_309
timestamp 0
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_321
timestamp 0
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_333
timestamp 0
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_345
timestamp 0
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_357
timestamp 0
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_363
timestamp 0
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_365
timestamp 0
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_377
timestamp 0
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_389
timestamp 0
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_401
timestamp 0
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_413
timestamp 0
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_419
timestamp 0
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_421
timestamp 0
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_433
timestamp 0
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_445
timestamp 0
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_457
timestamp 0
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_469
timestamp 0
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_475
timestamp 0
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_477
timestamp 0
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_489
timestamp 0
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_501
timestamp 0
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_513
timestamp 0
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_525
timestamp 0
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_531
timestamp 0
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_533
timestamp 0
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_545
timestamp 0
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_557
timestamp 0
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_569
timestamp 0
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_581
timestamp 0
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_587
timestamp 0
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_589
timestamp 0
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_601
timestamp 0
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82_613
timestamp 0
transform 1 0 57500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_621
timestamp 0
transform 1 0 58236 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_3
timestamp 0
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_15
timestamp 0
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_27
timestamp 0
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_39
timestamp 0
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_51
timestamp 0
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_55
timestamp 0
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_57
timestamp 0
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_69
timestamp 0
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_81
timestamp 0
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_93
timestamp 0
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_105
timestamp 0
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_111
timestamp 0
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_113
timestamp 0
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_125
timestamp 0
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_137
timestamp 0
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_149
timestamp 0
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_161
timestamp 0
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_167
timestamp 0
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_169
timestamp 0
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_181
timestamp 0
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_193
timestamp 0
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_205
timestamp 0
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_217
timestamp 0
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_223
timestamp 0
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_225
timestamp 0
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_237
timestamp 0
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_249
timestamp 0
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_261
timestamp 0
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_273
timestamp 0
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_279
timestamp 0
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_281
timestamp 0
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_293
timestamp 0
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_305
timestamp 0
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_317
timestamp 0
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_329
timestamp 0
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_335
timestamp 0
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_337
timestamp 0
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_349
timestamp 0
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_361
timestamp 0
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_373
timestamp 0
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_385
timestamp 0
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_391
timestamp 0
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_393
timestamp 0
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_405
timestamp 0
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_417
timestamp 0
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_429
timestamp 0
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_441
timestamp 0
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_447
timestamp 0
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_449
timestamp 0
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_461
timestamp 0
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_473
timestamp 0
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_485
timestamp 0
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_497
timestamp 0
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_503
timestamp 0
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_505
timestamp 0
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_517
timestamp 0
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_529
timestamp 0
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_541
timestamp 0
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_553
timestamp 0
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_559
timestamp 0
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_561
timestamp 0
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_573
timestamp 0
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_585
timestamp 0
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_597
timestamp 0
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_609
timestamp 0
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_615
timestamp 0
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_617
timestamp 0
transform 1 0 57868 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_621
timestamp 0
transform 1 0 58236 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_3
timestamp 0
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_15
timestamp 0
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 0
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_29
timestamp 0
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_41
timestamp 0
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_53
timestamp 0
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_65
timestamp 0
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 0
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 0
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_85
timestamp 0
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_97
timestamp 0
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_109
timestamp 0
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_121
timestamp 0
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_133
timestamp 0
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_139
timestamp 0
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_141
timestamp 0
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_153
timestamp 0
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_165
timestamp 0
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_177
timestamp 0
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_189
timestamp 0
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_195
timestamp 0
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_197
timestamp 0
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_209
timestamp 0
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_221
timestamp 0
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_233
timestamp 0
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_245
timestamp 0
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_251
timestamp 0
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_253
timestamp 0
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_265
timestamp 0
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_277
timestamp 0
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_289
timestamp 0
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_301
timestamp 0
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_307
timestamp 0
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_309
timestamp 0
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_321
timestamp 0
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_333
timestamp 0
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_345
timestamp 0
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_357
timestamp 0
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_363
timestamp 0
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_365
timestamp 0
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_377
timestamp 0
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_389
timestamp 0
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_401
timestamp 0
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_413
timestamp 0
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_419
timestamp 0
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_421
timestamp 0
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_433
timestamp 0
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_445
timestamp 0
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_457
timestamp 0
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_469
timestamp 0
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_475
timestamp 0
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_477
timestamp 0
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_489
timestamp 0
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_501
timestamp 0
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_513
timestamp 0
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_525
timestamp 0
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_531
timestamp 0
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_533
timestamp 0
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_545
timestamp 0
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_557
timestamp 0
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_569
timestamp 0
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_581
timestamp 0
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_587
timestamp 0
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_589
timestamp 0
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_601
timestamp 0
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_613
timestamp 0
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_3
timestamp 0
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_15
timestamp 0
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_27
timestamp 0
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_39
timestamp 0
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_51
timestamp 0
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_55
timestamp 0
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_57
timestamp 0
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 0
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 0
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_93
timestamp 0
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_105
timestamp 0
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_111
timestamp 0
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_113
timestamp 0
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_125
timestamp 0
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_137
timestamp 0
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_149
timestamp 0
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_161
timestamp 0
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_167
timestamp 0
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_169
timestamp 0
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_181
timestamp 0
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_193
timestamp 0
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_205
timestamp 0
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_217
timestamp 0
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_223
timestamp 0
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_225
timestamp 0
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_237
timestamp 0
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_249
timestamp 0
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_261
timestamp 0
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_273
timestamp 0
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_279
timestamp 0
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_281
timestamp 0
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_293
timestamp 0
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_305
timestamp 0
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_317
timestamp 0
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_329
timestamp 0
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_335
timestamp 0
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_337
timestamp 0
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_349
timestamp 0
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_361
timestamp 0
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_373
timestamp 0
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_385
timestamp 0
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_391
timestamp 0
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_393
timestamp 0
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_405
timestamp 0
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_417
timestamp 0
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_429
timestamp 0
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_441
timestamp 0
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_447
timestamp 0
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_449
timestamp 0
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_461
timestamp 0
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_473
timestamp 0
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_485
timestamp 0
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_497
timestamp 0
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_503
timestamp 0
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_505
timestamp 0
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_517
timestamp 0
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_529
timestamp 0
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_541
timestamp 0
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_553
timestamp 0
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_559
timestamp 0
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_561
timestamp 0
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_573
timestamp 0
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_585
timestamp 0
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_597
timestamp 0
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_609
timestamp 0
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_615
timestamp 0
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_617
timestamp 0
transform 1 0 57868 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_621
timestamp 0
transform 1 0 58236 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_3
timestamp 0
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_15
timestamp 0
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 0
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 0
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 0
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_53
timestamp 0
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_65
timestamp 0
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_77
timestamp 0
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_83
timestamp 0
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_85
timestamp 0
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_97
timestamp 0
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_109
timestamp 0
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_121
timestamp 0
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_133
timestamp 0
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_139
timestamp 0
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_141
timestamp 0
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_153
timestamp 0
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_165
timestamp 0
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_177
timestamp 0
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_189
timestamp 0
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_195
timestamp 0
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_197
timestamp 0
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_209
timestamp 0
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_221
timestamp 0
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_233
timestamp 0
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_245
timestamp 0
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_251
timestamp 0
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_253
timestamp 0
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_265
timestamp 0
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_277
timestamp 0
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_289
timestamp 0
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_301
timestamp 0
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_307
timestamp 0
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_309
timestamp 0
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_321
timestamp 0
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_333
timestamp 0
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_345
timestamp 0
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_357
timestamp 0
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_363
timestamp 0
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_365
timestamp 0
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_377
timestamp 0
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_389
timestamp 0
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_401
timestamp 0
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_413
timestamp 0
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_419
timestamp 0
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_421
timestamp 0
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_433
timestamp 0
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_445
timestamp 0
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_457
timestamp 0
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_469
timestamp 0
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_475
timestamp 0
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_477
timestamp 0
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_489
timestamp 0
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_501
timestamp 0
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_513
timestamp 0
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_525
timestamp 0
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_531
timestamp 0
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_533
timestamp 0
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_545
timestamp 0
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_557
timestamp 0
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_569
timestamp 0
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_581
timestamp 0
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_587
timestamp 0
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_589
timestamp 0
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_601
timestamp 0
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_613
timestamp 0
transform 1 0 57500 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_621
timestamp 0
transform 1 0 58236 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_3
timestamp 0
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_15
timestamp 0
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_27
timestamp 0
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_39
timestamp 0
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_51
timestamp 0
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_55
timestamp 0
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_57
timestamp 0
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_69
timestamp 0
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_81
timestamp 0
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_93
timestamp 0
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_105
timestamp 0
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_111
timestamp 0
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_113
timestamp 0
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_125
timestamp 0
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_137
timestamp 0
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_149
timestamp 0
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_161
timestamp 0
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_167
timestamp 0
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_169
timestamp 0
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_181
timestamp 0
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_193
timestamp 0
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_205
timestamp 0
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_217
timestamp 0
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_223
timestamp 0
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_225
timestamp 0
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_237
timestamp 0
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_249
timestamp 0
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_261
timestamp 0
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_273
timestamp 0
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_279
timestamp 0
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_281
timestamp 0
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_293
timestamp 0
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_305
timestamp 0
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_317
timestamp 0
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_329
timestamp 0
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_335
timestamp 0
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_337
timestamp 0
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_349
timestamp 0
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_361
timestamp 0
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_373
timestamp 0
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_385
timestamp 0
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_391
timestamp 0
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_393
timestamp 0
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_405
timestamp 0
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_417
timestamp 0
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_429
timestamp 0
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_441
timestamp 0
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_447
timestamp 0
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_449
timestamp 0
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_461
timestamp 0
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_473
timestamp 0
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_485
timestamp 0
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_497
timestamp 0
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_503
timestamp 0
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_505
timestamp 0
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_517
timestamp 0
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_529
timestamp 0
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_541
timestamp 0
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_553
timestamp 0
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_559
timestamp 0
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_561
timestamp 0
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_573
timestamp 0
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_585
timestamp 0
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_597
timestamp 0
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_609
timestamp 0
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_615
timestamp 0
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_617
timestamp 0
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_3
timestamp 0
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_15
timestamp 0
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 0
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 0
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 0
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_53
timestamp 0
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_65
timestamp 0
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_77
timestamp 0
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 0
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_85
timestamp 0
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_97
timestamp 0
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_109
timestamp 0
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_121
timestamp 0
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_133
timestamp 0
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_139
timestamp 0
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_141
timestamp 0
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_153
timestamp 0
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_165
timestamp 0
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_177
timestamp 0
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_189
timestamp 0
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_195
timestamp 0
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_197
timestamp 0
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_209
timestamp 0
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_221
timestamp 0
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_233
timestamp 0
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_245
timestamp 0
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_251
timestamp 0
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_253
timestamp 0
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_265
timestamp 0
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_277
timestamp 0
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_289
timestamp 0
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_301
timestamp 0
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_307
timestamp 0
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_309
timestamp 0
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_321
timestamp 0
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_333
timestamp 0
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_345
timestamp 0
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_357
timestamp 0
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_363
timestamp 0
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_365
timestamp 0
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_377
timestamp 0
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_389
timestamp 0
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_401
timestamp 0
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_413
timestamp 0
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_419
timestamp 0
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_421
timestamp 0
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_433
timestamp 0
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_445
timestamp 0
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_457
timestamp 0
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_469
timestamp 0
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_475
timestamp 0
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_477
timestamp 0
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_489
timestamp 0
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_501
timestamp 0
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_513
timestamp 0
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_525
timestamp 0
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_531
timestamp 0
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_533
timestamp 0
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_545
timestamp 0
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_557
timestamp 0
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_569
timestamp 0
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_581
timestamp 0
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_587
timestamp 0
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_589
timestamp 0
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_601
timestamp 0
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88_613
timestamp 0
transform 1 0 57500 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_621
timestamp 0
transform 1 0 58236 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_3
timestamp 0
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_15
timestamp 0
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_27
timestamp 0
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_39
timestamp 0
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_51
timestamp 0
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 0
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_57
timestamp 0
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_69
timestamp 0
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_81
timestamp 0
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_93
timestamp 0
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_105
timestamp 0
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_111
timestamp 0
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_113
timestamp 0
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_125
timestamp 0
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_137
timestamp 0
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_149
timestamp 0
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_161
timestamp 0
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_167
timestamp 0
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_169
timestamp 0
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_181
timestamp 0
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_193
timestamp 0
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_205
timestamp 0
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_217
timestamp 0
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_223
timestamp 0
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_225
timestamp 0
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_237
timestamp 0
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_249
timestamp 0
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_261
timestamp 0
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_273
timestamp 0
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_279
timestamp 0
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_281
timestamp 0
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_293
timestamp 0
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_305
timestamp 0
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_317
timestamp 0
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_329
timestamp 0
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_335
timestamp 0
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_337
timestamp 0
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_349
timestamp 0
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_361
timestamp 0
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_373
timestamp 0
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_385
timestamp 0
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_391
timestamp 0
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_393
timestamp 0
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_405
timestamp 0
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_417
timestamp 0
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_429
timestamp 0
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_441
timestamp 0
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_447
timestamp 0
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_449
timestamp 0
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_461
timestamp 0
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_473
timestamp 0
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_485
timestamp 0
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_497
timestamp 0
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_503
timestamp 0
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_505
timestamp 0
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_517
timestamp 0
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_529
timestamp 0
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_541
timestamp 0
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_553
timestamp 0
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_559
timestamp 0
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_561
timestamp 0
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_573
timestamp 0
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_585
timestamp 0
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_597
timestamp 0
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_609
timestamp 0
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_615
timestamp 0
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_617
timestamp 0
transform 1 0 57868 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_621
timestamp 0
transform 1 0 58236 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_3
timestamp 0
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_15
timestamp 0
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 0
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 0
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 0
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 0
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 0
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 0
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 0
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_85
timestamp 0
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_97
timestamp 0
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_109
timestamp 0
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_121
timestamp 0
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_133
timestamp 0
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_139
timestamp 0
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_141
timestamp 0
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_153
timestamp 0
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_165
timestamp 0
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_177
timestamp 0
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_189
timestamp 0
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_195
timestamp 0
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_197
timestamp 0
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_209
timestamp 0
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_221
timestamp 0
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_233
timestamp 0
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_245
timestamp 0
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_251
timestamp 0
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_253
timestamp 0
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_265
timestamp 0
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_277
timestamp 0
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_289
timestamp 0
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_301
timestamp 0
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_307
timestamp 0
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_309
timestamp 0
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_321
timestamp 0
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_333
timestamp 0
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_345
timestamp 0
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_357
timestamp 0
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_363
timestamp 0
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_365
timestamp 0
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_377
timestamp 0
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_389
timestamp 0
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_401
timestamp 0
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_413
timestamp 0
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_419
timestamp 0
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_421
timestamp 0
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_433
timestamp 0
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_445
timestamp 0
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_457
timestamp 0
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_469
timestamp 0
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_475
timestamp 0
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_477
timestamp 0
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_489
timestamp 0
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_501
timestamp 0
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_513
timestamp 0
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_525
timestamp 0
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_531
timestamp 0
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_533
timestamp 0
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_545
timestamp 0
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_557
timestamp 0
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_569
timestamp 0
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_581
timestamp 0
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_587
timestamp 0
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_589
timestamp 0
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_601
timestamp 0
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_613
timestamp 0
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 0
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 0
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_27
timestamp 0
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_39
timestamp 0
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_51
timestamp 0
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_55
timestamp 0
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_57
timestamp 0
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_69
timestamp 0
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_81
timestamp 0
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_93
timestamp 0
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_105
timestamp 0
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_111
timestamp 0
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_113
timestamp 0
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_125
timestamp 0
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_137
timestamp 0
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_149
timestamp 0
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_161
timestamp 0
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_167
timestamp 0
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_169
timestamp 0
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_181
timestamp 0
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_193
timestamp 0
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_205
timestamp 0
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_217
timestamp 0
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_223
timestamp 0
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_225
timestamp 0
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_237
timestamp 0
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_249
timestamp 0
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_261
timestamp 0
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_273
timestamp 0
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_279
timestamp 0
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_281
timestamp 0
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_293
timestamp 0
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_305
timestamp 0
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_317
timestamp 0
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_329
timestamp 0
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_335
timestamp 0
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_337
timestamp 0
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_349
timestamp 0
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_361
timestamp 0
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_373
timestamp 0
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_385
timestamp 0
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_391
timestamp 0
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_393
timestamp 0
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_405
timestamp 0
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_417
timestamp 0
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_429
timestamp 0
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_441
timestamp 0
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_447
timestamp 0
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_449
timestamp 0
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_461
timestamp 0
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_473
timestamp 0
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_485
timestamp 0
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_497
timestamp 0
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_503
timestamp 0
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_505
timestamp 0
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_517
timestamp 0
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_529
timestamp 0
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_541
timestamp 0
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_553
timestamp 0
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_559
timestamp 0
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_561
timestamp 0
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_573
timestamp 0
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_585
timestamp 0
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_597
timestamp 0
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_609
timestamp 0
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_615
timestamp 0
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_617
timestamp 0
transform 1 0 57868 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_621
timestamp 0
transform 1 0 58236 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_3
timestamp 0
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_15
timestamp 0
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 0
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_29
timestamp 0
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_41
timestamp 0
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_53
timestamp 0
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_65
timestamp 0
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_77
timestamp 0
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_83
timestamp 0
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_85
timestamp 0
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_97
timestamp 0
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_109
timestamp 0
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_121
timestamp 0
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_133
timestamp 0
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_139
timestamp 0
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_141
timestamp 0
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_153
timestamp 0
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_165
timestamp 0
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_177
timestamp 0
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_189
timestamp 0
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_195
timestamp 0
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_197
timestamp 0
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_209
timestamp 0
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_221
timestamp 0
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_233
timestamp 0
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_245
timestamp 0
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_251
timestamp 0
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_253
timestamp 0
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_265
timestamp 0
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_277
timestamp 0
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_289
timestamp 0
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_301
timestamp 0
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_307
timestamp 0
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_309
timestamp 0
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_321
timestamp 0
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_333
timestamp 0
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_345
timestamp 0
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_357
timestamp 0
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_363
timestamp 0
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_365
timestamp 0
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_377
timestamp 0
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_389
timestamp 0
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_401
timestamp 0
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_413
timestamp 0
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_419
timestamp 0
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_421
timestamp 0
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_433
timestamp 0
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_445
timestamp 0
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_457
timestamp 0
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_469
timestamp 0
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_475
timestamp 0
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_477
timestamp 0
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_489
timestamp 0
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_501
timestamp 0
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_513
timestamp 0
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_525
timestamp 0
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_531
timestamp 0
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_533
timestamp 0
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_545
timestamp 0
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_557
timestamp 0
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_569
timestamp 0
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_581
timestamp 0
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_587
timestamp 0
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_589
timestamp 0
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_601
timestamp 0
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_613
timestamp 0
transform 1 0 57500 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_621
timestamp 0
transform 1 0 58236 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 0
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 0
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_27
timestamp 0
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_39
timestamp 0
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_51
timestamp 0
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_55
timestamp 0
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_57
timestamp 0
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_69
timestamp 0
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_81
timestamp 0
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_93
timestamp 0
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_105
timestamp 0
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_111
timestamp 0
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_113
timestamp 0
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_125
timestamp 0
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_137
timestamp 0
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_149
timestamp 0
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_161
timestamp 0
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_167
timestamp 0
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_169
timestamp 0
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_181
timestamp 0
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_193
timestamp 0
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_205
timestamp 0
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_217
timestamp 0
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_223
timestamp 0
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_225
timestamp 0
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_237
timestamp 0
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_249
timestamp 0
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_261
timestamp 0
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_273
timestamp 0
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_279
timestamp 0
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_281
timestamp 0
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_293
timestamp 0
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_305
timestamp 0
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_317
timestamp 0
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_329
timestamp 0
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_335
timestamp 0
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_337
timestamp 0
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_349
timestamp 0
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_361
timestamp 0
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_373
timestamp 0
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_385
timestamp 0
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_391
timestamp 0
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_393
timestamp 0
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_405
timestamp 0
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_417
timestamp 0
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_429
timestamp 0
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_441
timestamp 0
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_447
timestamp 0
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_449
timestamp 0
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_461
timestamp 0
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_473
timestamp 0
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_485
timestamp 0
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_497
timestamp 0
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_503
timestamp 0
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_505
timestamp 0
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_517
timestamp 0
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_529
timestamp 0
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_541
timestamp 0
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_553
timestamp 0
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_559
timestamp 0
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_561
timestamp 0
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_573
timestamp 0
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_585
timestamp 0
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_597
timestamp 0
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_609
timestamp 0
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_615
timestamp 0
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_617
timestamp 0
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_3
timestamp 0
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_15
timestamp 0
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 0
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_29
timestamp 0
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_41
timestamp 0
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_53
timestamp 0
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_65
timestamp 0
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_77
timestamp 0
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_83
timestamp 0
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_85
timestamp 0
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_97
timestamp 0
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_109
timestamp 0
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_121
timestamp 0
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_133
timestamp 0
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_139
timestamp 0
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_141
timestamp 0
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_153
timestamp 0
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_165
timestamp 0
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_177
timestamp 0
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_189
timestamp 0
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_195
timestamp 0
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_197
timestamp 0
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_209
timestamp 0
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_221
timestamp 0
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_233
timestamp 0
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_245
timestamp 0
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_251
timestamp 0
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_253
timestamp 0
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_265
timestamp 0
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_277
timestamp 0
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_289
timestamp 0
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_301
timestamp 0
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_307
timestamp 0
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_309
timestamp 0
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_321
timestamp 0
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_333
timestamp 0
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_345
timestamp 0
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_357
timestamp 0
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_363
timestamp 0
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_365
timestamp 0
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_377
timestamp 0
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_389
timestamp 0
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_401
timestamp 0
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_413
timestamp 0
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_419
timestamp 0
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_421
timestamp 0
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_433
timestamp 0
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_445
timestamp 0
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_457
timestamp 0
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_469
timestamp 0
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_475
timestamp 0
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_477
timestamp 0
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_489
timestamp 0
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_501
timestamp 0
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_513
timestamp 0
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_525
timestamp 0
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_531
timestamp 0
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_533
timestamp 0
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_545
timestamp 0
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_557
timestamp 0
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_569
timestamp 0
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_581
timestamp 0
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_587
timestamp 0
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_589
timestamp 0
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_601
timestamp 0
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94_613
timestamp 0
transform 1 0 57500 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_621
timestamp 0
transform 1 0 58236 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_3
timestamp 0
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_15
timestamp 0
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_27
timestamp 0
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_39
timestamp 0
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_51
timestamp 0
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_55
timestamp 0
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_57
timestamp 0
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_69
timestamp 0
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_81
timestamp 0
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_93
timestamp 0
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_105
timestamp 0
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_111
timestamp 0
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_113
timestamp 0
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_125
timestamp 0
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_137
timestamp 0
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_149
timestamp 0
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_161
timestamp 0
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_167
timestamp 0
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_169
timestamp 0
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_181
timestamp 0
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_193
timestamp 0
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_205
timestamp 0
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_217
timestamp 0
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_223
timestamp 0
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_225
timestamp 0
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_237
timestamp 0
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_249
timestamp 0
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_261
timestamp 0
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_273
timestamp 0
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_279
timestamp 0
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_281
timestamp 0
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_293
timestamp 0
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_305
timestamp 0
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_317
timestamp 0
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_329
timestamp 0
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_335
timestamp 0
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_337
timestamp 0
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_349
timestamp 0
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_361
timestamp 0
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_373
timestamp 0
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_385
timestamp 0
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_391
timestamp 0
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_393
timestamp 0
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_405
timestamp 0
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_417
timestamp 0
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_429
timestamp 0
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_441
timestamp 0
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_447
timestamp 0
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_449
timestamp 0
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_461
timestamp 0
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_473
timestamp 0
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_485
timestamp 0
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_497
timestamp 0
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_503
timestamp 0
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_505
timestamp 0
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_517
timestamp 0
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_529
timestamp 0
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_541
timestamp 0
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_553
timestamp 0
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_559
timestamp 0
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_561
timestamp 0
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_573
timestamp 0
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_585
timestamp 0
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_597
timestamp 0
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_609
timestamp 0
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_615
timestamp 0
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_617
timestamp 0
transform 1 0 57868 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_621
timestamp 0
transform 1 0 58236 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 0
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 0
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 0
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_29
timestamp 0
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_41
timestamp 0
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_53
timestamp 0
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_65
timestamp 0
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_77
timestamp 0
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 0
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_85
timestamp 0
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_97
timestamp 0
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_109
timestamp 0
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_121
timestamp 0
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_133
timestamp 0
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_139
timestamp 0
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_141
timestamp 0
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_153
timestamp 0
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_165
timestamp 0
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_177
timestamp 0
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_189
timestamp 0
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_195
timestamp 0
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_197
timestamp 0
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_209
timestamp 0
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_221
timestamp 0
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_233
timestamp 0
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_245
timestamp 0
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_251
timestamp 0
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_253
timestamp 0
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_265
timestamp 0
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_277
timestamp 0
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_289
timestamp 0
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_301
timestamp 0
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_307
timestamp 0
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_309
timestamp 0
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_321
timestamp 0
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_333
timestamp 0
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_345
timestamp 0
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_357
timestamp 0
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_363
timestamp 0
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_365
timestamp 0
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_377
timestamp 0
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_389
timestamp 0
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_401
timestamp 0
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_413
timestamp 0
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_419
timestamp 0
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_421
timestamp 0
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_433
timestamp 0
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_445
timestamp 0
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_457
timestamp 0
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_469
timestamp 0
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_475
timestamp 0
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_477
timestamp 0
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_489
timestamp 0
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_501
timestamp 0
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_513
timestamp 0
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_525
timestamp 0
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_531
timestamp 0
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_533
timestamp 0
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_545
timestamp 0
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_557
timestamp 0
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_569
timestamp 0
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_581
timestamp 0
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_587
timestamp 0
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_589
timestamp 0
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_601
timestamp 0
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_613
timestamp 0
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_3
timestamp 0
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_15
timestamp 0
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_27
timestamp 0
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_39
timestamp 0
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_51
timestamp 0
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_55
timestamp 0
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_57
timestamp 0
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_69
timestamp 0
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_81
timestamp 0
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_93
timestamp 0
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_105
timestamp 0
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_111
timestamp 0
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_113
timestamp 0
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_125
timestamp 0
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_137
timestamp 0
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_149
timestamp 0
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_161
timestamp 0
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_167
timestamp 0
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_169
timestamp 0
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_181
timestamp 0
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_193
timestamp 0
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_205
timestamp 0
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_217
timestamp 0
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_223
timestamp 0
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_225
timestamp 0
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_237
timestamp 0
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_249
timestamp 0
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_261
timestamp 0
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_273
timestamp 0
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_279
timestamp 0
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_281
timestamp 0
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_293
timestamp 0
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_305
timestamp 0
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_317
timestamp 0
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_329
timestamp 0
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_335
timestamp 0
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_337
timestamp 0
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_349
timestamp 0
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_361
timestamp 0
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_373
timestamp 0
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_385
timestamp 0
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_391
timestamp 0
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_393
timestamp 0
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_405
timestamp 0
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_417
timestamp 0
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_429
timestamp 0
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_441
timestamp 0
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_447
timestamp 0
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_449
timestamp 0
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_461
timestamp 0
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_473
timestamp 0
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_485
timestamp 0
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_497
timestamp 0
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_503
timestamp 0
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_505
timestamp 0
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_517
timestamp 0
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_529
timestamp 0
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_541
timestamp 0
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_553
timestamp 0
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_559
timestamp 0
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_561
timestamp 0
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_573
timestamp 0
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_585
timestamp 0
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_597
timestamp 0
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_609
timestamp 0
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_615
timestamp 0
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_617
timestamp 0
transform 1 0 57868 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_621
timestamp 0
transform 1 0 58236 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_3
timestamp 0
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_15
timestamp 0
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 0
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_29
timestamp 0
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_41
timestamp 0
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_53
timestamp 0
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_65
timestamp 0
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_77
timestamp 0
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_83
timestamp 0
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_85
timestamp 0
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_97
timestamp 0
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_109
timestamp 0
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_121
timestamp 0
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_133
timestamp 0
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_139
timestamp 0
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_141
timestamp 0
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_153
timestamp 0
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_165
timestamp 0
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_177
timestamp 0
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_189
timestamp 0
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_195
timestamp 0
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_197
timestamp 0
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_209
timestamp 0
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_221
timestamp 0
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_233
timestamp 0
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_245
timestamp 0
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_251
timestamp 0
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_253
timestamp 0
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_265
timestamp 0
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_277
timestamp 0
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_289
timestamp 0
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_301
timestamp 0
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_307
timestamp 0
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_309
timestamp 0
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_321
timestamp 0
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_333
timestamp 0
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_345
timestamp 0
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_357
timestamp 0
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_363
timestamp 0
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_365
timestamp 0
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_377
timestamp 0
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_389
timestamp 0
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_401
timestamp 0
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_413
timestamp 0
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_419
timestamp 0
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_421
timestamp 0
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_433
timestamp 0
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_445
timestamp 0
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_457
timestamp 0
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_469
timestamp 0
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_475
timestamp 0
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_477
timestamp 0
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_489
timestamp 0
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_501
timestamp 0
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_513
timestamp 0
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_525
timestamp 0
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_531
timestamp 0
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_533
timestamp 0
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_545
timestamp 0
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_557
timestamp 0
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_569
timestamp 0
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_581
timestamp 0
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_587
timestamp 0
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_589
timestamp 0
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_601
timestamp 0
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_613
timestamp 0
transform 1 0 57500 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_621
timestamp 0
transform 1 0 58236 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_3
timestamp 0
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_15
timestamp 0
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_27
timestamp 0
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_39
timestamp 0
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_51
timestamp 0
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_55
timestamp 0
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 0
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 0
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 0
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_93
timestamp 0
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_105
timestamp 0
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_111
timestamp 0
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_113
timestamp 0
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_125
timestamp 0
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_137
timestamp 0
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_149
timestamp 0
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_161
timestamp 0
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_167
timestamp 0
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_169
timestamp 0
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_181
timestamp 0
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_193
timestamp 0
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_205
timestamp 0
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_217
timestamp 0
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_223
timestamp 0
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_225
timestamp 0
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_237
timestamp 0
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_249
timestamp 0
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_261
timestamp 0
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_273
timestamp 0
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_279
timestamp 0
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_281
timestamp 0
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_293
timestamp 0
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_305
timestamp 0
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_317
timestamp 0
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_329
timestamp 0
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_335
timestamp 0
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_337
timestamp 0
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_349
timestamp 0
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_361
timestamp 0
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_373
timestamp 0
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_385
timestamp 0
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_391
timestamp 0
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_393
timestamp 0
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_405
timestamp 0
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_417
timestamp 0
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_429
timestamp 0
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_441
timestamp 0
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_447
timestamp 0
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_449
timestamp 0
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_461
timestamp 0
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_473
timestamp 0
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_485
timestamp 0
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_497
timestamp 0
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_503
timestamp 0
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_505
timestamp 0
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_517
timestamp 0
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_529
timestamp 0
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_541
timestamp 0
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_553
timestamp 0
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_559
timestamp 0
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_561
timestamp 0
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_573
timestamp 0
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_585
timestamp 0
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_597
timestamp 0
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_609
timestamp 0
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_615
timestamp 0
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_617
timestamp 0
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_3
timestamp 0
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_15
timestamp 0
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 0
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_29
timestamp 0
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_41
timestamp 0
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_53
timestamp 0
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_65
timestamp 0
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_77
timestamp 0
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_83
timestamp 0
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_85
timestamp 0
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_97
timestamp 0
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_109
timestamp 0
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_121
timestamp 0
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_133
timestamp 0
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_139
timestamp 0
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_141
timestamp 0
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_153
timestamp 0
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_165
timestamp 0
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_177
timestamp 0
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_189
timestamp 0
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_195
timestamp 0
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_197
timestamp 0
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_209
timestamp 0
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_221
timestamp 0
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_233
timestamp 0
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_245
timestamp 0
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_251
timestamp 0
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_253
timestamp 0
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_265
timestamp 0
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_277
timestamp 0
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_289
timestamp 0
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_301
timestamp 0
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_307
timestamp 0
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_309
timestamp 0
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_321
timestamp 0
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_333
timestamp 0
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_345
timestamp 0
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_357
timestamp 0
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_363
timestamp 0
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_365
timestamp 0
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_377
timestamp 0
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_389
timestamp 0
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_401
timestamp 0
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_413
timestamp 0
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_419
timestamp 0
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_421
timestamp 0
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_433
timestamp 0
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_445
timestamp 0
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_457
timestamp 0
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_469
timestamp 0
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_475
timestamp 0
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_477
timestamp 0
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_489
timestamp 0
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_501
timestamp 0
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_513
timestamp 0
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_525
timestamp 0
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_531
timestamp 0
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_533
timestamp 0
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_545
timestamp 0
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_557
timestamp 0
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_569
timestamp 0
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_581
timestamp 0
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_587
timestamp 0
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_589
timestamp 0
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_601
timestamp 0
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_613
timestamp 0
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_3
timestamp 0
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_15
timestamp 0
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_27
timestamp 0
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_29
timestamp 0
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_41
timestamp 0
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_53
timestamp 0
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_57
timestamp 0
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_69
timestamp 0
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_81
timestamp 0
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_85
timestamp 0
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_97
timestamp 0
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_109
timestamp 0
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_113
timestamp 0
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_125
timestamp 0
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_137
timestamp 0
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_141
timestamp 0
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_153
timestamp 0
transform 1 0 15180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_165
timestamp 0
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_169
timestamp 0
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_181
timestamp 0
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_193
timestamp 0
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_197
timestamp 0
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_209
timestamp 0
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_221
timestamp 0
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_225
timestamp 0
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_237
timestamp 0
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_249
timestamp 0
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_253
timestamp 0
transform 1 0 24380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_265
timestamp 0
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_277
timestamp 0
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_281
timestamp 0
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_293
timestamp 0
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_305
timestamp 0
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_309
timestamp 0
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_321
timestamp 0
transform 1 0 30636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_333
timestamp 0
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_337
timestamp 0
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_349
timestamp 0
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_361
timestamp 0
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_365
timestamp 0
transform 1 0 34684 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_377
timestamp 0
transform 1 0 35788 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_389
timestamp 0
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_393
timestamp 0
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_405
timestamp 0
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_417
timestamp 0
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_421
timestamp 0
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_433
timestamp 0
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_445
timestamp 0
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_449
timestamp 0
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_461
timestamp 0
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_473
timestamp 0
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_477
timestamp 0
transform 1 0 44988 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_489
timestamp 0
transform 1 0 46092 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_501
timestamp 0
transform 1 0 47196 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_505
timestamp 0
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_517
timestamp 0
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_529
timestamp 0
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_533
timestamp 0
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_545
timestamp 0
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_557
timestamp 0
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_561
timestamp 0
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_573
timestamp 0
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_585
timestamp 0
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_589
timestamp 0
transform 1 0 55292 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_601
timestamp 0
transform 1 0 56396 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_613
timestamp 0
transform 1 0 57500 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_617
timestamp 0
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_102
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_103
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_104
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_105
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_106
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_107
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_108
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_109
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_110
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_111
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_112
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_113
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_114
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_115
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_116
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_117
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_118
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_119
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_120
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_121
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_122
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_123
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_124
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_125
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_126
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_127
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_128
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_129
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_130
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_131
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_132
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_133
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 0
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_134
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 0
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_135
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 0
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_136
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 0
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_137
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 0
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_138
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 0
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_139
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 0
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_140
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 0
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_141
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 0
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_142
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 0
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_143
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 0
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_144
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 0
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_145
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 0
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_146
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 0
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_147
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 0
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_148
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 0
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_149
timestamp 0
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 0
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_150
timestamp 0
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 0
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_151
timestamp 0
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 0
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_152
timestamp 0
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 0
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_153
timestamp 0
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 0
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_154
timestamp 0
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 0
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_155
timestamp 0
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 0
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_156
timestamp 0
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 0
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_157
timestamp 0
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 0
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_158
timestamp 0
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 0
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_159
timestamp 0
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 0
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_160
timestamp 0
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 0
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_161
timestamp 0
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 0
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_162
timestamp 0
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 0
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_163
timestamp 0
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 0
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_164
timestamp 0
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 0
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_165
timestamp 0
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 0
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_166
timestamp 0
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 0
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_167
timestamp 0
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 0
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_168
timestamp 0
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 0
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_169
timestamp 0
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 0
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_170
timestamp 0
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 0
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_171
timestamp 0
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 0
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_172
timestamp 0
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 0
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_173
timestamp 0
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 0
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_174
timestamp 0
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 0
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_175
timestamp 0
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 0
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_176
timestamp 0
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 0
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_177
timestamp 0
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 0
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_178
timestamp 0
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 0
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_179
timestamp 0
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 0
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_180
timestamp 0
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 0
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_181
timestamp 0
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 0
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_182
timestamp 0
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 0
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_183
timestamp 0
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 0
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_184
timestamp 0
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 0
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Left_185
timestamp 0
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Right_83
timestamp 0
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Left_186
timestamp 0
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Right_84
timestamp 0
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Left_187
timestamp 0
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Right_85
timestamp 0
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Left_188
timestamp 0
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Right_86
timestamp 0
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Left_189
timestamp 0
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Right_87
timestamp 0
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Left_190
timestamp 0
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Right_88
timestamp 0
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Left_191
timestamp 0
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Right_89
timestamp 0
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Left_192
timestamp 0
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Right_90
timestamp 0
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Left_193
timestamp 0
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Right_91
timestamp 0
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Left_194
timestamp 0
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Right_92
timestamp 0
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Left_195
timestamp 0
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Right_93
timestamp 0
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Left_196
timestamp 0
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Right_94
timestamp 0
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Left_197
timestamp 0
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Right_95
timestamp 0
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Left_198
timestamp 0
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Right_96
timestamp 0
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Left_199
timestamp 0
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Right_97
timestamp 0
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Left_200
timestamp 0
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Right_98
timestamp 0
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Left_201
timestamp 0
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Right_99
timestamp 0
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Left_202
timestamp 0
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Right_100
timestamp 0
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Left_203
timestamp 0
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Right_101
timestamp 0
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_204
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_205
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_206
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_207
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_208
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_209
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_210
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_211
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_212
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_213
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_214
timestamp 0
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_215
timestamp 0
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_216
timestamp 0
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_217
timestamp 0
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_218
timestamp 0
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_219
timestamp 0
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_220
timestamp 0
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_221
timestamp 0
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_222
timestamp 0
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_223
timestamp 0
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_224
timestamp 0
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_225
timestamp 0
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_226
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_227
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_228
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_229
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_230
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_231
timestamp 0
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_232
timestamp 0
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_233
timestamp 0
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_234
timestamp 0
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_235
timestamp 0
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_236
timestamp 0
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_237
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_238
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_239
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_240
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_241
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_242
timestamp 0
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_243
timestamp 0
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_244
timestamp 0
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_245
timestamp 0
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_246
timestamp 0
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_247
timestamp 0
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_248
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_249
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_250
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_251
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_252
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_253
timestamp 0
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_254
timestamp 0
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_255
timestamp 0
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_256
timestamp 0
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_257
timestamp 0
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_258
timestamp 0
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_259
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_260
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_261
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_262
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_263
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_264
timestamp 0
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_265
timestamp 0
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_266
timestamp 0
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_267
timestamp 0
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_268
timestamp 0
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_269
timestamp 0
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_270
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_271
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_272
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_273
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_274
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_275
timestamp 0
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_276
timestamp 0
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_277
timestamp 0
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_278
timestamp 0
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_279
timestamp 0
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_280
timestamp 0
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_281
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_282
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_283
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_284
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_285
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_286
timestamp 0
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_287
timestamp 0
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_288
timestamp 0
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_289
timestamp 0
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_290
timestamp 0
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_291
timestamp 0
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_292
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_293
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_294
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_295
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_296
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_297
timestamp 0
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_298
timestamp 0
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_299
timestamp 0
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_300
timestamp 0
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_301
timestamp 0
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_302
timestamp 0
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_303
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_304
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_305
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_306
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_307
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_308
timestamp 0
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_309
timestamp 0
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_310
timestamp 0
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_311
timestamp 0
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_312
timestamp 0
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_313
timestamp 0
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_314
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_315
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_316
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_317
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_318
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_319
timestamp 0
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_320
timestamp 0
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_321
timestamp 0
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_322
timestamp 0
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_323
timestamp 0
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_324
timestamp 0
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_325
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_326
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_327
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_328
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_329
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_330
timestamp 0
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_331
timestamp 0
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_332
timestamp 0
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_333
timestamp 0
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_334
timestamp 0
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_335
timestamp 0
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_336
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_337
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_338
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_339
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_340
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_341
timestamp 0
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_342
timestamp 0
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_343
timestamp 0
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_344
timestamp 0
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_345
timestamp 0
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_346
timestamp 0
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_347
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_348
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_349
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_350
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_351
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_352
timestamp 0
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_353
timestamp 0
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_354
timestamp 0
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_355
timestamp 0
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_356
timestamp 0
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_357
timestamp 0
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_358
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_359
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_360
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_361
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_362
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_363
timestamp 0
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_364
timestamp 0
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_365
timestamp 0
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_366
timestamp 0
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_367
timestamp 0
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_368
timestamp 0
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_369
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_370
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_371
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_372
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_373
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_374
timestamp 0
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_375
timestamp 0
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_376
timestamp 0
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_377
timestamp 0
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_378
timestamp 0
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_379
timestamp 0
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_380
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_381
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_382
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_383
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_384
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_385
timestamp 0
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_386
timestamp 0
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_387
timestamp 0
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_388
timestamp 0
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_389
timestamp 0
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_390
timestamp 0
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_391
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_392
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_393
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_394
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_395
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_396
timestamp 0
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_397
timestamp 0
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_398
timestamp 0
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_399
timestamp 0
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_400
timestamp 0
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_401
timestamp 0
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_402
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_403
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_404
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_405
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_406
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_407
timestamp 0
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_408
timestamp 0
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_409
timestamp 0
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_410
timestamp 0
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_411
timestamp 0
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_412
timestamp 0
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_413
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_414
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_415
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_416
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_417
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_418
timestamp 0
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_419
timestamp 0
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_420
timestamp 0
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_421
timestamp 0
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_422
timestamp 0
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_423
timestamp 0
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_424
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_425
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_426
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_427
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_428
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_429
timestamp 0
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_430
timestamp 0
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_431
timestamp 0
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_432
timestamp 0
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_433
timestamp 0
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_434
timestamp 0
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_435
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_436
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_437
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_438
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_439
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_440
timestamp 0
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_441
timestamp 0
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_442
timestamp 0
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_443
timestamp 0
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_444
timestamp 0
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_445
timestamp 0
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_446
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_447
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_448
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_449
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_450
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_451
timestamp 0
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_452
timestamp 0
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_453
timestamp 0
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_454
timestamp 0
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_455
timestamp 0
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_456
timestamp 0
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_457
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_458
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_459
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_460
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_461
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_462
timestamp 0
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_463
timestamp 0
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_464
timestamp 0
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_465
timestamp 0
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_466
timestamp 0
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_467
timestamp 0
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_468
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_469
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_470
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_471
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_472
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_473
timestamp 0
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_474
timestamp 0
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_475
timestamp 0
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_476
timestamp 0
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_477
timestamp 0
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_478
timestamp 0
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_479
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_480
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_481
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_482
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_483
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_484
timestamp 0
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_485
timestamp 0
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_486
timestamp 0
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_487
timestamp 0
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_488
timestamp 0
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_489
timestamp 0
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_490
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_491
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_492
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_493
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_494
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_495
timestamp 0
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_496
timestamp 0
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_497
timestamp 0
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_498
timestamp 0
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_499
timestamp 0
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_500
timestamp 0
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_501
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_502
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_503
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_504
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_505
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_506
timestamp 0
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_507
timestamp 0
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_508
timestamp 0
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_509
timestamp 0
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_510
timestamp 0
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_511
timestamp 0
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_512
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_513
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_514
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_515
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_516
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_517
timestamp 0
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_518
timestamp 0
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_519
timestamp 0
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_520
timestamp 0
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_521
timestamp 0
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_522
timestamp 0
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_523
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_524
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_525
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_526
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_527
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_528
timestamp 0
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_529
timestamp 0
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_530
timestamp 0
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_531
timestamp 0
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_532
timestamp 0
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_533
timestamp 0
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_534
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_535
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_536
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_537
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_538
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_539
timestamp 0
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_540
timestamp 0
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_541
timestamp 0
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_542
timestamp 0
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_543
timestamp 0
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_544
timestamp 0
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_545
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_546
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_547
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_548
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_549
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_550
timestamp 0
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_551
timestamp 0
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_552
timestamp 0
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_553
timestamp 0
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_554
timestamp 0
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_555
timestamp 0
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_556
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_557
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_558
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_559
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_560
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_561
timestamp 0
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_562
timestamp 0
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_563
timestamp 0
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_564
timestamp 0
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_565
timestamp 0
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_566
timestamp 0
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_567
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_568
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_569
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_570
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_571
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_572
timestamp 0
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_573
timestamp 0
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_574
timestamp 0
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_575
timestamp 0
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_576
timestamp 0
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_577
timestamp 0
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_578
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_579
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_580
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_581
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_582
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_583
timestamp 0
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_584
timestamp 0
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_585
timestamp 0
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_586
timestamp 0
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_587
timestamp 0
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_588
timestamp 0
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_589
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_590
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_591
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_592
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_593
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_594
timestamp 0
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_595
timestamp 0
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_596
timestamp 0
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_597
timestamp 0
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_598
timestamp 0
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_599
timestamp 0
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_600
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_601
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_602
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_603
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_604
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_605
timestamp 0
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_606
timestamp 0
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_607
timestamp 0
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_608
timestamp 0
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_609
timestamp 0
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_610
timestamp 0
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_611
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_612
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_613
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_614
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_615
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_616
timestamp 0
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_617
timestamp 0
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_618
timestamp 0
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_619
timestamp 0
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_620
timestamp 0
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_621
timestamp 0
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_622
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_623
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_624
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_625
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_626
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_627
timestamp 0
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_628
timestamp 0
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_629
timestamp 0
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_630
timestamp 0
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_631
timestamp 0
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_632
timestamp 0
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_633
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_634
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_635
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_636
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_637
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_638
timestamp 0
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_639
timestamp 0
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_640
timestamp 0
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_641
timestamp 0
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_642
timestamp 0
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_643
timestamp 0
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_644
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_645
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_646
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_647
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_648
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_649
timestamp 0
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_650
timestamp 0
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_651
timestamp 0
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_652
timestamp 0
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_653
timestamp 0
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_654
timestamp 0
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_655
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_656
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_657
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_658
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_659
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_660
timestamp 0
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_661
timestamp 0
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_662
timestamp 0
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_663
timestamp 0
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_664
timestamp 0
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_665
timestamp 0
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_666
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_667
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_668
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_669
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_670
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_671
timestamp 0
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_672
timestamp 0
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_673
timestamp 0
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_674
timestamp 0
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_675
timestamp 0
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_676
timestamp 0
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_677
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_678
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_679
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_680
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_681
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_682
timestamp 0
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_683
timestamp 0
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_684
timestamp 0
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_685
timestamp 0
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_686
timestamp 0
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_687
timestamp 0
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_688
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_689
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_690
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_691
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_692
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_693
timestamp 0
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_694
timestamp 0
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_695
timestamp 0
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_696
timestamp 0
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_697
timestamp 0
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_698
timestamp 0
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_699
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_700
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_701
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_702
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_703
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_704
timestamp 0
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_705
timestamp 0
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_706
timestamp 0
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_707
timestamp 0
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_708
timestamp 0
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_709
timestamp 0
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_710
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_711
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_712
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_713
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_714
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_715
timestamp 0
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_716
timestamp 0
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_717
timestamp 0
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_718
timestamp 0
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_719
timestamp 0
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_720
timestamp 0
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_721
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_722
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_723
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_724
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_725
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_726
timestamp 0
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_727
timestamp 0
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_728
timestamp 0
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_729
timestamp 0
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_730
timestamp 0
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_731
timestamp 0
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_732
timestamp 0
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_733
timestamp 0
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_734
timestamp 0
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_735
timestamp 0
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_736
timestamp 0
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_737
timestamp 0
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_738
timestamp 0
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_739
timestamp 0
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_740
timestamp 0
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_741
timestamp 0
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_742
timestamp 0
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_743
timestamp 0
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_744
timestamp 0
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_745
timestamp 0
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_746
timestamp 0
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_747
timestamp 0
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_748
timestamp 0
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_749
timestamp 0
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_750
timestamp 0
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_751
timestamp 0
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_752
timestamp 0
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_753
timestamp 0
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_754
timestamp 0
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_755
timestamp 0
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_756
timestamp 0
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_757
timestamp 0
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_758
timestamp 0
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_759
timestamp 0
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_760
timestamp 0
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_761
timestamp 0
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_762
timestamp 0
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_763
timestamp 0
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_764
timestamp 0
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_765
timestamp 0
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_766
timestamp 0
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_767
timestamp 0
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_768
timestamp 0
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_769
timestamp 0
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_770
timestamp 0
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_771
timestamp 0
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_772
timestamp 0
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_773
timestamp 0
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_774
timestamp 0
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_775
timestamp 0
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_776
timestamp 0
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_777
timestamp 0
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_778
timestamp 0
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_779
timestamp 0
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_780
timestamp 0
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_781
timestamp 0
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_782
timestamp 0
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_783
timestamp 0
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_784
timestamp 0
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_785
timestamp 0
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_786
timestamp 0
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_787
timestamp 0
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_788
timestamp 0
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_789
timestamp 0
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_790
timestamp 0
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_791
timestamp 0
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_792
timestamp 0
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_793
timestamp 0
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_794
timestamp 0
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_795
timestamp 0
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_796
timestamp 0
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_797
timestamp 0
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_798
timestamp 0
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_799
timestamp 0
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_800
timestamp 0
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_801
timestamp 0
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_802
timestamp 0
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_803
timestamp 0
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_804
timestamp 0
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_805
timestamp 0
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_806
timestamp 0
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_807
timestamp 0
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_808
timestamp 0
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_809
timestamp 0
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_810
timestamp 0
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_811
timestamp 0
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_812
timestamp 0
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_813
timestamp 0
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_814
timestamp 0
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_815
timestamp 0
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_816
timestamp 0
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_817
timestamp 0
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_818
timestamp 0
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_819
timestamp 0
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_820
timestamp 0
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_821
timestamp 0
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_822
timestamp 0
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_823
timestamp 0
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_824
timestamp 0
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_825
timestamp 0
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_826
timestamp 0
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_827
timestamp 0
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_828
timestamp 0
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_829
timestamp 0
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_830
timestamp 0
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_831
timestamp 0
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_832
timestamp 0
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_833
timestamp 0
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_834
timestamp 0
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_835
timestamp 0
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_836
timestamp 0
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_837
timestamp 0
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_838
timestamp 0
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_839
timestamp 0
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_840
timestamp 0
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_841
timestamp 0
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_842
timestamp 0
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_843
timestamp 0
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_844
timestamp 0
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_845
timestamp 0
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_846
timestamp 0
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_847
timestamp 0
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_848
timestamp 0
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_849
timestamp 0
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_850
timestamp 0
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_851
timestamp 0
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_852
timestamp 0
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_853
timestamp 0
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_854
timestamp 0
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_855
timestamp 0
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_856
timestamp 0
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_857
timestamp 0
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_858
timestamp 0
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_859
timestamp 0
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_860
timestamp 0
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_861
timestamp 0
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_862
timestamp 0
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_863
timestamp 0
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_864
timestamp 0
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_865
timestamp 0
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_866
timestamp 0
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_867
timestamp 0
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_868
timestamp 0
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_869
timestamp 0
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_870
timestamp 0
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_871
timestamp 0
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_872
timestamp 0
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_873
timestamp 0
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_874
timestamp 0
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_875
timestamp 0
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_876
timestamp 0
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_877
timestamp 0
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_878
timestamp 0
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_879
timestamp 0
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_880
timestamp 0
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_881
timestamp 0
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_882
timestamp 0
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_883
timestamp 0
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_884
timestamp 0
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_885
timestamp 0
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_886
timestamp 0
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_887
timestamp 0
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_888
timestamp 0
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_889
timestamp 0
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_890
timestamp 0
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_891
timestamp 0
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_892
timestamp 0
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_893
timestamp 0
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_894
timestamp 0
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_895
timestamp 0
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_896
timestamp 0
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_897
timestamp 0
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_898
timestamp 0
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_899
timestamp 0
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_900
timestamp 0
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_901
timestamp 0
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_902
timestamp 0
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_903
timestamp 0
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_904
timestamp 0
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_905
timestamp 0
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_906
timestamp 0
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_907
timestamp 0
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_908
timestamp 0
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_909
timestamp 0
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_910
timestamp 0
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_911
timestamp 0
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_912
timestamp 0
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_913
timestamp 0
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_914
timestamp 0
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_915
timestamp 0
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_916
timestamp 0
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_917
timestamp 0
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_918
timestamp 0
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_919
timestamp 0
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_920
timestamp 0
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_921
timestamp 0
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_922
timestamp 0
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_923
timestamp 0
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_924
timestamp 0
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_925
timestamp 0
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_926
timestamp 0
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_927
timestamp 0
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_928
timestamp 0
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_929
timestamp 0
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_930
timestamp 0
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_931
timestamp 0
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_932
timestamp 0
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_933
timestamp 0
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_934
timestamp 0
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_935
timestamp 0
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_936
timestamp 0
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_937
timestamp 0
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_938
timestamp 0
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_939
timestamp 0
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_940
timestamp 0
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_941
timestamp 0
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_942
timestamp 0
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_943
timestamp 0
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_944
timestamp 0
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_945
timestamp 0
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_946
timestamp 0
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_947
timestamp 0
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_948
timestamp 0
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_949
timestamp 0
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_950
timestamp 0
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_951
timestamp 0
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_952
timestamp 0
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_953
timestamp 0
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_954
timestamp 0
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_955
timestamp 0
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_956
timestamp 0
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_957
timestamp 0
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_958
timestamp 0
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_959
timestamp 0
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_960
timestamp 0
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_961
timestamp 0
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_962
timestamp 0
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_963
timestamp 0
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_964
timestamp 0
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_965
timestamp 0
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_966
timestamp 0
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_967
timestamp 0
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_968
timestamp 0
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_969
timestamp 0
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_970
timestamp 0
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_971
timestamp 0
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_972
timestamp 0
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_973
timestamp 0
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_974
timestamp 0
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_975
timestamp 0
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_976
timestamp 0
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_977
timestamp 0
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_978
timestamp 0
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_979
timestamp 0
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_980
timestamp 0
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_981
timestamp 0
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_982
timestamp 0
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_983
timestamp 0
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_984
timestamp 0
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_985
timestamp 0
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_986
timestamp 0
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_987
timestamp 0
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_988
timestamp 0
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_989
timestamp 0
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_990
timestamp 0
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_991
timestamp 0
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_992
timestamp 0
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_993
timestamp 0
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_994
timestamp 0
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_995
timestamp 0
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_996
timestamp 0
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_997
timestamp 0
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_998
timestamp 0
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_999
timestamp 0
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1000
timestamp 0
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1001
timestamp 0
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1002
timestamp 0
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1003
timestamp 0
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1004
timestamp 0
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1005
timestamp 0
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1006
timestamp 0
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1007
timestamp 0
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1008
timestamp 0
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1009
timestamp 0
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1010
timestamp 0
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1011
timestamp 0
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1012
timestamp 0
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1013
timestamp 0
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1014
timestamp 0
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1015
timestamp 0
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1016
timestamp 0
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1017
timestamp 0
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1018
timestamp 0
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1019
timestamp 0
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1020
timestamp 0
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1021
timestamp 0
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1022
timestamp 0
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1023
timestamp 0
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1024
timestamp 0
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1025
timestamp 0
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1026
timestamp 0
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1027
timestamp 0
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1028
timestamp 0
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1029
timestamp 0
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1030
timestamp 0
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1031
timestamp 0
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1032
timestamp 0
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1033
timestamp 0
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1034
timestamp 0
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1035
timestamp 0
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1036
timestamp 0
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1037
timestamp 0
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1038
timestamp 0
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1039
timestamp 0
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1040
timestamp 0
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1041
timestamp 0
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1042
timestamp 0
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1043
timestamp 0
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1044
timestamp 0
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1045
timestamp 0
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1046
timestamp 0
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1047
timestamp 0
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1048
timestamp 0
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1049
timestamp 0
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1050
timestamp 0
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1051
timestamp 0
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1052
timestamp 0
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1053
timestamp 0
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1054
timestamp 0
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1055
timestamp 0
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1056
timestamp 0
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1057
timestamp 0
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1058
timestamp 0
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1059
timestamp 0
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1060
timestamp 0
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1061
timestamp 0
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1062
timestamp 0
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1063
timestamp 0
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1064
timestamp 0
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1065
timestamp 0
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1066
timestamp 0
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1067
timestamp 0
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1068
timestamp 0
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1069
timestamp 0
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1070
timestamp 0
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1071
timestamp 0
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1072
timestamp 0
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1073
timestamp 0
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1074
timestamp 0
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1075
timestamp 0
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1076
timestamp 0
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1077
timestamp 0
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1078
timestamp 0
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1079
timestamp 0
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1080
timestamp 0
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1081
timestamp 0
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1082
timestamp 0
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1083
timestamp 0
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1084
timestamp 0
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1085
timestamp 0
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1086
timestamp 0
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1087
timestamp 0
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1088
timestamp 0
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1089
timestamp 0
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1090
timestamp 0
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1091
timestamp 0
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1092
timestamp 0
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1093
timestamp 0
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1094
timestamp 0
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1095
timestamp 0
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1096
timestamp 0
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1097
timestamp 0
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1098
timestamp 0
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1099
timestamp 0
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1100
timestamp 0
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1101
timestamp 0
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1102
timestamp 0
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1103
timestamp 0
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1104
timestamp 0
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1105
timestamp 0
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1106
timestamp 0
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1107
timestamp 0
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1108
timestamp 0
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1109
timestamp 0
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1110
timestamp 0
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1111
timestamp 0
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1112
timestamp 0
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1113
timestamp 0
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1114
timestamp 0
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1115
timestamp 0
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1116
timestamp 0
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1117
timestamp 0
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1118
timestamp 0
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1119
timestamp 0
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1120
timestamp 0
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1121
timestamp 0
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1122
timestamp 0
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1123
timestamp 0
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1124
timestamp 0
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1125
timestamp 0
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1126
timestamp 0
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1127
timestamp 0
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1128
timestamp 0
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1129
timestamp 0
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1130
timestamp 0
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1131
timestamp 0
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1132
timestamp 0
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1133
timestamp 0
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1134
timestamp 0
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1135
timestamp 0
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1136
timestamp 0
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1137
timestamp 0
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1138
timestamp 0
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1139
timestamp 0
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1140
timestamp 0
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1141
timestamp 0
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1142
timestamp 0
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1143
timestamp 0
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1144
timestamp 0
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1145
timestamp 0
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1146
timestamp 0
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1147
timestamp 0
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1148
timestamp 0
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1149
timestamp 0
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1150
timestamp 0
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1151
timestamp 0
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1152
timestamp 0
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1153
timestamp 0
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1154
timestamp 0
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1155
timestamp 0
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1156
timestamp 0
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1157
timestamp 0
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1158
timestamp 0
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1159
timestamp 0
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1160
timestamp 0
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1161
timestamp 0
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1162
timestamp 0
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1163
timestamp 0
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1164
timestamp 0
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1165
timestamp 0
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1166
timestamp 0
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1167
timestamp 0
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1168
timestamp 0
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1169
timestamp 0
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1170
timestamp 0
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1171
timestamp 0
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1172
timestamp 0
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1173
timestamp 0
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1174
timestamp 0
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1175
timestamp 0
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1176
timestamp 0
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1177
timestamp 0
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1178
timestamp 0
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1179
timestamp 0
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1180
timestamp 0
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1181
timestamp 0
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1182
timestamp 0
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1183
timestamp 0
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1184
timestamp 0
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1185
timestamp 0
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1186
timestamp 0
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1187
timestamp 0
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1188
timestamp 0
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1189
timestamp 0
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1190
timestamp 0
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1191
timestamp 0
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1192
timestamp 0
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1193
timestamp 0
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1194
timestamp 0
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1195
timestamp 0
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1196
timestamp 0
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1197
timestamp 0
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1198
timestamp 0
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1199
timestamp 0
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1200
timestamp 0
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1201
timestamp 0
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1202
timestamp 0
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1203
timestamp 0
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1204
timestamp 0
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1205
timestamp 0
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1206
timestamp 0
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1207
timestamp 0
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1208
timestamp 0
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1209
timestamp 0
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1210
timestamp 0
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1211
timestamp 0
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1212
timestamp 0
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1213
timestamp 0
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1214
timestamp 0
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1215
timestamp 0
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1216
timestamp 0
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1217
timestamp 0
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1218
timestamp 0
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1219
timestamp 0
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1220
timestamp 0
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1221
timestamp 0
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1222
timestamp 0
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1223
timestamp 0
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1224
timestamp 0
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1225
timestamp 0
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1226
timestamp 0
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1227
timestamp 0
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1228
timestamp 0
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1229
timestamp 0
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1230
timestamp 0
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1231
timestamp 0
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1232
timestamp 0
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1233
timestamp 0
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1234
timestamp 0
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1235
timestamp 0
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1236
timestamp 0
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1237
timestamp 0
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1238
timestamp 0
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1239
timestamp 0
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1240
timestamp 0
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1241
timestamp 0
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1242
timestamp 0
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1243
timestamp 0
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1244
timestamp 0
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1245
timestamp 0
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1246
timestamp 0
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1247
timestamp 0
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1248
timestamp 0
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1249
timestamp 0
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1250
timestamp 0
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1251
timestamp 0
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1252
timestamp 0
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1253
timestamp 0
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1254
timestamp 0
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1255
timestamp 0
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1256
timestamp 0
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1257
timestamp 0
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1258
timestamp 0
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1259
timestamp 0
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1260
timestamp 0
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1261
timestamp 0
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1262
timestamp 0
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1263
timestamp 0
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1264
timestamp 0
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1265
timestamp 0
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1266
timestamp 0
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1267
timestamp 0
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1268
timestamp 0
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1269
timestamp 0
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1270
timestamp 0
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1271
timestamp 0
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1272
timestamp 0
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1273
timestamp 0
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1274
timestamp 0
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1275
timestamp 0
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1276
timestamp 0
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1277
timestamp 0
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1278
timestamp 0
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1279
timestamp 0
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1280
timestamp 0
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1281
timestamp 0
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1282
timestamp 0
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1283
timestamp 0
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1284
timestamp 0
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1285
timestamp 0
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1286
timestamp 0
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1287
timestamp 0
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1288
timestamp 0
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1289
timestamp 0
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1290
timestamp 0
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1291
timestamp 0
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1292
timestamp 0
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1293
timestamp 0
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1294
timestamp 0
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1295
timestamp 0
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1296
timestamp 0
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1297
timestamp 0
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1298
timestamp 0
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1299
timestamp 0
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1300
timestamp 0
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1301
timestamp 0
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1302
timestamp 0
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1303
timestamp 0
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1304
timestamp 0
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1305
timestamp 0
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1306
timestamp 0
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1307
timestamp 0
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1308
timestamp 0
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1309
timestamp 0
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1310
timestamp 0
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1311
timestamp 0
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1312
timestamp 0
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1313
timestamp 0
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1314
timestamp 0
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1315
timestamp 0
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1316
timestamp 0
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1317
timestamp 0
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1318
timestamp 0
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1319
timestamp 0
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1320
timestamp 0
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1321
timestamp 0
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1322
timestamp 0
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1323
timestamp 0
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1324
timestamp 0
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1325
timestamp 0
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1326
timestamp 0
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1327
timestamp 0
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1328
timestamp 0
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1329
timestamp 0
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1330
timestamp 0
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1331
timestamp 0
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1332
timestamp 0
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1333
timestamp 0
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1334
timestamp 0
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1335
timestamp 0
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1336
timestamp 0
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1337
timestamp 0
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1338
timestamp 0
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1339
timestamp 0
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1340
timestamp 0
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1341
timestamp 0
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1342
timestamp 0
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1343
timestamp 0
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1344
timestamp 0
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1345
timestamp 0
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1346
timestamp 0
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1347
timestamp 0
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  top_module_1
timestamp 0
transform 1 0 58328 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_2
timestamp 0
transform 1 0 58328 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_3
timestamp 0
transform 1 0 58328 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_4
timestamp 0
transform 1 0 58328 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_5
timestamp 0
transform 1 0 58328 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_6
timestamp 0
transform 1 0 58328 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_7
timestamp 0
transform 1 0 58328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_8
timestamp 0
transform 1 0 58328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_9
timestamp 0
transform 1 0 58328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_10
timestamp 0
transform 1 0 58328 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_11
timestamp 0
transform 1 0 58328 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_12
timestamp 0
transform 1 0 58328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_13
timestamp 0
transform 1 0 58328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_14
timestamp 0
transform 1 0 58328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_15
timestamp 0
transform 1 0 58328 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_16
timestamp 0
transform 1 0 58328 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_17
timestamp 0
transform 1 0 58328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_18
timestamp 0
transform 1 0 58328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_19
timestamp 0
transform 1 0 58328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_20
timestamp 0
transform 1 0 58328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_21
timestamp 0
transform 1 0 58328 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_22
timestamp 0
transform 1 0 58328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_23
timestamp 0
transform 1 0 58328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_24
timestamp 0
transform 1 0 58328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_25
timestamp 0
transform 1 0 58328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_26
timestamp 0
transform 1 0 58328 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_27
timestamp 0
transform 1 0 58328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_28
timestamp 0
transform 1 0 58328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_29
timestamp 0
transform 1 0 58328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_30
timestamp 0
transform 1 0 58328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_31
timestamp 0
transform 1 0 58328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_32
timestamp 0
transform 1 0 58328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_33
timestamp 0
transform 1 0 58328 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_34
timestamp 0
transform 1 0 58328 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_35
timestamp 0
transform 1 0 58328 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_36
timestamp 0
transform 1 0 58328 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_37
timestamp 0
transform 1 0 58328 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_38
timestamp 0
transform 1 0 58328 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_39
timestamp 0
transform 1 0 58328 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_40
timestamp 0
transform 1 0 58328 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_41
timestamp 0
transform 1 0 58328 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_42
timestamp 0
transform 1 0 58328 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_43
timestamp 0
transform 1 0 58328 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_44
timestamp 0
transform 1 0 58328 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_45
timestamp 0
transform 1 0 58328 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_46
timestamp 0
transform 1 0 58328 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_47
timestamp 0
transform 1 0 58328 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_48
timestamp 0
transform 1 0 58328 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_49
timestamp 0
transform 1 0 58328 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_50
timestamp 0
transform 1 0 58328 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_51
timestamp 0
transform 1 0 58328 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_52
timestamp 0
transform 1 0 58328 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_53
timestamp 0
transform 1 0 58328 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_54
timestamp 0
transform 1 0 58328 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_55
timestamp 0
transform 1 0 58328 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_56
timestamp 0
transform 1 0 58328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_57
timestamp 0
transform 1 0 58328 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_58
timestamp 0
transform 1 0 58328 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_59
timestamp 0
transform 1 0 58328 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_60
timestamp 0
transform 1 0 58328 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_61
timestamp 0
transform 1 0 58328 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_62
timestamp 0
transform 1 0 58328 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_63
timestamp 0
transform 1 0 58328 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  top_module_64
timestamp 0
transform 1 0 58328 0 1 30464
box -38 -48 314 592
<< labels >>
rlabel metal1 s 29992 57664 29992 57664 4 VGND
rlabel metal1 s 29992 57120 29992 57120 4 VPWR
rlabel metal2 s 58558 29529 58558 29529 4 net1
rlabel metal2 s 58558 22253 58558 22253 4 net10
rlabel metal3 s 58558 21301 58558 21301 4 net11
rlabel metal2 s 58558 20689 58558 20689 4 net12
rlabel metal2 s 58558 19737 58558 19737 4 net13
rlabel metal2 s 58558 18989 58558 18989 4 net14
rlabel metal3 s 58558 18037 58558 18037 4 net15
rlabel metal2 s 58558 17425 58558 17425 4 net16
rlabel metal1 s 58282 16626 58282 16626 4 net17
rlabel metal2 s 58558 15725 58558 15725 4 net18
rlabel metal3 s 58558 14773 58558 14773 4 net19
rlabel metal2 s 58558 28815 58558 28815 4 net2
rlabel metal2 s 58558 14161 58558 14161 4 net20
rlabel metal2 s 58558 13209 58558 13209 4 net21
rlabel metal2 s 58558 12461 58558 12461 4 net22
rlabel metal3 s 58558 11509 58558 11509 4 net23
rlabel metal2 s 58558 10897 58558 10897 4 net24
rlabel metal2 s 58558 9945 58558 9945 4 net25
rlabel metal2 s 58558 9197 58558 9197 4 net26
rlabel metal2 s 58558 8279 58558 8279 4 net27
rlabel metal2 s 58558 7633 58558 7633 4 net28
rlabel metal2 s 58558 6681 58558 6681 4 net29
rlabel metal3 s 58558 27829 58558 27829 4 net3
rlabel metal2 s 58558 5933 58558 5933 4 net30
rlabel metal3 s 58558 4981 58558 4981 4 net31
rlabel metal2 s 58558 4369 58558 4369 4 net32
rlabel metal2 s 58558 55641 58558 55641 4 net33
rlabel metal2 s 58558 54893 58558 54893 4 net34
rlabel metal3 s 58558 53941 58558 53941 4 net35
rlabel metal2 s 58558 53329 58558 53329 4 net36
rlabel metal2 s 58558 52377 58558 52377 4 net37
rlabel metal2 s 58558 51629 58558 51629 4 net38
rlabel metal3 s 58558 50677 58558 50677 4 net39
rlabel metal2 s 58558 27217 58558 27217 4 net4
rlabel metal2 s 58558 50065 58558 50065 4 net40
rlabel metal2 s 58558 49113 58558 49113 4 net41
rlabel metal2 s 58558 48365 58558 48365 4 net42
rlabel metal3 s 58558 47413 58558 47413 4 net43
rlabel metal2 s 58558 46801 58558 46801 4 net44
rlabel metal2 s 58558 45849 58558 45849 4 net45
rlabel metal2 s 58558 45101 58558 45101 4 net46
rlabel metal3 s 58558 44149 58558 44149 4 net47
rlabel metal2 s 58558 43537 58558 43537 4 net48
rlabel metal2 s 58558 42585 58558 42585 4 net49
rlabel metal3 s 58842 26180 58842 26180 4 net5
rlabel metal2 s 58558 41837 58558 41837 4 net50
rlabel metal3 s 58558 40885 58558 40885 4 net51
rlabel metal2 s 58558 40273 58558 40273 4 net52
rlabel metal2 s 58558 39321 58558 39321 4 net53
rlabel metal2 s 58558 38573 58558 38573 4 net54
rlabel metal3 s 58558 37621 58558 37621 4 net55
rlabel metal2 s 58558 37043 58558 37043 4 net56
rlabel metal2 s 58558 36057 58558 36057 4 net57
rlabel metal2 s 58558 35309 58558 35309 4 net58
rlabel metal3 s 58558 34357 58558 34357 4 net59
rlabel metal2 s 58558 25517 58558 25517 4 net6
rlabel metal2 s 58558 33745 58558 33745 4 net60
rlabel metal2 s 58558 32793 58558 32793 4 net61
rlabel metal2 s 58558 32045 58558 32045 4 net62
rlabel metal3 s 58558 31093 58558 31093 4 net63
rlabel metal2 s 58558 30481 58558 30481 4 net64
rlabel metal3 s 58558 24565 58558 24565 4 net7
rlabel metal2 s 58558 23953 58558 23953 4 net8
rlabel metal2 s 58558 23001 58558 23001 4 net9
flabel metal5 s 1056 53676 58928 53996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 48676 58928 48996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 43676 58928 43996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 38676 58928 38996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 33676 58928 33996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 28676 58928 28996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 23676 58928 23996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 18676 58928 18996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 13676 58928 13996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8676 58928 8996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3676 58928 3996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 57604 2128 57924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 52604 2128 52924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 47604 2128 47924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 42604 2128 42924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 37604 2128 37924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 32604 2128 32924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 27604 2128 27924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 22604 2128 22924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 17604 2128 17924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 12604 2128 12924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7604 2128 7924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2604 2128 2924 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 53016 58928 53336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 48016 58928 48336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 43016 58928 43336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 38016 58928 38336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 33016 58928 33336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 28016 58928 28336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 23016 58928 23336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 18016 58928 18336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 13016 58928 13336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 8016 58928 8336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3016 58928 3336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 56944 2128 57264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 51944 2128 52264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 46944 2128 47264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 41944 2128 42264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 36944 2128 37264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 31944 2128 32264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 26944 2128 27264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 21944 2128 22264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 16944 2128 17264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 11944 2128 12264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 6944 2128 7264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1944 2128 2264 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 10072 800 10192 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 0 49784 800 49904 0 FreeSans 600 0 0 0 control
port 4 nsew
flabel metal3 s 0 29928 800 30048 0 FreeSans 600 0 0 0 reset
port 5 nsew
flabel metal3 s 59200 29384 60000 29504 0 FreeSans 600 0 0 0 result1[0]
port 6 nsew
flabel metal3 s 59200 21224 60000 21344 0 FreeSans 600 0 0 0 result1[10]
port 7 nsew
flabel metal3 s 59200 20408 60000 20528 0 FreeSans 600 0 0 0 result1[11]
port 8 nsew
flabel metal3 s 59200 19592 60000 19712 0 FreeSans 600 0 0 0 result1[12]
port 9 nsew
flabel metal3 s 59200 18776 60000 18896 0 FreeSans 600 0 0 0 result1[13]
port 10 nsew
flabel metal3 s 59200 17960 60000 18080 0 FreeSans 600 0 0 0 result1[14]
port 11 nsew
flabel metal3 s 59200 17144 60000 17264 0 FreeSans 600 0 0 0 result1[15]
port 12 nsew
flabel metal3 s 59200 16328 60000 16448 0 FreeSans 600 0 0 0 result1[16]
port 13 nsew
flabel metal3 s 59200 15512 60000 15632 0 FreeSans 600 0 0 0 result1[17]
port 14 nsew
flabel metal3 s 59200 14696 60000 14816 0 FreeSans 600 0 0 0 result1[18]
port 15 nsew
flabel metal3 s 59200 13880 60000 14000 0 FreeSans 600 0 0 0 result1[19]
port 16 nsew
flabel metal3 s 59200 28568 60000 28688 0 FreeSans 600 0 0 0 result1[1]
port 17 nsew
flabel metal3 s 59200 13064 60000 13184 0 FreeSans 600 0 0 0 result1[20]
port 18 nsew
flabel metal3 s 59200 12248 60000 12368 0 FreeSans 600 0 0 0 result1[21]
port 19 nsew
flabel metal3 s 59200 11432 60000 11552 0 FreeSans 600 0 0 0 result1[22]
port 20 nsew
flabel metal3 s 59200 10616 60000 10736 0 FreeSans 600 0 0 0 result1[23]
port 21 nsew
flabel metal3 s 59200 9800 60000 9920 0 FreeSans 600 0 0 0 result1[24]
port 22 nsew
flabel metal3 s 59200 8984 60000 9104 0 FreeSans 600 0 0 0 result1[25]
port 23 nsew
flabel metal3 s 59200 8168 60000 8288 0 FreeSans 600 0 0 0 result1[26]
port 24 nsew
flabel metal3 s 59200 7352 60000 7472 0 FreeSans 600 0 0 0 result1[27]
port 25 nsew
flabel metal3 s 59200 6536 60000 6656 0 FreeSans 600 0 0 0 result1[28]
port 26 nsew
flabel metal3 s 59200 5720 60000 5840 0 FreeSans 600 0 0 0 result1[29]
port 27 nsew
flabel metal3 s 59200 27752 60000 27872 0 FreeSans 600 0 0 0 result1[2]
port 28 nsew
flabel metal3 s 59200 4904 60000 5024 0 FreeSans 600 0 0 0 result1[30]
port 29 nsew
flabel metal3 s 59200 4088 60000 4208 0 FreeSans 600 0 0 0 result1[31]
port 30 nsew
flabel metal3 s 59200 26936 60000 27056 0 FreeSans 600 0 0 0 result1[3]
port 31 nsew
flabel metal3 s 59200 26120 60000 26240 0 FreeSans 600 0 0 0 result1[4]
port 32 nsew
flabel metal3 s 59200 25304 60000 25424 0 FreeSans 600 0 0 0 result1[5]
port 33 nsew
flabel metal3 s 59200 24488 60000 24608 0 FreeSans 600 0 0 0 result1[6]
port 34 nsew
flabel metal3 s 59200 23672 60000 23792 0 FreeSans 600 0 0 0 result1[7]
port 35 nsew
flabel metal3 s 59200 22856 60000 22976 0 FreeSans 600 0 0 0 result1[8]
port 36 nsew
flabel metal3 s 59200 22040 60000 22160 0 FreeSans 600 0 0 0 result1[9]
port 37 nsew
flabel metal3 s 59200 55496 60000 55616 0 FreeSans 600 0 0 0 result2[0]
port 38 nsew
flabel metal3 s 59200 47336 60000 47456 0 FreeSans 600 0 0 0 result2[10]
port 39 nsew
flabel metal3 s 59200 46520 60000 46640 0 FreeSans 600 0 0 0 result2[11]
port 40 nsew
flabel metal3 s 59200 45704 60000 45824 0 FreeSans 600 0 0 0 result2[12]
port 41 nsew
flabel metal3 s 59200 44888 60000 45008 0 FreeSans 600 0 0 0 result2[13]
port 42 nsew
flabel metal3 s 59200 44072 60000 44192 0 FreeSans 600 0 0 0 result2[14]
port 43 nsew
flabel metal3 s 59200 43256 60000 43376 0 FreeSans 600 0 0 0 result2[15]
port 44 nsew
flabel metal3 s 59200 42440 60000 42560 0 FreeSans 600 0 0 0 result2[16]
port 45 nsew
flabel metal3 s 59200 41624 60000 41744 0 FreeSans 600 0 0 0 result2[17]
port 46 nsew
flabel metal3 s 59200 40808 60000 40928 0 FreeSans 600 0 0 0 result2[18]
port 47 nsew
flabel metal3 s 59200 39992 60000 40112 0 FreeSans 600 0 0 0 result2[19]
port 48 nsew
flabel metal3 s 59200 54680 60000 54800 0 FreeSans 600 0 0 0 result2[1]
port 49 nsew
flabel metal3 s 59200 39176 60000 39296 0 FreeSans 600 0 0 0 result2[20]
port 50 nsew
flabel metal3 s 59200 38360 60000 38480 0 FreeSans 600 0 0 0 result2[21]
port 51 nsew
flabel metal3 s 59200 37544 60000 37664 0 FreeSans 600 0 0 0 result2[22]
port 52 nsew
flabel metal3 s 59200 36728 60000 36848 0 FreeSans 600 0 0 0 result2[23]
port 53 nsew
flabel metal3 s 59200 35912 60000 36032 0 FreeSans 600 0 0 0 result2[24]
port 54 nsew
flabel metal3 s 59200 35096 60000 35216 0 FreeSans 600 0 0 0 result2[25]
port 55 nsew
flabel metal3 s 59200 34280 60000 34400 0 FreeSans 600 0 0 0 result2[26]
port 56 nsew
flabel metal3 s 59200 33464 60000 33584 0 FreeSans 600 0 0 0 result2[27]
port 57 nsew
flabel metal3 s 59200 32648 60000 32768 0 FreeSans 600 0 0 0 result2[28]
port 58 nsew
flabel metal3 s 59200 31832 60000 31952 0 FreeSans 600 0 0 0 result2[29]
port 59 nsew
flabel metal3 s 59200 53864 60000 53984 0 FreeSans 600 0 0 0 result2[2]
port 60 nsew
flabel metal3 s 59200 31016 60000 31136 0 FreeSans 600 0 0 0 result2[30]
port 61 nsew
flabel metal3 s 59200 30200 60000 30320 0 FreeSans 600 0 0 0 result2[31]
port 62 nsew
flabel metal3 s 59200 53048 60000 53168 0 FreeSans 600 0 0 0 result2[3]
port 63 nsew
flabel metal3 s 59200 52232 60000 52352 0 FreeSans 600 0 0 0 result2[4]
port 64 nsew
flabel metal3 s 59200 51416 60000 51536 0 FreeSans 600 0 0 0 result2[5]
port 65 nsew
flabel metal3 s 59200 50600 60000 50720 0 FreeSans 600 0 0 0 result2[6]
port 66 nsew
flabel metal3 s 59200 49784 60000 49904 0 FreeSans 600 0 0 0 result2[7]
port 67 nsew
flabel metal3 s 59200 48968 60000 49088 0 FreeSans 600 0 0 0 result2[8]
port 68 nsew
flabel metal3 s 59200 48152 60000 48272 0 FreeSans 600 0 0 0 result2[9]
port 69 nsew
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
